// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_ddr_east
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_ddr_east_p (
    output logic [182:0]                                 o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data,
    output logic                                         o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head,
    input  logic                                         i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy,
    output logic                                         o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail,
    output logic                                         o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld,
    input  logic [182:0]                                 i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data,
    input  logic                                         i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head,
    output logic                                         o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy,
    input  logic                                         i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail,
    input  logic                                         i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld,
    input  logic [398:0]                                 i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld,
    output logic [398:0]                                 o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld,
    input  logic [398:0]                                 i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld,
    output logic [398:0]                                 o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld,
    input  logic [398:0]                                 i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld,
    output logic [398:0]                                 o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld,
    input  logic [398:0]                                 i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld,
    output logic [398:0]                                 o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld,
    input  logic [182:0]                                 i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld,
    output logic [182:0]                                 o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld,
    input  logic                                         i_l2_addr_mode_port_b0,
    input  logic                                         i_l2_addr_mode_port_b1,
    input  logic                                         i_l2_intr_mode_port_b0,
    input  logic                                         i_l2_intr_mode_port_b1,
    input  logic                                         i_lpddr_graph_addr_mode_port_b0,
    input  logic                                         i_lpddr_graph_addr_mode_port_b1,
    input  logic                                         i_lpddr_graph_intr_mode_port_b0,
    input  logic                                         i_lpddr_graph_intr_mode_port_b1,
    input  wire                                          i_lpddr_ppp_0_aon_clk,
    input  wire                                          i_lpddr_ppp_0_aon_rst_n,
    output logic                                         o_lpddr_ppp_0_cfg_pwr_idle_val,
    output logic                                         o_lpddr_ppp_0_cfg_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_0_cfg_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_0_clk,
    input  wire                                          i_lpddr_ppp_0_clken,
    output logic                                         o_lpddr_ppp_0_pwr_idle_val,
    output logic                                         o_lpddr_ppp_0_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_0_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_0_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t     o_lpddr_ppp_0_targ_cfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_0_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_0_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     i_lpddr_ppp_0_targ_cfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_0_targ_cfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_0_targ_cfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_0_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                   o_lpddr_ppp_0_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     o_lpddr_ppp_0_targ_cfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_0_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_0_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_0_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_0_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_0_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_0_targ_mt_axi_m_arlen,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_0_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_0_targ_mt_axi_m_arqos,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_0_targ_mt_axi_m_arsize,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_0_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_0_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_0_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_0_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_0_targ_mt_axi_m_awlen,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_0_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_0_targ_mt_axi_m_awqos,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_0_targ_mt_axi_m_awsize,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_0_targ_mt_axi_m_bid,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_0_targ_mt_axi_m_bresp,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       i_lpddr_ppp_0_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_0_targ_mt_axi_m_rid,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_rlast,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_0_targ_mt_axi_m_rresp,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       o_lpddr_ppp_0_targ_mt_axi_m_wdata,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_wlast,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t       o_lpddr_ppp_0_targ_mt_axi_m_wstrb,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_lpddr_ppp_0_targ_syscfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_lpddr_ppp_0_targ_syscfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_0_targ_syscfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_0_targ_syscfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_lpddr_ppp_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_lpddr_ppp_0_targ_syscfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_0_targ_syscfg_apb_m_pwrite,
    input  wire                                          i_lpddr_ppp_1_aon_clk,
    input  wire                                          i_lpddr_ppp_1_aon_rst_n,
    output logic                                         o_lpddr_ppp_1_cfg_pwr_idle_val,
    output logic                                         o_lpddr_ppp_1_cfg_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_1_cfg_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_1_clk,
    input  wire                                          i_lpddr_ppp_1_clken,
    output logic                                         o_lpddr_ppp_1_pwr_idle_val,
    output logic                                         o_lpddr_ppp_1_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_1_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_1_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t     o_lpddr_ppp_1_targ_cfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_1_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_1_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     i_lpddr_ppp_1_targ_cfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_1_targ_cfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_1_targ_cfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_1_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                   o_lpddr_ppp_1_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     o_lpddr_ppp_1_targ_cfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_1_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_1_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_1_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_1_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_1_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_1_targ_mt_axi_m_arlen,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_1_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_1_targ_mt_axi_m_arqos,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_1_targ_mt_axi_m_arsize,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_1_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_1_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_1_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_1_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_1_targ_mt_axi_m_awlen,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_1_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_1_targ_mt_axi_m_awqos,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_1_targ_mt_axi_m_awsize,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_1_targ_mt_axi_m_bid,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_1_targ_mt_axi_m_bresp,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       i_lpddr_ppp_1_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_1_targ_mt_axi_m_rid,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_rlast,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_1_targ_mt_axi_m_rresp,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       o_lpddr_ppp_1_targ_mt_axi_m_wdata,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_wlast,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t       o_lpddr_ppp_1_targ_mt_axi_m_wstrb,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_lpddr_ppp_1_targ_syscfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_lpddr_ppp_1_targ_syscfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_1_targ_syscfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_1_targ_syscfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_lpddr_ppp_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_lpddr_ppp_1_targ_syscfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_1_targ_syscfg_apb_m_pwrite,
    input  wire                                          i_lpddr_ppp_2_aon_clk,
    input  wire                                          i_lpddr_ppp_2_aon_rst_n,
    output logic                                         o_lpddr_ppp_2_cfg_pwr_idle_val,
    output logic                                         o_lpddr_ppp_2_cfg_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_2_cfg_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_2_clk,
    input  wire                                          i_lpddr_ppp_2_clken,
    output logic                                         o_lpddr_ppp_2_pwr_idle_val,
    output logic                                         o_lpddr_ppp_2_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_2_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_2_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t     o_lpddr_ppp_2_targ_cfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_2_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_2_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     i_lpddr_ppp_2_targ_cfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_2_targ_cfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_2_targ_cfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_2_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                   o_lpddr_ppp_2_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     o_lpddr_ppp_2_targ_cfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_2_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_2_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_2_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_2_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_2_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_2_targ_mt_axi_m_arlen,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_2_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_2_targ_mt_axi_m_arqos,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_2_targ_mt_axi_m_arsize,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_2_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_2_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_2_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_2_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_2_targ_mt_axi_m_awlen,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_2_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_2_targ_mt_axi_m_awqos,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_2_targ_mt_axi_m_awsize,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_2_targ_mt_axi_m_bid,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_2_targ_mt_axi_m_bresp,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       i_lpddr_ppp_2_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_2_targ_mt_axi_m_rid,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_rlast,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_2_targ_mt_axi_m_rresp,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       o_lpddr_ppp_2_targ_mt_axi_m_wdata,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_wlast,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t       o_lpddr_ppp_2_targ_mt_axi_m_wstrb,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_lpddr_ppp_2_targ_syscfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_lpddr_ppp_2_targ_syscfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_2_targ_syscfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_2_targ_syscfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_lpddr_ppp_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_lpddr_ppp_2_targ_syscfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_2_targ_syscfg_apb_m_pwrite,
    input  wire                                          i_lpddr_ppp_3_aon_clk,
    input  wire                                          i_lpddr_ppp_3_aon_rst_n,
    output logic                                         o_lpddr_ppp_3_cfg_pwr_idle_val,
    output logic                                         o_lpddr_ppp_3_cfg_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_3_cfg_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_3_clk,
    input  wire                                          i_lpddr_ppp_3_clken,
    output logic                                         o_lpddr_ppp_3_pwr_idle_val,
    output logic                                         o_lpddr_ppp_3_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_3_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_3_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t     o_lpddr_ppp_3_targ_cfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_3_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_3_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     i_lpddr_ppp_3_targ_cfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_3_targ_cfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_3_targ_cfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_3_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                   o_lpddr_ppp_3_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     o_lpddr_ppp_3_targ_cfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_3_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_3_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_3_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_3_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_3_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_3_targ_mt_axi_m_arlen,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_3_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_3_targ_mt_axi_m_arqos,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_3_targ_mt_axi_m_arsize,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_3_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_3_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_3_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_3_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_3_targ_mt_axi_m_awlen,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_3_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_3_targ_mt_axi_m_awqos,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_3_targ_mt_axi_m_awsize,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_3_targ_mt_axi_m_bid,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_3_targ_mt_axi_m_bresp,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       i_lpddr_ppp_3_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_3_targ_mt_axi_m_rid,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_rlast,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_3_targ_mt_axi_m_rresp,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       o_lpddr_ppp_3_targ_mt_axi_m_wdata,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_wlast,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t       o_lpddr_ppp_3_targ_mt_axi_m_wstrb,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_lpddr_ppp_3_targ_syscfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_lpddr_ppp_3_targ_syscfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_3_targ_syscfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_3_targ_syscfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_lpddr_ppp_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_lpddr_ppp_3_targ_syscfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_3_targ_syscfg_apb_m_pwrite,
    input  logic                                         i_lpddr_ppp_addr_mode_port_b0,
    input  logic                                         i_lpddr_ppp_addr_mode_port_b1,
    input  logic                                         i_lpddr_ppp_intr_mode_port_b0,
    input  logic                                         i_lpddr_ppp_intr_mode_port_b1,
    input  wire                                          i_noc_clk,
    input  wire                                          i_noc_rst_n,
    input  wire                                          i_soc_periph_aon_clk,
    input  wire                                          i_soc_periph_aon_rst_n,
    input  wire                                          i_soc_periph_clk,
    input  wire                                          i_soc_periph_clken,
    input  chip_pkg::chip_axi_addr_t                     i_soc_periph_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                          i_soc_periph_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                          i_soc_periph_init_lt_axi_s_arcache,
    input  soc_periph_pkg::soc_periph_init_lt_axi_id_t   i_soc_periph_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                            i_soc_periph_init_lt_axi_s_arlen,
    input  logic                                         i_soc_periph_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                           i_soc_periph_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                            i_soc_periph_init_lt_axi_s_arqos,
    output logic                                         o_soc_periph_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                           i_soc_periph_init_lt_axi_s_arsize,
    input  logic                                         i_soc_periph_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                     i_soc_periph_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                          i_soc_periph_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                          i_soc_periph_init_lt_axi_s_awcache,
    input  soc_periph_pkg::soc_periph_init_lt_axi_id_t   i_soc_periph_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                            i_soc_periph_init_lt_axi_s_awlen,
    input  logic                                         i_soc_periph_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                           i_soc_periph_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                            i_soc_periph_init_lt_axi_s_awqos,
    output logic                                         o_soc_periph_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                           i_soc_periph_init_lt_axi_s_awsize,
    input  logic                                         i_soc_periph_init_lt_axi_s_awvalid,
    output soc_periph_pkg::soc_periph_init_lt_axi_id_t   o_soc_periph_init_lt_axi_s_bid,
    input  logic                                         i_soc_periph_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                           o_soc_periph_init_lt_axi_s_bresp,
    output logic                                         o_soc_periph_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                  o_soc_periph_init_lt_axi_s_rdata,
    output soc_periph_pkg::soc_periph_init_lt_axi_id_t   o_soc_periph_init_lt_axi_s_rid,
    output logic                                         o_soc_periph_init_lt_axi_s_rlast,
    input  logic                                         i_soc_periph_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                           o_soc_periph_init_lt_axi_s_rresp,
    output logic                                         o_soc_periph_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                  i_soc_periph_init_lt_axi_s_wdata,
    input  logic                                         i_soc_periph_init_lt_axi_s_wlast,
    output logic                                         o_soc_periph_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                 i_soc_periph_init_lt_axi_s_wstrb,
    input  logic                                         i_soc_periph_init_lt_axi_s_wvalid,
    output logic                                         o_soc_periph_pwr_idle_val,
    output logic                                         o_soc_periph_pwr_idle_ack,
    input  logic                                         i_soc_periph_pwr_idle_req,
    input  wire                                          i_soc_periph_rst_n,
    output chip_pkg::chip_axi_addr_t                     o_soc_periph_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_soc_periph_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_soc_periph_targ_lt_axi_m_arcache,
    output soc_periph_pkg::soc_periph_targ_lt_axi_id_t   o_soc_periph_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_soc_periph_targ_lt_axi_m_arlen,
    output logic                                         o_soc_periph_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_soc_periph_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_soc_periph_targ_lt_axi_m_arqos,
    input  logic                                         i_soc_periph_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_soc_periph_targ_lt_axi_m_arsize,
    output logic                                         o_soc_periph_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_soc_periph_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_soc_periph_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_soc_periph_targ_lt_axi_m_awcache,
    output soc_periph_pkg::soc_periph_targ_lt_axi_id_t   o_soc_periph_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_soc_periph_targ_lt_axi_m_awlen,
    output logic                                         o_soc_periph_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_soc_periph_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_soc_periph_targ_lt_axi_m_awqos,
    input  logic                                         i_soc_periph_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_soc_periph_targ_lt_axi_m_awsize,
    output logic                                         o_soc_periph_targ_lt_axi_m_awvalid,
    input  soc_periph_pkg::soc_periph_targ_lt_axi_id_t   i_soc_periph_targ_lt_axi_m_bid,
    output logic                                         o_soc_periph_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_soc_periph_targ_lt_axi_m_bresp,
    input  logic                                         i_soc_periph_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                  i_soc_periph_targ_lt_axi_m_rdata,
    input  soc_periph_pkg::soc_periph_targ_lt_axi_id_t   i_soc_periph_targ_lt_axi_m_rid,
    input  logic                                         i_soc_periph_targ_lt_axi_m_rlast,
    output logic                                         o_soc_periph_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_soc_periph_targ_lt_axi_m_rresp,
    input  logic                                         i_soc_periph_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                  o_soc_periph_targ_lt_axi_m_wdata,
    output logic                                         o_soc_periph_targ_lt_axi_m_wlast,
    input  logic                                         i_soc_periph_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                 o_soc_periph_targ_lt_axi_m_wstrb,
    output logic                                         o_soc_periph_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_soc_periph_targ_syscfg_apb_m_paddr,
    output logic                                         o_soc_periph_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_soc_periph_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_soc_periph_targ_syscfg_apb_m_prdata,
    input  logic                                         i_soc_periph_targ_syscfg_apb_m_pready,
    output logic                                         o_soc_periph_targ_syscfg_apb_m_psel,
    input  logic                                         i_soc_periph_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_soc_periph_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_soc_periph_targ_syscfg_apb_m_pwdata,
    output logic                                         o_soc_periph_targ_syscfg_apb_m_pwrite,
    // DFT Interface
    input  wire           tck,
    input  wire           trst,
    input  logic          tms,
    input  logic          tdi,
    output logic          tdo_en,
    output logic          tdo,
    input  wire           test_clk,
    input  logic          test_mode,
    input  logic          edt_update,
    input  logic          scan_en,
    input  logic [12-1:0] scan_in,
    output logic [12-1:0] scan_out
);
    // -- Automatically-generated Reset Synchronizers -- //
    wire lpddr_ppp_0_aon_rst_n_synced;
    wire lpddr_ppp_1_aon_rst_n_synced;
    wire lpddr_ppp_2_aon_rst_n_synced;
    wire lpddr_ppp_3_aon_rst_n_synced;
    wire soc_periph_aon_rst_n_synced;

    // LPDDR PPP 0 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_lpddr_ppp_0_aon_rst_n_sync (
        .i_clk          (i_lpddr_ppp_0_aon_clk),
        .i_rst_n        (i_lpddr_ppp_0_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (lpddr_ppp_0_aon_rst_n_synced)
    );

    // LPDDR PPP 1 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_lpddr_ppp_1_aon_rst_n_sync (
        .i_clk          (i_lpddr_ppp_1_aon_clk),
        .i_rst_n        (i_lpddr_ppp_1_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (lpddr_ppp_1_aon_rst_n_synced)
    );

    // LPDDR PPP 2 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_lpddr_ppp_2_aon_rst_n_sync (
        .i_clk          (i_lpddr_ppp_2_aon_clk),
        .i_rst_n        (i_lpddr_ppp_2_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (lpddr_ppp_2_aon_rst_n_synced)
    );

    // LPDDR PPP 3 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_lpddr_ppp_3_aon_rst_n_sync (
        .i_clk          (i_lpddr_ppp_3_aon_clk),
        .i_rst_n        (i_lpddr_ppp_3_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (lpddr_ppp_3_aon_rst_n_synced)
    );

    // SOC PERIPH AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_soc_periph_aon_rst_n_sync (
        .i_clk          (i_soc_periph_aon_clk),
        .i_rst_n        (i_soc_periph_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (soc_periph_aon_rst_n_synced)
    );

    noc_ddr_east u_noc_ddr_east (
    .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data),
    .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head),
    .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy),
    .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail),
    .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld),
    .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data),
    .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head),
    .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy),
    .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail),
    .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data),
    .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head),
    .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data),
    .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head),
    .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld),
    .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .i_lpddr_ppp_0_aon_clk(i_lpddr_ppp_0_aon_clk),
    .i_lpddr_ppp_0_aon_rst_n(lpddr_ppp_0_aon_rst_n_synced),
    .o_lpddr_ppp_0_cfg_pwr_idle_val(o_lpddr_ppp_0_cfg_pwr_idle_val),
    .o_lpddr_ppp_0_cfg_pwr_idle_ack(o_lpddr_ppp_0_cfg_pwr_idle_ack),
    .i_lpddr_ppp_0_cfg_pwr_idle_req(i_lpddr_ppp_0_cfg_pwr_idle_req),
    .i_lpddr_ppp_0_clk(i_lpddr_ppp_0_clk),
    .i_lpddr_ppp_0_clken(i_lpddr_ppp_0_clken),
    .o_lpddr_ppp_0_pwr_idle_val(o_lpddr_ppp_0_pwr_idle_val),
    .o_lpddr_ppp_0_pwr_idle_ack(o_lpddr_ppp_0_pwr_idle_ack),
    .i_lpddr_ppp_0_pwr_idle_req(i_lpddr_ppp_0_pwr_idle_req),
    .i_lpddr_ppp_0_rst_n(i_lpddr_ppp_0_rst_n),
    .o_lpddr_ppp_0_targ_cfg_apb_m_paddr(o_lpddr_ppp_0_targ_cfg_apb_m_paddr),
    .o_lpddr_ppp_0_targ_cfg_apb_m_penable(o_lpddr_ppp_0_targ_cfg_apb_m_penable),
    .o_lpddr_ppp_0_targ_cfg_apb_m_pprot(o_lpddr_ppp_0_targ_cfg_apb_m_pprot),
    .i_lpddr_ppp_0_targ_cfg_apb_m_prdata(i_lpddr_ppp_0_targ_cfg_apb_m_prdata),
    .i_lpddr_ppp_0_targ_cfg_apb_m_pready(i_lpddr_ppp_0_targ_cfg_apb_m_pready),
    .o_lpddr_ppp_0_targ_cfg_apb_m_psel(o_lpddr_ppp_0_targ_cfg_apb_m_psel),
    .i_lpddr_ppp_0_targ_cfg_apb_m_pslverr(i_lpddr_ppp_0_targ_cfg_apb_m_pslverr),
    .o_lpddr_ppp_0_targ_cfg_apb_m_pstrb(o_lpddr_ppp_0_targ_cfg_apb_m_pstrb),
    .o_lpddr_ppp_0_targ_cfg_apb_m_pwdata(o_lpddr_ppp_0_targ_cfg_apb_m_pwdata),
    .o_lpddr_ppp_0_targ_cfg_apb_m_pwrite(o_lpddr_ppp_0_targ_cfg_apb_m_pwrite),
    .o_lpddr_ppp_0_targ_mt_axi_m_araddr(o_lpddr_ppp_0_targ_mt_axi_m_araddr),
    .o_lpddr_ppp_0_targ_mt_axi_m_arburst(o_lpddr_ppp_0_targ_mt_axi_m_arburst),
    .o_lpddr_ppp_0_targ_mt_axi_m_arcache(o_lpddr_ppp_0_targ_mt_axi_m_arcache),
    .o_lpddr_ppp_0_targ_mt_axi_m_arid(o_lpddr_ppp_0_targ_mt_axi_m_arid),
    .o_lpddr_ppp_0_targ_mt_axi_m_arlen(o_lpddr_ppp_0_targ_mt_axi_m_arlen),
    .o_lpddr_ppp_0_targ_mt_axi_m_arlock(o_lpddr_ppp_0_targ_mt_axi_m_arlock),
    .o_lpddr_ppp_0_targ_mt_axi_m_arprot(o_lpddr_ppp_0_targ_mt_axi_m_arprot),
    .o_lpddr_ppp_0_targ_mt_axi_m_arqos(o_lpddr_ppp_0_targ_mt_axi_m_arqos),
    .i_lpddr_ppp_0_targ_mt_axi_m_arready(i_lpddr_ppp_0_targ_mt_axi_m_arready),
    .o_lpddr_ppp_0_targ_mt_axi_m_arsize(o_lpddr_ppp_0_targ_mt_axi_m_arsize),
    .o_lpddr_ppp_0_targ_mt_axi_m_arvalid(o_lpddr_ppp_0_targ_mt_axi_m_arvalid),
    .o_lpddr_ppp_0_targ_mt_axi_m_awaddr(o_lpddr_ppp_0_targ_mt_axi_m_awaddr),
    .o_lpddr_ppp_0_targ_mt_axi_m_awburst(o_lpddr_ppp_0_targ_mt_axi_m_awburst),
    .o_lpddr_ppp_0_targ_mt_axi_m_awcache(o_lpddr_ppp_0_targ_mt_axi_m_awcache),
    .o_lpddr_ppp_0_targ_mt_axi_m_awid(o_lpddr_ppp_0_targ_mt_axi_m_awid),
    .o_lpddr_ppp_0_targ_mt_axi_m_awlen(o_lpddr_ppp_0_targ_mt_axi_m_awlen),
    .o_lpddr_ppp_0_targ_mt_axi_m_awlock(o_lpddr_ppp_0_targ_mt_axi_m_awlock),
    .o_lpddr_ppp_0_targ_mt_axi_m_awprot(o_lpddr_ppp_0_targ_mt_axi_m_awprot),
    .o_lpddr_ppp_0_targ_mt_axi_m_awqos(o_lpddr_ppp_0_targ_mt_axi_m_awqos),
    .i_lpddr_ppp_0_targ_mt_axi_m_awready(i_lpddr_ppp_0_targ_mt_axi_m_awready),
    .o_lpddr_ppp_0_targ_mt_axi_m_awsize(o_lpddr_ppp_0_targ_mt_axi_m_awsize),
    .o_lpddr_ppp_0_targ_mt_axi_m_awvalid(o_lpddr_ppp_0_targ_mt_axi_m_awvalid),
    .i_lpddr_ppp_0_targ_mt_axi_m_bid(i_lpddr_ppp_0_targ_mt_axi_m_bid),
    .o_lpddr_ppp_0_targ_mt_axi_m_bready(o_lpddr_ppp_0_targ_mt_axi_m_bready),
    .i_lpddr_ppp_0_targ_mt_axi_m_bresp(i_lpddr_ppp_0_targ_mt_axi_m_bresp),
    .i_lpddr_ppp_0_targ_mt_axi_m_bvalid(i_lpddr_ppp_0_targ_mt_axi_m_bvalid),
    .i_lpddr_ppp_0_targ_mt_axi_m_rdata(i_lpddr_ppp_0_targ_mt_axi_m_rdata),
    .i_lpddr_ppp_0_targ_mt_axi_m_rid(i_lpddr_ppp_0_targ_mt_axi_m_rid),
    .i_lpddr_ppp_0_targ_mt_axi_m_rlast(i_lpddr_ppp_0_targ_mt_axi_m_rlast),
    .o_lpddr_ppp_0_targ_mt_axi_m_rready(o_lpddr_ppp_0_targ_mt_axi_m_rready),
    .i_lpddr_ppp_0_targ_mt_axi_m_rresp(i_lpddr_ppp_0_targ_mt_axi_m_rresp),
    .i_lpddr_ppp_0_targ_mt_axi_m_rvalid(i_lpddr_ppp_0_targ_mt_axi_m_rvalid),
    .o_lpddr_ppp_0_targ_mt_axi_m_wdata(o_lpddr_ppp_0_targ_mt_axi_m_wdata),
    .o_lpddr_ppp_0_targ_mt_axi_m_wlast(o_lpddr_ppp_0_targ_mt_axi_m_wlast),
    .i_lpddr_ppp_0_targ_mt_axi_m_wready(i_lpddr_ppp_0_targ_mt_axi_m_wready),
    .o_lpddr_ppp_0_targ_mt_axi_m_wstrb(o_lpddr_ppp_0_targ_mt_axi_m_wstrb),
    .o_lpddr_ppp_0_targ_mt_axi_m_wvalid(o_lpddr_ppp_0_targ_mt_axi_m_wvalid),
    .o_lpddr_ppp_0_targ_syscfg_apb_m_paddr(o_lpddr_ppp_0_targ_syscfg_apb_m_paddr),
    .o_lpddr_ppp_0_targ_syscfg_apb_m_penable(o_lpddr_ppp_0_targ_syscfg_apb_m_penable),
    .o_lpddr_ppp_0_targ_syscfg_apb_m_pprot(o_lpddr_ppp_0_targ_syscfg_apb_m_pprot),
    .i_lpddr_ppp_0_targ_syscfg_apb_m_prdata(i_lpddr_ppp_0_targ_syscfg_apb_m_prdata),
    .i_lpddr_ppp_0_targ_syscfg_apb_m_pready(i_lpddr_ppp_0_targ_syscfg_apb_m_pready),
    .o_lpddr_ppp_0_targ_syscfg_apb_m_psel(o_lpddr_ppp_0_targ_syscfg_apb_m_psel),
    .i_lpddr_ppp_0_targ_syscfg_apb_m_pslverr(i_lpddr_ppp_0_targ_syscfg_apb_m_pslverr),
    .o_lpddr_ppp_0_targ_syscfg_apb_m_pstrb(o_lpddr_ppp_0_targ_syscfg_apb_m_pstrb),
    .o_lpddr_ppp_0_targ_syscfg_apb_m_pwdata(o_lpddr_ppp_0_targ_syscfg_apb_m_pwdata),
    .o_lpddr_ppp_0_targ_syscfg_apb_m_pwrite(o_lpddr_ppp_0_targ_syscfg_apb_m_pwrite),
    .i_lpddr_ppp_1_aon_clk(i_lpddr_ppp_1_aon_clk),
    .i_lpddr_ppp_1_aon_rst_n(lpddr_ppp_1_aon_rst_n_synced),
    .o_lpddr_ppp_1_cfg_pwr_idle_val(o_lpddr_ppp_1_cfg_pwr_idle_val),
    .o_lpddr_ppp_1_cfg_pwr_idle_ack(o_lpddr_ppp_1_cfg_pwr_idle_ack),
    .i_lpddr_ppp_1_cfg_pwr_idle_req(i_lpddr_ppp_1_cfg_pwr_idle_req),
    .i_lpddr_ppp_1_clk(i_lpddr_ppp_1_clk),
    .i_lpddr_ppp_1_clken(i_lpddr_ppp_1_clken),
    .o_lpddr_ppp_1_pwr_idle_val(o_lpddr_ppp_1_pwr_idle_val),
    .o_lpddr_ppp_1_pwr_idle_ack(o_lpddr_ppp_1_pwr_idle_ack),
    .i_lpddr_ppp_1_pwr_idle_req(i_lpddr_ppp_1_pwr_idle_req),
    .i_lpddr_ppp_1_rst_n(i_lpddr_ppp_1_rst_n),
    .o_lpddr_ppp_1_targ_cfg_apb_m_paddr(o_lpddr_ppp_1_targ_cfg_apb_m_paddr),
    .o_lpddr_ppp_1_targ_cfg_apb_m_penable(o_lpddr_ppp_1_targ_cfg_apb_m_penable),
    .o_lpddr_ppp_1_targ_cfg_apb_m_pprot(o_lpddr_ppp_1_targ_cfg_apb_m_pprot),
    .i_lpddr_ppp_1_targ_cfg_apb_m_prdata(i_lpddr_ppp_1_targ_cfg_apb_m_prdata),
    .i_lpddr_ppp_1_targ_cfg_apb_m_pready(i_lpddr_ppp_1_targ_cfg_apb_m_pready),
    .o_lpddr_ppp_1_targ_cfg_apb_m_psel(o_lpddr_ppp_1_targ_cfg_apb_m_psel),
    .i_lpddr_ppp_1_targ_cfg_apb_m_pslverr(i_lpddr_ppp_1_targ_cfg_apb_m_pslverr),
    .o_lpddr_ppp_1_targ_cfg_apb_m_pstrb(o_lpddr_ppp_1_targ_cfg_apb_m_pstrb),
    .o_lpddr_ppp_1_targ_cfg_apb_m_pwdata(o_lpddr_ppp_1_targ_cfg_apb_m_pwdata),
    .o_lpddr_ppp_1_targ_cfg_apb_m_pwrite(o_lpddr_ppp_1_targ_cfg_apb_m_pwrite),
    .o_lpddr_ppp_1_targ_mt_axi_m_araddr(o_lpddr_ppp_1_targ_mt_axi_m_araddr),
    .o_lpddr_ppp_1_targ_mt_axi_m_arburst(o_lpddr_ppp_1_targ_mt_axi_m_arburst),
    .o_lpddr_ppp_1_targ_mt_axi_m_arcache(o_lpddr_ppp_1_targ_mt_axi_m_arcache),
    .o_lpddr_ppp_1_targ_mt_axi_m_arid(o_lpddr_ppp_1_targ_mt_axi_m_arid),
    .o_lpddr_ppp_1_targ_mt_axi_m_arlen(o_lpddr_ppp_1_targ_mt_axi_m_arlen),
    .o_lpddr_ppp_1_targ_mt_axi_m_arlock(o_lpddr_ppp_1_targ_mt_axi_m_arlock),
    .o_lpddr_ppp_1_targ_mt_axi_m_arprot(o_lpddr_ppp_1_targ_mt_axi_m_arprot),
    .o_lpddr_ppp_1_targ_mt_axi_m_arqos(o_lpddr_ppp_1_targ_mt_axi_m_arqos),
    .i_lpddr_ppp_1_targ_mt_axi_m_arready(i_lpddr_ppp_1_targ_mt_axi_m_arready),
    .o_lpddr_ppp_1_targ_mt_axi_m_arsize(o_lpddr_ppp_1_targ_mt_axi_m_arsize),
    .o_lpddr_ppp_1_targ_mt_axi_m_arvalid(o_lpddr_ppp_1_targ_mt_axi_m_arvalid),
    .o_lpddr_ppp_1_targ_mt_axi_m_awaddr(o_lpddr_ppp_1_targ_mt_axi_m_awaddr),
    .o_lpddr_ppp_1_targ_mt_axi_m_awburst(o_lpddr_ppp_1_targ_mt_axi_m_awburst),
    .o_lpddr_ppp_1_targ_mt_axi_m_awcache(o_lpddr_ppp_1_targ_mt_axi_m_awcache),
    .o_lpddr_ppp_1_targ_mt_axi_m_awid(o_lpddr_ppp_1_targ_mt_axi_m_awid),
    .o_lpddr_ppp_1_targ_mt_axi_m_awlen(o_lpddr_ppp_1_targ_mt_axi_m_awlen),
    .o_lpddr_ppp_1_targ_mt_axi_m_awlock(o_lpddr_ppp_1_targ_mt_axi_m_awlock),
    .o_lpddr_ppp_1_targ_mt_axi_m_awprot(o_lpddr_ppp_1_targ_mt_axi_m_awprot),
    .o_lpddr_ppp_1_targ_mt_axi_m_awqos(o_lpddr_ppp_1_targ_mt_axi_m_awqos),
    .i_lpddr_ppp_1_targ_mt_axi_m_awready(i_lpddr_ppp_1_targ_mt_axi_m_awready),
    .o_lpddr_ppp_1_targ_mt_axi_m_awsize(o_lpddr_ppp_1_targ_mt_axi_m_awsize),
    .o_lpddr_ppp_1_targ_mt_axi_m_awvalid(o_lpddr_ppp_1_targ_mt_axi_m_awvalid),
    .i_lpddr_ppp_1_targ_mt_axi_m_bid(i_lpddr_ppp_1_targ_mt_axi_m_bid),
    .o_lpddr_ppp_1_targ_mt_axi_m_bready(o_lpddr_ppp_1_targ_mt_axi_m_bready),
    .i_lpddr_ppp_1_targ_mt_axi_m_bresp(i_lpddr_ppp_1_targ_mt_axi_m_bresp),
    .i_lpddr_ppp_1_targ_mt_axi_m_bvalid(i_lpddr_ppp_1_targ_mt_axi_m_bvalid),
    .i_lpddr_ppp_1_targ_mt_axi_m_rdata(i_lpddr_ppp_1_targ_mt_axi_m_rdata),
    .i_lpddr_ppp_1_targ_mt_axi_m_rid(i_lpddr_ppp_1_targ_mt_axi_m_rid),
    .i_lpddr_ppp_1_targ_mt_axi_m_rlast(i_lpddr_ppp_1_targ_mt_axi_m_rlast),
    .o_lpddr_ppp_1_targ_mt_axi_m_rready(o_lpddr_ppp_1_targ_mt_axi_m_rready),
    .i_lpddr_ppp_1_targ_mt_axi_m_rresp(i_lpddr_ppp_1_targ_mt_axi_m_rresp),
    .i_lpddr_ppp_1_targ_mt_axi_m_rvalid(i_lpddr_ppp_1_targ_mt_axi_m_rvalid),
    .o_lpddr_ppp_1_targ_mt_axi_m_wdata(o_lpddr_ppp_1_targ_mt_axi_m_wdata),
    .o_lpddr_ppp_1_targ_mt_axi_m_wlast(o_lpddr_ppp_1_targ_mt_axi_m_wlast),
    .i_lpddr_ppp_1_targ_mt_axi_m_wready(i_lpddr_ppp_1_targ_mt_axi_m_wready),
    .o_lpddr_ppp_1_targ_mt_axi_m_wstrb(o_lpddr_ppp_1_targ_mt_axi_m_wstrb),
    .o_lpddr_ppp_1_targ_mt_axi_m_wvalid(o_lpddr_ppp_1_targ_mt_axi_m_wvalid),
    .o_lpddr_ppp_1_targ_syscfg_apb_m_paddr(o_lpddr_ppp_1_targ_syscfg_apb_m_paddr),
    .o_lpddr_ppp_1_targ_syscfg_apb_m_penable(o_lpddr_ppp_1_targ_syscfg_apb_m_penable),
    .o_lpddr_ppp_1_targ_syscfg_apb_m_pprot(o_lpddr_ppp_1_targ_syscfg_apb_m_pprot),
    .i_lpddr_ppp_1_targ_syscfg_apb_m_prdata(i_lpddr_ppp_1_targ_syscfg_apb_m_prdata),
    .i_lpddr_ppp_1_targ_syscfg_apb_m_pready(i_lpddr_ppp_1_targ_syscfg_apb_m_pready),
    .o_lpddr_ppp_1_targ_syscfg_apb_m_psel(o_lpddr_ppp_1_targ_syscfg_apb_m_psel),
    .i_lpddr_ppp_1_targ_syscfg_apb_m_pslverr(i_lpddr_ppp_1_targ_syscfg_apb_m_pslverr),
    .o_lpddr_ppp_1_targ_syscfg_apb_m_pstrb(o_lpddr_ppp_1_targ_syscfg_apb_m_pstrb),
    .o_lpddr_ppp_1_targ_syscfg_apb_m_pwdata(o_lpddr_ppp_1_targ_syscfg_apb_m_pwdata),
    .o_lpddr_ppp_1_targ_syscfg_apb_m_pwrite(o_lpddr_ppp_1_targ_syscfg_apb_m_pwrite),
    .i_lpddr_ppp_2_aon_clk(i_lpddr_ppp_2_aon_clk),
    .i_lpddr_ppp_2_aon_rst_n(lpddr_ppp_2_aon_rst_n_synced),
    .o_lpddr_ppp_2_cfg_pwr_idle_val(o_lpddr_ppp_2_cfg_pwr_idle_val),
    .o_lpddr_ppp_2_cfg_pwr_idle_ack(o_lpddr_ppp_2_cfg_pwr_idle_ack),
    .i_lpddr_ppp_2_cfg_pwr_idle_req(i_lpddr_ppp_2_cfg_pwr_idle_req),
    .i_lpddr_ppp_2_clk(i_lpddr_ppp_2_clk),
    .i_lpddr_ppp_2_clken(i_lpddr_ppp_2_clken),
    .o_lpddr_ppp_2_pwr_idle_val(o_lpddr_ppp_2_pwr_idle_val),
    .o_lpddr_ppp_2_pwr_idle_ack(o_lpddr_ppp_2_pwr_idle_ack),
    .i_lpddr_ppp_2_pwr_idle_req(i_lpddr_ppp_2_pwr_idle_req),
    .i_lpddr_ppp_2_rst_n(i_lpddr_ppp_2_rst_n),
    .o_lpddr_ppp_2_targ_cfg_apb_m_paddr(o_lpddr_ppp_2_targ_cfg_apb_m_paddr),
    .o_lpddr_ppp_2_targ_cfg_apb_m_penable(o_lpddr_ppp_2_targ_cfg_apb_m_penable),
    .o_lpddr_ppp_2_targ_cfg_apb_m_pprot(o_lpddr_ppp_2_targ_cfg_apb_m_pprot),
    .i_lpddr_ppp_2_targ_cfg_apb_m_prdata(i_lpddr_ppp_2_targ_cfg_apb_m_prdata),
    .i_lpddr_ppp_2_targ_cfg_apb_m_pready(i_lpddr_ppp_2_targ_cfg_apb_m_pready),
    .o_lpddr_ppp_2_targ_cfg_apb_m_psel(o_lpddr_ppp_2_targ_cfg_apb_m_psel),
    .i_lpddr_ppp_2_targ_cfg_apb_m_pslverr(i_lpddr_ppp_2_targ_cfg_apb_m_pslverr),
    .o_lpddr_ppp_2_targ_cfg_apb_m_pstrb(o_lpddr_ppp_2_targ_cfg_apb_m_pstrb),
    .o_lpddr_ppp_2_targ_cfg_apb_m_pwdata(o_lpddr_ppp_2_targ_cfg_apb_m_pwdata),
    .o_lpddr_ppp_2_targ_cfg_apb_m_pwrite(o_lpddr_ppp_2_targ_cfg_apb_m_pwrite),
    .o_lpddr_ppp_2_targ_mt_axi_m_araddr(o_lpddr_ppp_2_targ_mt_axi_m_araddr),
    .o_lpddr_ppp_2_targ_mt_axi_m_arburst(o_lpddr_ppp_2_targ_mt_axi_m_arburst),
    .o_lpddr_ppp_2_targ_mt_axi_m_arcache(o_lpddr_ppp_2_targ_mt_axi_m_arcache),
    .o_lpddr_ppp_2_targ_mt_axi_m_arid(o_lpddr_ppp_2_targ_mt_axi_m_arid),
    .o_lpddr_ppp_2_targ_mt_axi_m_arlen(o_lpddr_ppp_2_targ_mt_axi_m_arlen),
    .o_lpddr_ppp_2_targ_mt_axi_m_arlock(o_lpddr_ppp_2_targ_mt_axi_m_arlock),
    .o_lpddr_ppp_2_targ_mt_axi_m_arprot(o_lpddr_ppp_2_targ_mt_axi_m_arprot),
    .o_lpddr_ppp_2_targ_mt_axi_m_arqos(o_lpddr_ppp_2_targ_mt_axi_m_arqos),
    .i_lpddr_ppp_2_targ_mt_axi_m_arready(i_lpddr_ppp_2_targ_mt_axi_m_arready),
    .o_lpddr_ppp_2_targ_mt_axi_m_arsize(o_lpddr_ppp_2_targ_mt_axi_m_arsize),
    .o_lpddr_ppp_2_targ_mt_axi_m_arvalid(o_lpddr_ppp_2_targ_mt_axi_m_arvalid),
    .o_lpddr_ppp_2_targ_mt_axi_m_awaddr(o_lpddr_ppp_2_targ_mt_axi_m_awaddr),
    .o_lpddr_ppp_2_targ_mt_axi_m_awburst(o_lpddr_ppp_2_targ_mt_axi_m_awburst),
    .o_lpddr_ppp_2_targ_mt_axi_m_awcache(o_lpddr_ppp_2_targ_mt_axi_m_awcache),
    .o_lpddr_ppp_2_targ_mt_axi_m_awid(o_lpddr_ppp_2_targ_mt_axi_m_awid),
    .o_lpddr_ppp_2_targ_mt_axi_m_awlen(o_lpddr_ppp_2_targ_mt_axi_m_awlen),
    .o_lpddr_ppp_2_targ_mt_axi_m_awlock(o_lpddr_ppp_2_targ_mt_axi_m_awlock),
    .o_lpddr_ppp_2_targ_mt_axi_m_awprot(o_lpddr_ppp_2_targ_mt_axi_m_awprot),
    .o_lpddr_ppp_2_targ_mt_axi_m_awqos(o_lpddr_ppp_2_targ_mt_axi_m_awqos),
    .i_lpddr_ppp_2_targ_mt_axi_m_awready(i_lpddr_ppp_2_targ_mt_axi_m_awready),
    .o_lpddr_ppp_2_targ_mt_axi_m_awsize(o_lpddr_ppp_2_targ_mt_axi_m_awsize),
    .o_lpddr_ppp_2_targ_mt_axi_m_awvalid(o_lpddr_ppp_2_targ_mt_axi_m_awvalid),
    .i_lpddr_ppp_2_targ_mt_axi_m_bid(i_lpddr_ppp_2_targ_mt_axi_m_bid),
    .o_lpddr_ppp_2_targ_mt_axi_m_bready(o_lpddr_ppp_2_targ_mt_axi_m_bready),
    .i_lpddr_ppp_2_targ_mt_axi_m_bresp(i_lpddr_ppp_2_targ_mt_axi_m_bresp),
    .i_lpddr_ppp_2_targ_mt_axi_m_bvalid(i_lpddr_ppp_2_targ_mt_axi_m_bvalid),
    .i_lpddr_ppp_2_targ_mt_axi_m_rdata(i_lpddr_ppp_2_targ_mt_axi_m_rdata),
    .i_lpddr_ppp_2_targ_mt_axi_m_rid(i_lpddr_ppp_2_targ_mt_axi_m_rid),
    .i_lpddr_ppp_2_targ_mt_axi_m_rlast(i_lpddr_ppp_2_targ_mt_axi_m_rlast),
    .o_lpddr_ppp_2_targ_mt_axi_m_rready(o_lpddr_ppp_2_targ_mt_axi_m_rready),
    .i_lpddr_ppp_2_targ_mt_axi_m_rresp(i_lpddr_ppp_2_targ_mt_axi_m_rresp),
    .i_lpddr_ppp_2_targ_mt_axi_m_rvalid(i_lpddr_ppp_2_targ_mt_axi_m_rvalid),
    .o_lpddr_ppp_2_targ_mt_axi_m_wdata(o_lpddr_ppp_2_targ_mt_axi_m_wdata),
    .o_lpddr_ppp_2_targ_mt_axi_m_wlast(o_lpddr_ppp_2_targ_mt_axi_m_wlast),
    .i_lpddr_ppp_2_targ_mt_axi_m_wready(i_lpddr_ppp_2_targ_mt_axi_m_wready),
    .o_lpddr_ppp_2_targ_mt_axi_m_wstrb(o_lpddr_ppp_2_targ_mt_axi_m_wstrb),
    .o_lpddr_ppp_2_targ_mt_axi_m_wvalid(o_lpddr_ppp_2_targ_mt_axi_m_wvalid),
    .o_lpddr_ppp_2_targ_syscfg_apb_m_paddr(o_lpddr_ppp_2_targ_syscfg_apb_m_paddr),
    .o_lpddr_ppp_2_targ_syscfg_apb_m_penable(o_lpddr_ppp_2_targ_syscfg_apb_m_penable),
    .o_lpddr_ppp_2_targ_syscfg_apb_m_pprot(o_lpddr_ppp_2_targ_syscfg_apb_m_pprot),
    .i_lpddr_ppp_2_targ_syscfg_apb_m_prdata(i_lpddr_ppp_2_targ_syscfg_apb_m_prdata),
    .i_lpddr_ppp_2_targ_syscfg_apb_m_pready(i_lpddr_ppp_2_targ_syscfg_apb_m_pready),
    .o_lpddr_ppp_2_targ_syscfg_apb_m_psel(o_lpddr_ppp_2_targ_syscfg_apb_m_psel),
    .i_lpddr_ppp_2_targ_syscfg_apb_m_pslverr(i_lpddr_ppp_2_targ_syscfg_apb_m_pslverr),
    .o_lpddr_ppp_2_targ_syscfg_apb_m_pstrb(o_lpddr_ppp_2_targ_syscfg_apb_m_pstrb),
    .o_lpddr_ppp_2_targ_syscfg_apb_m_pwdata(o_lpddr_ppp_2_targ_syscfg_apb_m_pwdata),
    .o_lpddr_ppp_2_targ_syscfg_apb_m_pwrite(o_lpddr_ppp_2_targ_syscfg_apb_m_pwrite),
    .i_lpddr_ppp_3_aon_clk(i_lpddr_ppp_3_aon_clk),
    .i_lpddr_ppp_3_aon_rst_n(lpddr_ppp_3_aon_rst_n_synced),
    .o_lpddr_ppp_3_cfg_pwr_idle_val(o_lpddr_ppp_3_cfg_pwr_idle_val),
    .o_lpddr_ppp_3_cfg_pwr_idle_ack(o_lpddr_ppp_3_cfg_pwr_idle_ack),
    .i_lpddr_ppp_3_cfg_pwr_idle_req(i_lpddr_ppp_3_cfg_pwr_idle_req),
    .i_lpddr_ppp_3_clk(i_lpddr_ppp_3_clk),
    .i_lpddr_ppp_3_clken(i_lpddr_ppp_3_clken),
    .o_lpddr_ppp_3_pwr_idle_val(o_lpddr_ppp_3_pwr_idle_val),
    .o_lpddr_ppp_3_pwr_idle_ack(o_lpddr_ppp_3_pwr_idle_ack),
    .i_lpddr_ppp_3_pwr_idle_req(i_lpddr_ppp_3_pwr_idle_req),
    .i_lpddr_ppp_3_rst_n(i_lpddr_ppp_3_rst_n),
    .o_lpddr_ppp_3_targ_cfg_apb_m_paddr(o_lpddr_ppp_3_targ_cfg_apb_m_paddr),
    .o_lpddr_ppp_3_targ_cfg_apb_m_penable(o_lpddr_ppp_3_targ_cfg_apb_m_penable),
    .o_lpddr_ppp_3_targ_cfg_apb_m_pprot(o_lpddr_ppp_3_targ_cfg_apb_m_pprot),
    .i_lpddr_ppp_3_targ_cfg_apb_m_prdata(i_lpddr_ppp_3_targ_cfg_apb_m_prdata),
    .i_lpddr_ppp_3_targ_cfg_apb_m_pready(i_lpddr_ppp_3_targ_cfg_apb_m_pready),
    .o_lpddr_ppp_3_targ_cfg_apb_m_psel(o_lpddr_ppp_3_targ_cfg_apb_m_psel),
    .i_lpddr_ppp_3_targ_cfg_apb_m_pslverr(i_lpddr_ppp_3_targ_cfg_apb_m_pslverr),
    .o_lpddr_ppp_3_targ_cfg_apb_m_pstrb(o_lpddr_ppp_3_targ_cfg_apb_m_pstrb),
    .o_lpddr_ppp_3_targ_cfg_apb_m_pwdata(o_lpddr_ppp_3_targ_cfg_apb_m_pwdata),
    .o_lpddr_ppp_3_targ_cfg_apb_m_pwrite(o_lpddr_ppp_3_targ_cfg_apb_m_pwrite),
    .o_lpddr_ppp_3_targ_mt_axi_m_araddr(o_lpddr_ppp_3_targ_mt_axi_m_araddr),
    .o_lpddr_ppp_3_targ_mt_axi_m_arburst(o_lpddr_ppp_3_targ_mt_axi_m_arburst),
    .o_lpddr_ppp_3_targ_mt_axi_m_arcache(o_lpddr_ppp_3_targ_mt_axi_m_arcache),
    .o_lpddr_ppp_3_targ_mt_axi_m_arid(o_lpddr_ppp_3_targ_mt_axi_m_arid),
    .o_lpddr_ppp_3_targ_mt_axi_m_arlen(o_lpddr_ppp_3_targ_mt_axi_m_arlen),
    .o_lpddr_ppp_3_targ_mt_axi_m_arlock(o_lpddr_ppp_3_targ_mt_axi_m_arlock),
    .o_lpddr_ppp_3_targ_mt_axi_m_arprot(o_lpddr_ppp_3_targ_mt_axi_m_arprot),
    .o_lpddr_ppp_3_targ_mt_axi_m_arqos(o_lpddr_ppp_3_targ_mt_axi_m_arqos),
    .i_lpddr_ppp_3_targ_mt_axi_m_arready(i_lpddr_ppp_3_targ_mt_axi_m_arready),
    .o_lpddr_ppp_3_targ_mt_axi_m_arsize(o_lpddr_ppp_3_targ_mt_axi_m_arsize),
    .o_lpddr_ppp_3_targ_mt_axi_m_arvalid(o_lpddr_ppp_3_targ_mt_axi_m_arvalid),
    .o_lpddr_ppp_3_targ_mt_axi_m_awaddr(o_lpddr_ppp_3_targ_mt_axi_m_awaddr),
    .o_lpddr_ppp_3_targ_mt_axi_m_awburst(o_lpddr_ppp_3_targ_mt_axi_m_awburst),
    .o_lpddr_ppp_3_targ_mt_axi_m_awcache(o_lpddr_ppp_3_targ_mt_axi_m_awcache),
    .o_lpddr_ppp_3_targ_mt_axi_m_awid(o_lpddr_ppp_3_targ_mt_axi_m_awid),
    .o_lpddr_ppp_3_targ_mt_axi_m_awlen(o_lpddr_ppp_3_targ_mt_axi_m_awlen),
    .o_lpddr_ppp_3_targ_mt_axi_m_awlock(o_lpddr_ppp_3_targ_mt_axi_m_awlock),
    .o_lpddr_ppp_3_targ_mt_axi_m_awprot(o_lpddr_ppp_3_targ_mt_axi_m_awprot),
    .o_lpddr_ppp_3_targ_mt_axi_m_awqos(o_lpddr_ppp_3_targ_mt_axi_m_awqos),
    .i_lpddr_ppp_3_targ_mt_axi_m_awready(i_lpddr_ppp_3_targ_mt_axi_m_awready),
    .o_lpddr_ppp_3_targ_mt_axi_m_awsize(o_lpddr_ppp_3_targ_mt_axi_m_awsize),
    .o_lpddr_ppp_3_targ_mt_axi_m_awvalid(o_lpddr_ppp_3_targ_mt_axi_m_awvalid),
    .i_lpddr_ppp_3_targ_mt_axi_m_bid(i_lpddr_ppp_3_targ_mt_axi_m_bid),
    .o_lpddr_ppp_3_targ_mt_axi_m_bready(o_lpddr_ppp_3_targ_mt_axi_m_bready),
    .i_lpddr_ppp_3_targ_mt_axi_m_bresp(i_lpddr_ppp_3_targ_mt_axi_m_bresp),
    .i_lpddr_ppp_3_targ_mt_axi_m_bvalid(i_lpddr_ppp_3_targ_mt_axi_m_bvalid),
    .i_lpddr_ppp_3_targ_mt_axi_m_rdata(i_lpddr_ppp_3_targ_mt_axi_m_rdata),
    .i_lpddr_ppp_3_targ_mt_axi_m_rid(i_lpddr_ppp_3_targ_mt_axi_m_rid),
    .i_lpddr_ppp_3_targ_mt_axi_m_rlast(i_lpddr_ppp_3_targ_mt_axi_m_rlast),
    .o_lpddr_ppp_3_targ_mt_axi_m_rready(o_lpddr_ppp_3_targ_mt_axi_m_rready),
    .i_lpddr_ppp_3_targ_mt_axi_m_rresp(i_lpddr_ppp_3_targ_mt_axi_m_rresp),
    .i_lpddr_ppp_3_targ_mt_axi_m_rvalid(i_lpddr_ppp_3_targ_mt_axi_m_rvalid),
    .o_lpddr_ppp_3_targ_mt_axi_m_wdata(o_lpddr_ppp_3_targ_mt_axi_m_wdata),
    .o_lpddr_ppp_3_targ_mt_axi_m_wlast(o_lpddr_ppp_3_targ_mt_axi_m_wlast),
    .i_lpddr_ppp_3_targ_mt_axi_m_wready(i_lpddr_ppp_3_targ_mt_axi_m_wready),
    .o_lpddr_ppp_3_targ_mt_axi_m_wstrb(o_lpddr_ppp_3_targ_mt_axi_m_wstrb),
    .o_lpddr_ppp_3_targ_mt_axi_m_wvalid(o_lpddr_ppp_3_targ_mt_axi_m_wvalid),
    .o_lpddr_ppp_3_targ_syscfg_apb_m_paddr(o_lpddr_ppp_3_targ_syscfg_apb_m_paddr),
    .o_lpddr_ppp_3_targ_syscfg_apb_m_penable(o_lpddr_ppp_3_targ_syscfg_apb_m_penable),
    .o_lpddr_ppp_3_targ_syscfg_apb_m_pprot(o_lpddr_ppp_3_targ_syscfg_apb_m_pprot),
    .i_lpddr_ppp_3_targ_syscfg_apb_m_prdata(i_lpddr_ppp_3_targ_syscfg_apb_m_prdata),
    .i_lpddr_ppp_3_targ_syscfg_apb_m_pready(i_lpddr_ppp_3_targ_syscfg_apb_m_pready),
    .o_lpddr_ppp_3_targ_syscfg_apb_m_psel(o_lpddr_ppp_3_targ_syscfg_apb_m_psel),
    .i_lpddr_ppp_3_targ_syscfg_apb_m_pslverr(i_lpddr_ppp_3_targ_syscfg_apb_m_pslverr),
    .o_lpddr_ppp_3_targ_syscfg_apb_m_pstrb(o_lpddr_ppp_3_targ_syscfg_apb_m_pstrb),
    .o_lpddr_ppp_3_targ_syscfg_apb_m_pwdata(o_lpddr_ppp_3_targ_syscfg_apb_m_pwdata),
    .o_lpddr_ppp_3_targ_syscfg_apb_m_pwrite(o_lpddr_ppp_3_targ_syscfg_apb_m_pwrite),
    .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .i_noc_clk(i_noc_clk),
    .i_noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en),
    .i_soc_periph_aon_clk(i_soc_periph_aon_clk),
    .i_soc_periph_aon_rst_n(soc_periph_aon_rst_n_synced),
    .i_soc_periph_clk(i_soc_periph_clk),
    .i_soc_periph_clken(i_soc_periph_clken),
    .i_soc_periph_init_lt_axi_s_araddr(i_soc_periph_init_lt_axi_s_araddr),
    .i_soc_periph_init_lt_axi_s_arburst(i_soc_periph_init_lt_axi_s_arburst),
    .i_soc_periph_init_lt_axi_s_arcache(i_soc_periph_init_lt_axi_s_arcache),
    .i_soc_periph_init_lt_axi_s_arid(i_soc_periph_init_lt_axi_s_arid),
    .i_soc_periph_init_lt_axi_s_arlen(i_soc_periph_init_lt_axi_s_arlen),
    .i_soc_periph_init_lt_axi_s_arlock(i_soc_periph_init_lt_axi_s_arlock),
    .i_soc_periph_init_lt_axi_s_arprot(i_soc_periph_init_lt_axi_s_arprot),
    .i_soc_periph_init_lt_axi_s_arqos(i_soc_periph_init_lt_axi_s_arqos),
    .o_soc_periph_init_lt_axi_s_arready(o_soc_periph_init_lt_axi_s_arready),
    .i_soc_periph_init_lt_axi_s_arsize(i_soc_periph_init_lt_axi_s_arsize),
    .i_soc_periph_init_lt_axi_s_arvalid(i_soc_periph_init_lt_axi_s_arvalid),
    .i_soc_periph_init_lt_axi_s_awaddr(i_soc_periph_init_lt_axi_s_awaddr),
    .i_soc_periph_init_lt_axi_s_awburst(i_soc_periph_init_lt_axi_s_awburst),
    .i_soc_periph_init_lt_axi_s_awcache(i_soc_periph_init_lt_axi_s_awcache),
    .i_soc_periph_init_lt_axi_s_awid(i_soc_periph_init_lt_axi_s_awid),
    .i_soc_periph_init_lt_axi_s_awlen(i_soc_periph_init_lt_axi_s_awlen),
    .i_soc_periph_init_lt_axi_s_awlock(i_soc_periph_init_lt_axi_s_awlock),
    .i_soc_periph_init_lt_axi_s_awprot(i_soc_periph_init_lt_axi_s_awprot),
    .i_soc_periph_init_lt_axi_s_awqos(i_soc_periph_init_lt_axi_s_awqos),
    .o_soc_periph_init_lt_axi_s_awready(o_soc_periph_init_lt_axi_s_awready),
    .i_soc_periph_init_lt_axi_s_awsize(i_soc_periph_init_lt_axi_s_awsize),
    .i_soc_periph_init_lt_axi_s_awvalid(i_soc_periph_init_lt_axi_s_awvalid),
    .o_soc_periph_init_lt_axi_s_bid(o_soc_periph_init_lt_axi_s_bid),
    .i_soc_periph_init_lt_axi_s_bready(i_soc_periph_init_lt_axi_s_bready),
    .o_soc_periph_init_lt_axi_s_bresp(o_soc_periph_init_lt_axi_s_bresp),
    .o_soc_periph_init_lt_axi_s_bvalid(o_soc_periph_init_lt_axi_s_bvalid),
    .o_soc_periph_init_lt_axi_s_rdata(o_soc_periph_init_lt_axi_s_rdata),
    .o_soc_periph_init_lt_axi_s_rid(o_soc_periph_init_lt_axi_s_rid),
    .o_soc_periph_init_lt_axi_s_rlast(o_soc_periph_init_lt_axi_s_rlast),
    .i_soc_periph_init_lt_axi_s_rready(i_soc_periph_init_lt_axi_s_rready),
    .o_soc_periph_init_lt_axi_s_rresp(o_soc_periph_init_lt_axi_s_rresp),
    .o_soc_periph_init_lt_axi_s_rvalid(o_soc_periph_init_lt_axi_s_rvalid),
    .i_soc_periph_init_lt_axi_s_wdata(i_soc_periph_init_lt_axi_s_wdata),
    .i_soc_periph_init_lt_axi_s_wlast(i_soc_periph_init_lt_axi_s_wlast),
    .o_soc_periph_init_lt_axi_s_wready(o_soc_periph_init_lt_axi_s_wready),
    .i_soc_periph_init_lt_axi_s_wstrb(i_soc_periph_init_lt_axi_s_wstrb),
    .i_soc_periph_init_lt_axi_s_wvalid(i_soc_periph_init_lt_axi_s_wvalid),
    .o_soc_periph_pwr_idle_val(o_soc_periph_pwr_idle_val),
    .o_soc_periph_pwr_idle_ack(o_soc_periph_pwr_idle_ack),
    .i_soc_periph_pwr_idle_req(i_soc_periph_pwr_idle_req),
    .i_soc_periph_rst_n(i_soc_periph_rst_n),
    .o_soc_periph_targ_lt_axi_m_araddr(o_soc_periph_targ_lt_axi_m_araddr),
    .o_soc_periph_targ_lt_axi_m_arburst(o_soc_periph_targ_lt_axi_m_arburst),
    .o_soc_periph_targ_lt_axi_m_arcache(o_soc_periph_targ_lt_axi_m_arcache),
    .o_soc_periph_targ_lt_axi_m_arid(o_soc_periph_targ_lt_axi_m_arid),
    .o_soc_periph_targ_lt_axi_m_arlen(o_soc_periph_targ_lt_axi_m_arlen),
    .o_soc_periph_targ_lt_axi_m_arlock(o_soc_periph_targ_lt_axi_m_arlock),
    .o_soc_periph_targ_lt_axi_m_arprot(o_soc_periph_targ_lt_axi_m_arprot),
    .o_soc_periph_targ_lt_axi_m_arqos(o_soc_periph_targ_lt_axi_m_arqos),
    .i_soc_periph_targ_lt_axi_m_arready(i_soc_periph_targ_lt_axi_m_arready),
    .o_soc_periph_targ_lt_axi_m_arsize(o_soc_periph_targ_lt_axi_m_arsize),
    .o_soc_periph_targ_lt_axi_m_arvalid(o_soc_periph_targ_lt_axi_m_arvalid),
    .o_soc_periph_targ_lt_axi_m_awaddr(o_soc_periph_targ_lt_axi_m_awaddr),
    .o_soc_periph_targ_lt_axi_m_awburst(o_soc_periph_targ_lt_axi_m_awburst),
    .o_soc_periph_targ_lt_axi_m_awcache(o_soc_periph_targ_lt_axi_m_awcache),
    .o_soc_periph_targ_lt_axi_m_awid(o_soc_periph_targ_lt_axi_m_awid),
    .o_soc_periph_targ_lt_axi_m_awlen(o_soc_periph_targ_lt_axi_m_awlen),
    .o_soc_periph_targ_lt_axi_m_awlock(o_soc_periph_targ_lt_axi_m_awlock),
    .o_soc_periph_targ_lt_axi_m_awprot(o_soc_periph_targ_lt_axi_m_awprot),
    .o_soc_periph_targ_lt_axi_m_awqos(o_soc_periph_targ_lt_axi_m_awqos),
    .i_soc_periph_targ_lt_axi_m_awready(i_soc_periph_targ_lt_axi_m_awready),
    .o_soc_periph_targ_lt_axi_m_awsize(o_soc_periph_targ_lt_axi_m_awsize),
    .o_soc_periph_targ_lt_axi_m_awvalid(o_soc_periph_targ_lt_axi_m_awvalid),
    .i_soc_periph_targ_lt_axi_m_bid(i_soc_periph_targ_lt_axi_m_bid),
    .o_soc_periph_targ_lt_axi_m_bready(o_soc_periph_targ_lt_axi_m_bready),
    .i_soc_periph_targ_lt_axi_m_bresp(i_soc_periph_targ_lt_axi_m_bresp),
    .i_soc_periph_targ_lt_axi_m_bvalid(i_soc_periph_targ_lt_axi_m_bvalid),
    .i_soc_periph_targ_lt_axi_m_rdata(i_soc_periph_targ_lt_axi_m_rdata),
    .i_soc_periph_targ_lt_axi_m_rid(i_soc_periph_targ_lt_axi_m_rid),
    .i_soc_periph_targ_lt_axi_m_rlast(i_soc_periph_targ_lt_axi_m_rlast),
    .o_soc_periph_targ_lt_axi_m_rready(o_soc_periph_targ_lt_axi_m_rready),
    .i_soc_periph_targ_lt_axi_m_rresp(i_soc_periph_targ_lt_axi_m_rresp),
    .i_soc_periph_targ_lt_axi_m_rvalid(i_soc_periph_targ_lt_axi_m_rvalid),
    .o_soc_periph_targ_lt_axi_m_wdata(o_soc_periph_targ_lt_axi_m_wdata),
    .o_soc_periph_targ_lt_axi_m_wlast(o_soc_periph_targ_lt_axi_m_wlast),
    .i_soc_periph_targ_lt_axi_m_wready(i_soc_periph_targ_lt_axi_m_wready),
    .o_soc_periph_targ_lt_axi_m_wstrb(o_soc_periph_targ_lt_axi_m_wstrb),
    .o_soc_periph_targ_lt_axi_m_wvalid(o_soc_periph_targ_lt_axi_m_wvalid),
    .o_soc_periph_targ_syscfg_apb_m_paddr(o_soc_periph_targ_syscfg_apb_m_paddr),
    .o_soc_periph_targ_syscfg_apb_m_penable(o_soc_periph_targ_syscfg_apb_m_penable),
    .o_soc_periph_targ_syscfg_apb_m_pprot(o_soc_periph_targ_syscfg_apb_m_pprot),
    .i_soc_periph_targ_syscfg_apb_m_prdata(i_soc_periph_targ_syscfg_apb_m_prdata),
    .i_soc_periph_targ_syscfg_apb_m_pready(i_soc_periph_targ_syscfg_apb_m_pready),
    .o_soc_periph_targ_syscfg_apb_m_psel(o_soc_periph_targ_syscfg_apb_m_psel),
    .i_soc_periph_targ_syscfg_apb_m_pslverr(i_soc_periph_targ_syscfg_apb_m_pslverr),
    .o_soc_periph_targ_syscfg_apb_m_pstrb(o_soc_periph_targ_syscfg_apb_m_pstrb),
    .o_soc_periph_targ_syscfg_apb_m_pwdata(o_soc_periph_targ_syscfg_apb_m_pwdata),
    .o_soc_periph_targ_syscfg_apb_m_pwrite(o_soc_periph_targ_syscfg_apb_m_pwrite)
);

endmodule
