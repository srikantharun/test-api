package spike_top_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;
  import svt_uvm_pkg::*;
  import svt_axi_uvm_pkg::*;
  import spike_seq_pkg::*;

  `include "spike_top_config.sv"
  `include "spike_top_env.sv"

endpackage : spike_top_pkg
