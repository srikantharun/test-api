// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_ddr_west
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_ddr_west (
    input  wire                                        i_ddr_wpll_aon_clk,
    input  wire                                        i_ddr_wpll_aon_rst_n,
    output chip_pkg::chip_syscfg_addr_t                o_ddr_wpll_targ_syscfg_apb_m_paddr,
    output logic                                       o_ddr_wpll_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_ddr_wpll_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_ddr_wpll_targ_syscfg_apb_m_prdata,
    input  logic                                       i_ddr_wpll_targ_syscfg_apb_m_pready,
    output logic                                       o_ddr_wpll_targ_syscfg_apb_m_psel,
    input  logic                                       i_ddr_wpll_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_ddr_wpll_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_ddr_wpll_targ_syscfg_apb_m_pwdata,
    output logic                                       o_ddr_wpll_targ_syscfg_apb_m_pwrite,
    input  logic [398:0]                               i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld,
    output logic [398:0]                               o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld,
    input  logic [398:0]                               i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld,
    output logic [398:0]                               o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld,
    input  logic [398:0]                               i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld,
    output logic [398:0]                               o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld,
    input  logic [398:0]                               i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld,
    output logic [398:0]                               o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld,
    input  logic [146:0]                               i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld,
    output logic [146:0]                               o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld,
    input  wire                                        i_lpddr_graph_0_aon_clk,
    input  wire                                        i_lpddr_graph_0_aon_rst_n,
    output logic                                       o_lpddr_graph_0_cfg_pwr_idle_val,
    output logic                                       o_lpddr_graph_0_cfg_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_0_cfg_pwr_idle_req,
    input  wire                                        i_lpddr_graph_0_clk,
    input  wire                                        i_lpddr_graph_0_clken,
    output logic                                       o_lpddr_graph_0_pwr_idle_val,
    output logic                                       o_lpddr_graph_0_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_0_pwr_idle_req,
    input  wire                                        i_lpddr_graph_0_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t   o_lpddr_graph_0_targ_cfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_0_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_0_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   i_lpddr_graph_0_targ_cfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_0_targ_cfg_apb_m_pready,
    output logic                                       o_lpddr_graph_0_targ_cfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_0_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                 o_lpddr_graph_0_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   o_lpddr_graph_0_targ_cfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_0_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_0_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_0_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_0_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_0_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_0_targ_ht_axi_m_arlen,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_0_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_0_targ_ht_axi_m_arqos,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_0_targ_ht_axi_m_arsize,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_0_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_0_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_0_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_0_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_0_targ_ht_axi_m_awlen,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_0_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_0_targ_ht_axi_m_awqos,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_0_targ_ht_axi_m_awsize,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_0_targ_ht_axi_m_bid,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_0_targ_ht_axi_m_bresp,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   i_lpddr_graph_0_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_0_targ_ht_axi_m_rid,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_rlast,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_0_targ_ht_axi_m_rresp,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   o_lpddr_graph_0_targ_ht_axi_m_wdata,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_wlast,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t   o_lpddr_graph_0_targ_ht_axi_m_wstrb,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                o_lpddr_graph_0_targ_syscfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_lpddr_graph_0_targ_syscfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_0_targ_syscfg_apb_m_pready,
    output logic                                       o_lpddr_graph_0_targ_syscfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_lpddr_graph_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_lpddr_graph_0_targ_syscfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_0_targ_syscfg_apb_m_pwrite,
    input  wire                                        i_lpddr_graph_1_aon_clk,
    input  wire                                        i_lpddr_graph_1_aon_rst_n,
    output logic                                       o_lpddr_graph_1_cfg_pwr_idle_val,
    output logic                                       o_lpddr_graph_1_cfg_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_1_cfg_pwr_idle_req,
    input  wire                                        i_lpddr_graph_1_clk,
    input  wire                                        i_lpddr_graph_1_clken,
    output logic                                       o_lpddr_graph_1_pwr_idle_val,
    output logic                                       o_lpddr_graph_1_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_1_pwr_idle_req,
    input  wire                                        i_lpddr_graph_1_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t   o_lpddr_graph_1_targ_cfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_1_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_1_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   i_lpddr_graph_1_targ_cfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_1_targ_cfg_apb_m_pready,
    output logic                                       o_lpddr_graph_1_targ_cfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_1_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                 o_lpddr_graph_1_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   o_lpddr_graph_1_targ_cfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_1_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_1_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_1_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_1_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_1_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_1_targ_ht_axi_m_arlen,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_1_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_1_targ_ht_axi_m_arqos,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_1_targ_ht_axi_m_arsize,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_1_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_1_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_1_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_1_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_1_targ_ht_axi_m_awlen,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_1_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_1_targ_ht_axi_m_awqos,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_1_targ_ht_axi_m_awsize,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_1_targ_ht_axi_m_bid,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_1_targ_ht_axi_m_bresp,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   i_lpddr_graph_1_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_1_targ_ht_axi_m_rid,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_rlast,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_1_targ_ht_axi_m_rresp,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   o_lpddr_graph_1_targ_ht_axi_m_wdata,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_wlast,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t   o_lpddr_graph_1_targ_ht_axi_m_wstrb,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                o_lpddr_graph_1_targ_syscfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_lpddr_graph_1_targ_syscfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_1_targ_syscfg_apb_m_pready,
    output logic                                       o_lpddr_graph_1_targ_syscfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_lpddr_graph_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_lpddr_graph_1_targ_syscfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_1_targ_syscfg_apb_m_pwrite,
    input  wire                                        i_lpddr_graph_2_aon_clk,
    input  wire                                        i_lpddr_graph_2_aon_rst_n,
    output logic                                       o_lpddr_graph_2_cfg_pwr_idle_val,
    output logic                                       o_lpddr_graph_2_cfg_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_2_cfg_pwr_idle_req,
    input  wire                                        i_lpddr_graph_2_clk,
    input  wire                                        i_lpddr_graph_2_clken,
    output logic                                       o_lpddr_graph_2_pwr_idle_val,
    output logic                                       o_lpddr_graph_2_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_2_pwr_idle_req,
    input  wire                                        i_lpddr_graph_2_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t   o_lpddr_graph_2_targ_cfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_2_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_2_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   i_lpddr_graph_2_targ_cfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_2_targ_cfg_apb_m_pready,
    output logic                                       o_lpddr_graph_2_targ_cfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_2_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                 o_lpddr_graph_2_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   o_lpddr_graph_2_targ_cfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_2_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_2_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_2_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_2_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_2_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_2_targ_ht_axi_m_arlen,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_2_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_2_targ_ht_axi_m_arqos,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_2_targ_ht_axi_m_arsize,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_2_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_2_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_2_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_2_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_2_targ_ht_axi_m_awlen,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_2_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_2_targ_ht_axi_m_awqos,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_2_targ_ht_axi_m_awsize,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_2_targ_ht_axi_m_bid,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_2_targ_ht_axi_m_bresp,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   i_lpddr_graph_2_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_2_targ_ht_axi_m_rid,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_rlast,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_2_targ_ht_axi_m_rresp,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   o_lpddr_graph_2_targ_ht_axi_m_wdata,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_wlast,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t   o_lpddr_graph_2_targ_ht_axi_m_wstrb,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                o_lpddr_graph_2_targ_syscfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_lpddr_graph_2_targ_syscfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_2_targ_syscfg_apb_m_pready,
    output logic                                       o_lpddr_graph_2_targ_syscfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_lpddr_graph_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_lpddr_graph_2_targ_syscfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_2_targ_syscfg_apb_m_pwrite,
    input  wire                                        i_lpddr_graph_3_aon_clk,
    input  wire                                        i_lpddr_graph_3_aon_rst_n,
    output logic                                       o_lpddr_graph_3_cfg_pwr_idle_val,
    output logic                                       o_lpddr_graph_3_cfg_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_3_cfg_pwr_idle_req,
    input  wire                                        i_lpddr_graph_3_clk,
    input  wire                                        i_lpddr_graph_3_clken,
    output logic                                       o_lpddr_graph_3_pwr_idle_val,
    output logic                                       o_lpddr_graph_3_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_3_pwr_idle_req,
    input  wire                                        i_lpddr_graph_3_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t   o_lpddr_graph_3_targ_cfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_3_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_3_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   i_lpddr_graph_3_targ_cfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_3_targ_cfg_apb_m_pready,
    output logic                                       o_lpddr_graph_3_targ_cfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_3_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                 o_lpddr_graph_3_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   o_lpddr_graph_3_targ_cfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_3_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_3_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_3_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_3_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_3_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_3_targ_ht_axi_m_arlen,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_3_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_3_targ_ht_axi_m_arqos,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_3_targ_ht_axi_m_arsize,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_3_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_3_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_3_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_3_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_3_targ_ht_axi_m_awlen,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_3_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_3_targ_ht_axi_m_awqos,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_3_targ_ht_axi_m_awsize,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_3_targ_ht_axi_m_bid,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_3_targ_ht_axi_m_bresp,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   i_lpddr_graph_3_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_3_targ_ht_axi_m_rid,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_rlast,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_3_targ_ht_axi_m_rresp,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   o_lpddr_graph_3_targ_ht_axi_m_wdata,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_wlast,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t   o_lpddr_graph_3_targ_ht_axi_m_wstrb,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                o_lpddr_graph_3_targ_syscfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_lpddr_graph_3_targ_syscfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_3_targ_syscfg_apb_m_pready,
    output logic                                       o_lpddr_graph_3_targ_syscfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_lpddr_graph_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_lpddr_graph_3_targ_syscfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_3_targ_syscfg_apb_m_pwrite,
    input  wire                                        i_noc_clk,
    input  wire                                        i_noc_rst_n,
    input  logic                                       scan_en
);

    // Automated Address MSB fix: extra nets declaration
    logic[40:0] lpddr_graph_0_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] lpddr_graph_0_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] lpddr_graph_1_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] lpddr_graph_1_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] lpddr_graph_2_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] lpddr_graph_2_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] lpddr_graph_3_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] lpddr_graph_3_targ_ht_axi_m_awaddr_msb_fixed;

    // Automated Address MSB fix: Initiator-side assignments to extend addresses by 1 bit

    // Automated Address MSB fix: Target-side assignments to drop unused MSB
    assign o_lpddr_graph_0_targ_ht_axi_m_araddr = lpddr_graph_0_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_lpddr_graph_0_targ_ht_axi_m_awaddr = lpddr_graph_0_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_lpddr_graph_1_targ_ht_axi_m_araddr = lpddr_graph_1_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_lpddr_graph_1_targ_ht_axi_m_awaddr = lpddr_graph_1_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_lpddr_graph_2_targ_ht_axi_m_araddr = lpddr_graph_2_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_lpddr_graph_2_targ_ht_axi_m_awaddr = lpddr_graph_2_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_lpddr_graph_3_targ_ht_axi_m_araddr = lpddr_graph_3_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_lpddr_graph_3_targ_ht_axi_m_awaddr = lpddr_graph_3_targ_ht_axi_m_awaddr_msb_fixed[39:0];


    noc_art_ddr_west u_noc_art_ddr_west (
    .ddr_wpll_aon_clk(i_ddr_wpll_aon_clk),
    .ddr_wpll_aon_rst_n(i_ddr_wpll_aon_rst_n),
    .ddr_wpll_targ_syscfg_PAddr(o_ddr_wpll_targ_syscfg_apb_m_paddr),
    .ddr_wpll_targ_syscfg_PEnable(o_ddr_wpll_targ_syscfg_apb_m_penable),
    .ddr_wpll_targ_syscfg_PProt(o_ddr_wpll_targ_syscfg_apb_m_pprot),
    .ddr_wpll_targ_syscfg_PRData(i_ddr_wpll_targ_syscfg_apb_m_prdata),
    .ddr_wpll_targ_syscfg_PReady(i_ddr_wpll_targ_syscfg_apb_m_pready),
    .ddr_wpll_targ_syscfg_PSel(o_ddr_wpll_targ_syscfg_apb_m_psel),
    .ddr_wpll_targ_syscfg_PSlvErr(i_ddr_wpll_targ_syscfg_apb_m_pslverr),
    .ddr_wpll_targ_syscfg_PStrb(o_ddr_wpll_targ_syscfg_apb_m_pstrb),
    .ddr_wpll_targ_syscfg_PWData(o_ddr_wpll_targ_syscfg_apb_m_pwdata),
    .ddr_wpll_targ_syscfg_PWrite(o_ddr_wpll_targ_syscfg_apb_m_pwrite),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Data(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Head(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Rdy(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Tail(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Vld(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Data(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Head(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Rdy(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Tail(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Vld(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Data(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Head(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Rdy(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Tail(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Vld(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Data(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Head(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Rdy(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Tail(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Vld(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Data(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Head(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Rdy(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Tail(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Vld(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Data(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Head(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Rdy(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Tail(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Vld(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Data(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Head(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Rdy(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Tail(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Vld(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Data(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Head(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Rdy(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Tail(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Vld(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Data(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Head(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Rdy(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Tail(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Vld(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Data(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Head(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Rdy(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Tail(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Vld(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld),
    .lpddr_graph_0_aon_clk(i_lpddr_graph_0_aon_clk),
    .lpddr_graph_0_aon_rst_n(i_lpddr_graph_0_aon_rst_n),
    .lpddr_graph_0_cfg_pwr_Idle(o_lpddr_graph_0_cfg_pwr_idle_val),
    .lpddr_graph_0_cfg_pwr_IdleAck(o_lpddr_graph_0_cfg_pwr_idle_ack),
    .lpddr_graph_0_cfg_pwr_IdleReq(i_lpddr_graph_0_cfg_pwr_idle_req),
    .lpddr_graph_0_clk(i_lpddr_graph_0_clk),
    .lpddr_graph_0_clken(i_lpddr_graph_0_clken),
    .lpddr_graph_0_pwr_Idle(o_lpddr_graph_0_pwr_idle_val),
    .lpddr_graph_0_pwr_IdleAck(o_lpddr_graph_0_pwr_idle_ack),
    .lpddr_graph_0_pwr_IdleReq(i_lpddr_graph_0_pwr_idle_req),
    .lpddr_graph_0_rst_n(i_lpddr_graph_0_rst_n),
    .lpddr_graph_0_targ_cfg_PAddr(o_lpddr_graph_0_targ_cfg_apb_m_paddr),
    .lpddr_graph_0_targ_cfg_PEnable(o_lpddr_graph_0_targ_cfg_apb_m_penable),
    .lpddr_graph_0_targ_cfg_PProt(o_lpddr_graph_0_targ_cfg_apb_m_pprot),
    .lpddr_graph_0_targ_cfg_PRData(i_lpddr_graph_0_targ_cfg_apb_m_prdata),
    .lpddr_graph_0_targ_cfg_PReady(i_lpddr_graph_0_targ_cfg_apb_m_pready),
    .lpddr_graph_0_targ_cfg_PSel(o_lpddr_graph_0_targ_cfg_apb_m_psel),
    .lpddr_graph_0_targ_cfg_PSlvErr(i_lpddr_graph_0_targ_cfg_apb_m_pslverr),
    .lpddr_graph_0_targ_cfg_PStrb(o_lpddr_graph_0_targ_cfg_apb_m_pstrb),
    .lpddr_graph_0_targ_cfg_PWData(o_lpddr_graph_0_targ_cfg_apb_m_pwdata),
    .lpddr_graph_0_targ_cfg_PWrite(o_lpddr_graph_0_targ_cfg_apb_m_pwrite),
    .lpddr_graph_0_targ_ht_Ar_Addr(lpddr_graph_0_targ_ht_axi_m_araddr_msb_fixed),
    .lpddr_graph_0_targ_ht_Ar_Burst(o_lpddr_graph_0_targ_ht_axi_m_arburst),
    .lpddr_graph_0_targ_ht_Ar_Cache(o_lpddr_graph_0_targ_ht_axi_m_arcache),
    .lpddr_graph_0_targ_ht_Ar_Id(o_lpddr_graph_0_targ_ht_axi_m_arid),
    .lpddr_graph_0_targ_ht_Ar_Len(o_lpddr_graph_0_targ_ht_axi_m_arlen),
    .lpddr_graph_0_targ_ht_Ar_Lock(o_lpddr_graph_0_targ_ht_axi_m_arlock),
    .lpddr_graph_0_targ_ht_Ar_Prot(o_lpddr_graph_0_targ_ht_axi_m_arprot),
    .lpddr_graph_0_targ_ht_Ar_Qos(o_lpddr_graph_0_targ_ht_axi_m_arqos),
    .lpddr_graph_0_targ_ht_Ar_Ready(i_lpddr_graph_0_targ_ht_axi_m_arready),
    .lpddr_graph_0_targ_ht_Ar_Size(o_lpddr_graph_0_targ_ht_axi_m_arsize),
    .lpddr_graph_0_targ_ht_Ar_Valid(o_lpddr_graph_0_targ_ht_axi_m_arvalid),
    .lpddr_graph_0_targ_ht_Aw_Addr(lpddr_graph_0_targ_ht_axi_m_awaddr_msb_fixed),
    .lpddr_graph_0_targ_ht_Aw_Burst(o_lpddr_graph_0_targ_ht_axi_m_awburst),
    .lpddr_graph_0_targ_ht_Aw_Cache(o_lpddr_graph_0_targ_ht_axi_m_awcache),
    .lpddr_graph_0_targ_ht_Aw_Id(o_lpddr_graph_0_targ_ht_axi_m_awid),
    .lpddr_graph_0_targ_ht_Aw_Len(o_lpddr_graph_0_targ_ht_axi_m_awlen),
    .lpddr_graph_0_targ_ht_Aw_Lock(o_lpddr_graph_0_targ_ht_axi_m_awlock),
    .lpddr_graph_0_targ_ht_Aw_Prot(o_lpddr_graph_0_targ_ht_axi_m_awprot),
    .lpddr_graph_0_targ_ht_Aw_Qos(o_lpddr_graph_0_targ_ht_axi_m_awqos),
    .lpddr_graph_0_targ_ht_Aw_Ready(i_lpddr_graph_0_targ_ht_axi_m_awready),
    .lpddr_graph_0_targ_ht_Aw_Size(o_lpddr_graph_0_targ_ht_axi_m_awsize),
    .lpddr_graph_0_targ_ht_Aw_Valid(o_lpddr_graph_0_targ_ht_axi_m_awvalid),
    .lpddr_graph_0_targ_ht_B_Id(i_lpddr_graph_0_targ_ht_axi_m_bid),
    .lpddr_graph_0_targ_ht_B_Ready(o_lpddr_graph_0_targ_ht_axi_m_bready),
    .lpddr_graph_0_targ_ht_B_Resp(i_lpddr_graph_0_targ_ht_axi_m_bresp),
    .lpddr_graph_0_targ_ht_B_Valid(i_lpddr_graph_0_targ_ht_axi_m_bvalid),
    .lpddr_graph_0_targ_ht_R_Data(i_lpddr_graph_0_targ_ht_axi_m_rdata),
    .lpddr_graph_0_targ_ht_R_Id(i_lpddr_graph_0_targ_ht_axi_m_rid),
    .lpddr_graph_0_targ_ht_R_Last(i_lpddr_graph_0_targ_ht_axi_m_rlast),
    .lpddr_graph_0_targ_ht_R_Ready(o_lpddr_graph_0_targ_ht_axi_m_rready),
    .lpddr_graph_0_targ_ht_R_Resp(i_lpddr_graph_0_targ_ht_axi_m_rresp),
    .lpddr_graph_0_targ_ht_R_Valid(i_lpddr_graph_0_targ_ht_axi_m_rvalid),
    .lpddr_graph_0_targ_ht_W_Data(o_lpddr_graph_0_targ_ht_axi_m_wdata),
    .lpddr_graph_0_targ_ht_W_Last(o_lpddr_graph_0_targ_ht_axi_m_wlast),
    .lpddr_graph_0_targ_ht_W_Ready(i_lpddr_graph_0_targ_ht_axi_m_wready),
    .lpddr_graph_0_targ_ht_W_Strb(o_lpddr_graph_0_targ_ht_axi_m_wstrb),
    .lpddr_graph_0_targ_ht_W_Valid(o_lpddr_graph_0_targ_ht_axi_m_wvalid),
    .lpddr_graph_0_targ_syscfg_PAddr(o_lpddr_graph_0_targ_syscfg_apb_m_paddr),
    .lpddr_graph_0_targ_syscfg_PEnable(o_lpddr_graph_0_targ_syscfg_apb_m_penable),
    .lpddr_graph_0_targ_syscfg_PProt(o_lpddr_graph_0_targ_syscfg_apb_m_pprot),
    .lpddr_graph_0_targ_syscfg_PRData(i_lpddr_graph_0_targ_syscfg_apb_m_prdata),
    .lpddr_graph_0_targ_syscfg_PReady(i_lpddr_graph_0_targ_syscfg_apb_m_pready),
    .lpddr_graph_0_targ_syscfg_PSel(o_lpddr_graph_0_targ_syscfg_apb_m_psel),
    .lpddr_graph_0_targ_syscfg_PSlvErr(i_lpddr_graph_0_targ_syscfg_apb_m_pslverr),
    .lpddr_graph_0_targ_syscfg_PStrb(o_lpddr_graph_0_targ_syscfg_apb_m_pstrb),
    .lpddr_graph_0_targ_syscfg_PWData(o_lpddr_graph_0_targ_syscfg_apb_m_pwdata),
    .lpddr_graph_0_targ_syscfg_PWrite(o_lpddr_graph_0_targ_syscfg_apb_m_pwrite),
    .lpddr_graph_1_aon_clk(i_lpddr_graph_1_aon_clk),
    .lpddr_graph_1_aon_rst_n(i_lpddr_graph_1_aon_rst_n),
    .lpddr_graph_1_cfg_pwr_Idle(o_lpddr_graph_1_cfg_pwr_idle_val),
    .lpddr_graph_1_cfg_pwr_IdleAck(o_lpddr_graph_1_cfg_pwr_idle_ack),
    .lpddr_graph_1_cfg_pwr_IdleReq(i_lpddr_graph_1_cfg_pwr_idle_req),
    .lpddr_graph_1_clk(i_lpddr_graph_1_clk),
    .lpddr_graph_1_clken(i_lpddr_graph_1_clken),
    .lpddr_graph_1_pwr_Idle(o_lpddr_graph_1_pwr_idle_val),
    .lpddr_graph_1_pwr_IdleAck(o_lpddr_graph_1_pwr_idle_ack),
    .lpddr_graph_1_pwr_IdleReq(i_lpddr_graph_1_pwr_idle_req),
    .lpddr_graph_1_rst_n(i_lpddr_graph_1_rst_n),
    .lpddr_graph_1_targ_cfg_PAddr(o_lpddr_graph_1_targ_cfg_apb_m_paddr),
    .lpddr_graph_1_targ_cfg_PEnable(o_lpddr_graph_1_targ_cfg_apb_m_penable),
    .lpddr_graph_1_targ_cfg_PProt(o_lpddr_graph_1_targ_cfg_apb_m_pprot),
    .lpddr_graph_1_targ_cfg_PRData(i_lpddr_graph_1_targ_cfg_apb_m_prdata),
    .lpddr_graph_1_targ_cfg_PReady(i_lpddr_graph_1_targ_cfg_apb_m_pready),
    .lpddr_graph_1_targ_cfg_PSel(o_lpddr_graph_1_targ_cfg_apb_m_psel),
    .lpddr_graph_1_targ_cfg_PSlvErr(i_lpddr_graph_1_targ_cfg_apb_m_pslverr),
    .lpddr_graph_1_targ_cfg_PStrb(o_lpddr_graph_1_targ_cfg_apb_m_pstrb),
    .lpddr_graph_1_targ_cfg_PWData(o_lpddr_graph_1_targ_cfg_apb_m_pwdata),
    .lpddr_graph_1_targ_cfg_PWrite(o_lpddr_graph_1_targ_cfg_apb_m_pwrite),
    .lpddr_graph_1_targ_ht_Ar_Addr(lpddr_graph_1_targ_ht_axi_m_araddr_msb_fixed),
    .lpddr_graph_1_targ_ht_Ar_Burst(o_lpddr_graph_1_targ_ht_axi_m_arburst),
    .lpddr_graph_1_targ_ht_Ar_Cache(o_lpddr_graph_1_targ_ht_axi_m_arcache),
    .lpddr_graph_1_targ_ht_Ar_Id(o_lpddr_graph_1_targ_ht_axi_m_arid),
    .lpddr_graph_1_targ_ht_Ar_Len(o_lpddr_graph_1_targ_ht_axi_m_arlen),
    .lpddr_graph_1_targ_ht_Ar_Lock(o_lpddr_graph_1_targ_ht_axi_m_arlock),
    .lpddr_graph_1_targ_ht_Ar_Prot(o_lpddr_graph_1_targ_ht_axi_m_arprot),
    .lpddr_graph_1_targ_ht_Ar_Qos(o_lpddr_graph_1_targ_ht_axi_m_arqos),
    .lpddr_graph_1_targ_ht_Ar_Ready(i_lpddr_graph_1_targ_ht_axi_m_arready),
    .lpddr_graph_1_targ_ht_Ar_Size(o_lpddr_graph_1_targ_ht_axi_m_arsize),
    .lpddr_graph_1_targ_ht_Ar_Valid(o_lpddr_graph_1_targ_ht_axi_m_arvalid),
    .lpddr_graph_1_targ_ht_Aw_Addr(lpddr_graph_1_targ_ht_axi_m_awaddr_msb_fixed),
    .lpddr_graph_1_targ_ht_Aw_Burst(o_lpddr_graph_1_targ_ht_axi_m_awburst),
    .lpddr_graph_1_targ_ht_Aw_Cache(o_lpddr_graph_1_targ_ht_axi_m_awcache),
    .lpddr_graph_1_targ_ht_Aw_Id(o_lpddr_graph_1_targ_ht_axi_m_awid),
    .lpddr_graph_1_targ_ht_Aw_Len(o_lpddr_graph_1_targ_ht_axi_m_awlen),
    .lpddr_graph_1_targ_ht_Aw_Lock(o_lpddr_graph_1_targ_ht_axi_m_awlock),
    .lpddr_graph_1_targ_ht_Aw_Prot(o_lpddr_graph_1_targ_ht_axi_m_awprot),
    .lpddr_graph_1_targ_ht_Aw_Qos(o_lpddr_graph_1_targ_ht_axi_m_awqos),
    .lpddr_graph_1_targ_ht_Aw_Ready(i_lpddr_graph_1_targ_ht_axi_m_awready),
    .lpddr_graph_1_targ_ht_Aw_Size(o_lpddr_graph_1_targ_ht_axi_m_awsize),
    .lpddr_graph_1_targ_ht_Aw_Valid(o_lpddr_graph_1_targ_ht_axi_m_awvalid),
    .lpddr_graph_1_targ_ht_B_Id(i_lpddr_graph_1_targ_ht_axi_m_bid),
    .lpddr_graph_1_targ_ht_B_Ready(o_lpddr_graph_1_targ_ht_axi_m_bready),
    .lpddr_graph_1_targ_ht_B_Resp(i_lpddr_graph_1_targ_ht_axi_m_bresp),
    .lpddr_graph_1_targ_ht_B_Valid(i_lpddr_graph_1_targ_ht_axi_m_bvalid),
    .lpddr_graph_1_targ_ht_R_Data(i_lpddr_graph_1_targ_ht_axi_m_rdata),
    .lpddr_graph_1_targ_ht_R_Id(i_lpddr_graph_1_targ_ht_axi_m_rid),
    .lpddr_graph_1_targ_ht_R_Last(i_lpddr_graph_1_targ_ht_axi_m_rlast),
    .lpddr_graph_1_targ_ht_R_Ready(o_lpddr_graph_1_targ_ht_axi_m_rready),
    .lpddr_graph_1_targ_ht_R_Resp(i_lpddr_graph_1_targ_ht_axi_m_rresp),
    .lpddr_graph_1_targ_ht_R_Valid(i_lpddr_graph_1_targ_ht_axi_m_rvalid),
    .lpddr_graph_1_targ_ht_W_Data(o_lpddr_graph_1_targ_ht_axi_m_wdata),
    .lpddr_graph_1_targ_ht_W_Last(o_lpddr_graph_1_targ_ht_axi_m_wlast),
    .lpddr_graph_1_targ_ht_W_Ready(i_lpddr_graph_1_targ_ht_axi_m_wready),
    .lpddr_graph_1_targ_ht_W_Strb(o_lpddr_graph_1_targ_ht_axi_m_wstrb),
    .lpddr_graph_1_targ_ht_W_Valid(o_lpddr_graph_1_targ_ht_axi_m_wvalid),
    .lpddr_graph_1_targ_syscfg_PAddr(o_lpddr_graph_1_targ_syscfg_apb_m_paddr),
    .lpddr_graph_1_targ_syscfg_PEnable(o_lpddr_graph_1_targ_syscfg_apb_m_penable),
    .lpddr_graph_1_targ_syscfg_PProt(o_lpddr_graph_1_targ_syscfg_apb_m_pprot),
    .lpddr_graph_1_targ_syscfg_PRData(i_lpddr_graph_1_targ_syscfg_apb_m_prdata),
    .lpddr_graph_1_targ_syscfg_PReady(i_lpddr_graph_1_targ_syscfg_apb_m_pready),
    .lpddr_graph_1_targ_syscfg_PSel(o_lpddr_graph_1_targ_syscfg_apb_m_psel),
    .lpddr_graph_1_targ_syscfg_PSlvErr(i_lpddr_graph_1_targ_syscfg_apb_m_pslverr),
    .lpddr_graph_1_targ_syscfg_PStrb(o_lpddr_graph_1_targ_syscfg_apb_m_pstrb),
    .lpddr_graph_1_targ_syscfg_PWData(o_lpddr_graph_1_targ_syscfg_apb_m_pwdata),
    .lpddr_graph_1_targ_syscfg_PWrite(o_lpddr_graph_1_targ_syscfg_apb_m_pwrite),
    .lpddr_graph_2_aon_clk(i_lpddr_graph_2_aon_clk),
    .lpddr_graph_2_aon_rst_n(i_lpddr_graph_2_aon_rst_n),
    .lpddr_graph_2_cfg_pwr_Idle(o_lpddr_graph_2_cfg_pwr_idle_val),
    .lpddr_graph_2_cfg_pwr_IdleAck(o_lpddr_graph_2_cfg_pwr_idle_ack),
    .lpddr_graph_2_cfg_pwr_IdleReq(i_lpddr_graph_2_cfg_pwr_idle_req),
    .lpddr_graph_2_clk(i_lpddr_graph_2_clk),
    .lpddr_graph_2_clken(i_lpddr_graph_2_clken),
    .lpddr_graph_2_pwr_Idle(o_lpddr_graph_2_pwr_idle_val),
    .lpddr_graph_2_pwr_IdleAck(o_lpddr_graph_2_pwr_idle_ack),
    .lpddr_graph_2_pwr_IdleReq(i_lpddr_graph_2_pwr_idle_req),
    .lpddr_graph_2_rst_n(i_lpddr_graph_2_rst_n),
    .lpddr_graph_2_targ_cfg_PAddr(o_lpddr_graph_2_targ_cfg_apb_m_paddr),
    .lpddr_graph_2_targ_cfg_PEnable(o_lpddr_graph_2_targ_cfg_apb_m_penable),
    .lpddr_graph_2_targ_cfg_PProt(o_lpddr_graph_2_targ_cfg_apb_m_pprot),
    .lpddr_graph_2_targ_cfg_PRData(i_lpddr_graph_2_targ_cfg_apb_m_prdata),
    .lpddr_graph_2_targ_cfg_PReady(i_lpddr_graph_2_targ_cfg_apb_m_pready),
    .lpddr_graph_2_targ_cfg_PSel(o_lpddr_graph_2_targ_cfg_apb_m_psel),
    .lpddr_graph_2_targ_cfg_PSlvErr(i_lpddr_graph_2_targ_cfg_apb_m_pslverr),
    .lpddr_graph_2_targ_cfg_PStrb(o_lpddr_graph_2_targ_cfg_apb_m_pstrb),
    .lpddr_graph_2_targ_cfg_PWData(o_lpddr_graph_2_targ_cfg_apb_m_pwdata),
    .lpddr_graph_2_targ_cfg_PWrite(o_lpddr_graph_2_targ_cfg_apb_m_pwrite),
    .lpddr_graph_2_targ_ht_Ar_Addr(lpddr_graph_2_targ_ht_axi_m_araddr_msb_fixed),
    .lpddr_graph_2_targ_ht_Ar_Burst(o_lpddr_graph_2_targ_ht_axi_m_arburst),
    .lpddr_graph_2_targ_ht_Ar_Cache(o_lpddr_graph_2_targ_ht_axi_m_arcache),
    .lpddr_graph_2_targ_ht_Ar_Id(o_lpddr_graph_2_targ_ht_axi_m_arid),
    .lpddr_graph_2_targ_ht_Ar_Len(o_lpddr_graph_2_targ_ht_axi_m_arlen),
    .lpddr_graph_2_targ_ht_Ar_Lock(o_lpddr_graph_2_targ_ht_axi_m_arlock),
    .lpddr_graph_2_targ_ht_Ar_Prot(o_lpddr_graph_2_targ_ht_axi_m_arprot),
    .lpddr_graph_2_targ_ht_Ar_Qos(o_lpddr_graph_2_targ_ht_axi_m_arqos),
    .lpddr_graph_2_targ_ht_Ar_Ready(i_lpddr_graph_2_targ_ht_axi_m_arready),
    .lpddr_graph_2_targ_ht_Ar_Size(o_lpddr_graph_2_targ_ht_axi_m_arsize),
    .lpddr_graph_2_targ_ht_Ar_Valid(o_lpddr_graph_2_targ_ht_axi_m_arvalid),
    .lpddr_graph_2_targ_ht_Aw_Addr(lpddr_graph_2_targ_ht_axi_m_awaddr_msb_fixed),
    .lpddr_graph_2_targ_ht_Aw_Burst(o_lpddr_graph_2_targ_ht_axi_m_awburst),
    .lpddr_graph_2_targ_ht_Aw_Cache(o_lpddr_graph_2_targ_ht_axi_m_awcache),
    .lpddr_graph_2_targ_ht_Aw_Id(o_lpddr_graph_2_targ_ht_axi_m_awid),
    .lpddr_graph_2_targ_ht_Aw_Len(o_lpddr_graph_2_targ_ht_axi_m_awlen),
    .lpddr_graph_2_targ_ht_Aw_Lock(o_lpddr_graph_2_targ_ht_axi_m_awlock),
    .lpddr_graph_2_targ_ht_Aw_Prot(o_lpddr_graph_2_targ_ht_axi_m_awprot),
    .lpddr_graph_2_targ_ht_Aw_Qos(o_lpddr_graph_2_targ_ht_axi_m_awqos),
    .lpddr_graph_2_targ_ht_Aw_Ready(i_lpddr_graph_2_targ_ht_axi_m_awready),
    .lpddr_graph_2_targ_ht_Aw_Size(o_lpddr_graph_2_targ_ht_axi_m_awsize),
    .lpddr_graph_2_targ_ht_Aw_Valid(o_lpddr_graph_2_targ_ht_axi_m_awvalid),
    .lpddr_graph_2_targ_ht_B_Id(i_lpddr_graph_2_targ_ht_axi_m_bid),
    .lpddr_graph_2_targ_ht_B_Ready(o_lpddr_graph_2_targ_ht_axi_m_bready),
    .lpddr_graph_2_targ_ht_B_Resp(i_lpddr_graph_2_targ_ht_axi_m_bresp),
    .lpddr_graph_2_targ_ht_B_Valid(i_lpddr_graph_2_targ_ht_axi_m_bvalid),
    .lpddr_graph_2_targ_ht_R_Data(i_lpddr_graph_2_targ_ht_axi_m_rdata),
    .lpddr_graph_2_targ_ht_R_Id(i_lpddr_graph_2_targ_ht_axi_m_rid),
    .lpddr_graph_2_targ_ht_R_Last(i_lpddr_graph_2_targ_ht_axi_m_rlast),
    .lpddr_graph_2_targ_ht_R_Ready(o_lpddr_graph_2_targ_ht_axi_m_rready),
    .lpddr_graph_2_targ_ht_R_Resp(i_lpddr_graph_2_targ_ht_axi_m_rresp),
    .lpddr_graph_2_targ_ht_R_Valid(i_lpddr_graph_2_targ_ht_axi_m_rvalid),
    .lpddr_graph_2_targ_ht_W_Data(o_lpddr_graph_2_targ_ht_axi_m_wdata),
    .lpddr_graph_2_targ_ht_W_Last(o_lpddr_graph_2_targ_ht_axi_m_wlast),
    .lpddr_graph_2_targ_ht_W_Ready(i_lpddr_graph_2_targ_ht_axi_m_wready),
    .lpddr_graph_2_targ_ht_W_Strb(o_lpddr_graph_2_targ_ht_axi_m_wstrb),
    .lpddr_graph_2_targ_ht_W_Valid(o_lpddr_graph_2_targ_ht_axi_m_wvalid),
    .lpddr_graph_2_targ_syscfg_PAddr(o_lpddr_graph_2_targ_syscfg_apb_m_paddr),
    .lpddr_graph_2_targ_syscfg_PEnable(o_lpddr_graph_2_targ_syscfg_apb_m_penable),
    .lpddr_graph_2_targ_syscfg_PProt(o_lpddr_graph_2_targ_syscfg_apb_m_pprot),
    .lpddr_graph_2_targ_syscfg_PRData(i_lpddr_graph_2_targ_syscfg_apb_m_prdata),
    .lpddr_graph_2_targ_syscfg_PReady(i_lpddr_graph_2_targ_syscfg_apb_m_pready),
    .lpddr_graph_2_targ_syscfg_PSel(o_lpddr_graph_2_targ_syscfg_apb_m_psel),
    .lpddr_graph_2_targ_syscfg_PSlvErr(i_lpddr_graph_2_targ_syscfg_apb_m_pslverr),
    .lpddr_graph_2_targ_syscfg_PStrb(o_lpddr_graph_2_targ_syscfg_apb_m_pstrb),
    .lpddr_graph_2_targ_syscfg_PWData(o_lpddr_graph_2_targ_syscfg_apb_m_pwdata),
    .lpddr_graph_2_targ_syscfg_PWrite(o_lpddr_graph_2_targ_syscfg_apb_m_pwrite),
    .lpddr_graph_3_aon_clk(i_lpddr_graph_3_aon_clk),
    .lpddr_graph_3_aon_rst_n(i_lpddr_graph_3_aon_rst_n),
    .lpddr_graph_3_cfg_pwr_Idle(o_lpddr_graph_3_cfg_pwr_idle_val),
    .lpddr_graph_3_cfg_pwr_IdleAck(o_lpddr_graph_3_cfg_pwr_idle_ack),
    .lpddr_graph_3_cfg_pwr_IdleReq(i_lpddr_graph_3_cfg_pwr_idle_req),
    .lpddr_graph_3_clk(i_lpddr_graph_3_clk),
    .lpddr_graph_3_clken(i_lpddr_graph_3_clken),
    .lpddr_graph_3_pwr_Idle(o_lpddr_graph_3_pwr_idle_val),
    .lpddr_graph_3_pwr_IdleAck(o_lpddr_graph_3_pwr_idle_ack),
    .lpddr_graph_3_pwr_IdleReq(i_lpddr_graph_3_pwr_idle_req),
    .lpddr_graph_3_rst_n(i_lpddr_graph_3_rst_n),
    .lpddr_graph_3_targ_cfg_PAddr(o_lpddr_graph_3_targ_cfg_apb_m_paddr),
    .lpddr_graph_3_targ_cfg_PEnable(o_lpddr_graph_3_targ_cfg_apb_m_penable),
    .lpddr_graph_3_targ_cfg_PProt(o_lpddr_graph_3_targ_cfg_apb_m_pprot),
    .lpddr_graph_3_targ_cfg_PRData(i_lpddr_graph_3_targ_cfg_apb_m_prdata),
    .lpddr_graph_3_targ_cfg_PReady(i_lpddr_graph_3_targ_cfg_apb_m_pready),
    .lpddr_graph_3_targ_cfg_PSel(o_lpddr_graph_3_targ_cfg_apb_m_psel),
    .lpddr_graph_3_targ_cfg_PSlvErr(i_lpddr_graph_3_targ_cfg_apb_m_pslverr),
    .lpddr_graph_3_targ_cfg_PStrb(o_lpddr_graph_3_targ_cfg_apb_m_pstrb),
    .lpddr_graph_3_targ_cfg_PWData(o_lpddr_graph_3_targ_cfg_apb_m_pwdata),
    .lpddr_graph_3_targ_cfg_PWrite(o_lpddr_graph_3_targ_cfg_apb_m_pwrite),
    .lpddr_graph_3_targ_ht_Ar_Addr(lpddr_graph_3_targ_ht_axi_m_araddr_msb_fixed),
    .lpddr_graph_3_targ_ht_Ar_Burst(o_lpddr_graph_3_targ_ht_axi_m_arburst),
    .lpddr_graph_3_targ_ht_Ar_Cache(o_lpddr_graph_3_targ_ht_axi_m_arcache),
    .lpddr_graph_3_targ_ht_Ar_Id(o_lpddr_graph_3_targ_ht_axi_m_arid),
    .lpddr_graph_3_targ_ht_Ar_Len(o_lpddr_graph_3_targ_ht_axi_m_arlen),
    .lpddr_graph_3_targ_ht_Ar_Lock(o_lpddr_graph_3_targ_ht_axi_m_arlock),
    .lpddr_graph_3_targ_ht_Ar_Prot(o_lpddr_graph_3_targ_ht_axi_m_arprot),
    .lpddr_graph_3_targ_ht_Ar_Qos(o_lpddr_graph_3_targ_ht_axi_m_arqos),
    .lpddr_graph_3_targ_ht_Ar_Ready(i_lpddr_graph_3_targ_ht_axi_m_arready),
    .lpddr_graph_3_targ_ht_Ar_Size(o_lpddr_graph_3_targ_ht_axi_m_arsize),
    .lpddr_graph_3_targ_ht_Ar_Valid(o_lpddr_graph_3_targ_ht_axi_m_arvalid),
    .lpddr_graph_3_targ_ht_Aw_Addr(lpddr_graph_3_targ_ht_axi_m_awaddr_msb_fixed),
    .lpddr_graph_3_targ_ht_Aw_Burst(o_lpddr_graph_3_targ_ht_axi_m_awburst),
    .lpddr_graph_3_targ_ht_Aw_Cache(o_lpddr_graph_3_targ_ht_axi_m_awcache),
    .lpddr_graph_3_targ_ht_Aw_Id(o_lpddr_graph_3_targ_ht_axi_m_awid),
    .lpddr_graph_3_targ_ht_Aw_Len(o_lpddr_graph_3_targ_ht_axi_m_awlen),
    .lpddr_graph_3_targ_ht_Aw_Lock(o_lpddr_graph_3_targ_ht_axi_m_awlock),
    .lpddr_graph_3_targ_ht_Aw_Prot(o_lpddr_graph_3_targ_ht_axi_m_awprot),
    .lpddr_graph_3_targ_ht_Aw_Qos(o_lpddr_graph_3_targ_ht_axi_m_awqos),
    .lpddr_graph_3_targ_ht_Aw_Ready(i_lpddr_graph_3_targ_ht_axi_m_awready),
    .lpddr_graph_3_targ_ht_Aw_Size(o_lpddr_graph_3_targ_ht_axi_m_awsize),
    .lpddr_graph_3_targ_ht_Aw_Valid(o_lpddr_graph_3_targ_ht_axi_m_awvalid),
    .lpddr_graph_3_targ_ht_B_Id(i_lpddr_graph_3_targ_ht_axi_m_bid),
    .lpddr_graph_3_targ_ht_B_Ready(o_lpddr_graph_3_targ_ht_axi_m_bready),
    .lpddr_graph_3_targ_ht_B_Resp(i_lpddr_graph_3_targ_ht_axi_m_bresp),
    .lpddr_graph_3_targ_ht_B_Valid(i_lpddr_graph_3_targ_ht_axi_m_bvalid),
    .lpddr_graph_3_targ_ht_R_Data(i_lpddr_graph_3_targ_ht_axi_m_rdata),
    .lpddr_graph_3_targ_ht_R_Id(i_lpddr_graph_3_targ_ht_axi_m_rid),
    .lpddr_graph_3_targ_ht_R_Last(i_lpddr_graph_3_targ_ht_axi_m_rlast),
    .lpddr_graph_3_targ_ht_R_Ready(o_lpddr_graph_3_targ_ht_axi_m_rready),
    .lpddr_graph_3_targ_ht_R_Resp(i_lpddr_graph_3_targ_ht_axi_m_rresp),
    .lpddr_graph_3_targ_ht_R_Valid(i_lpddr_graph_3_targ_ht_axi_m_rvalid),
    .lpddr_graph_3_targ_ht_W_Data(o_lpddr_graph_3_targ_ht_axi_m_wdata),
    .lpddr_graph_3_targ_ht_W_Last(o_lpddr_graph_3_targ_ht_axi_m_wlast),
    .lpddr_graph_3_targ_ht_W_Ready(i_lpddr_graph_3_targ_ht_axi_m_wready),
    .lpddr_graph_3_targ_ht_W_Strb(o_lpddr_graph_3_targ_ht_axi_m_wstrb),
    .lpddr_graph_3_targ_ht_W_Valid(o_lpddr_graph_3_targ_ht_axi_m_wvalid),
    .lpddr_graph_3_targ_syscfg_PAddr(o_lpddr_graph_3_targ_syscfg_apb_m_paddr),
    .lpddr_graph_3_targ_syscfg_PEnable(o_lpddr_graph_3_targ_syscfg_apb_m_penable),
    .lpddr_graph_3_targ_syscfg_PProt(o_lpddr_graph_3_targ_syscfg_apb_m_pprot),
    .lpddr_graph_3_targ_syscfg_PRData(i_lpddr_graph_3_targ_syscfg_apb_m_prdata),
    .lpddr_graph_3_targ_syscfg_PReady(i_lpddr_graph_3_targ_syscfg_apb_m_pready),
    .lpddr_graph_3_targ_syscfg_PSel(o_lpddr_graph_3_targ_syscfg_apb_m_psel),
    .lpddr_graph_3_targ_syscfg_PSlvErr(i_lpddr_graph_3_targ_syscfg_apb_m_pslverr),
    .lpddr_graph_3_targ_syscfg_PStrb(o_lpddr_graph_3_targ_syscfg_apb_m_pstrb),
    .lpddr_graph_3_targ_syscfg_PWData(o_lpddr_graph_3_targ_syscfg_apb_m_pwdata),
    .lpddr_graph_3_targ_syscfg_PWrite(o_lpddr_graph_3_targ_syscfg_apb_m_pwrite),
    .noc_clk(i_noc_clk),
    .noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
);

endmodule
