// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: {{ cookiecutter.author_full_name }} <{{ cookiecutter.author_email }}>


/// TODO:__one_line_summary_of_{{ cookiecutter.ip_name }}_pkg__
///
package {{ cookiecutter.ip_name }}_pkg;

endpackage
