`ifndef RAL_DWC_DDRPHYA_PPGC0_P0_PKG
`define RAL_DWC_DDRPHYA_PPGC0_P0_PKG

package ral_DWC_DDRPHYA_PPGC0_p0_pkg;
import uvm_pkg::*;

class ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenCtrl extends uvm_reg;
	rand uvm_reg_field PpgcGenCtrl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PpgcGenCtrl: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PpgcGenCtrl");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PpgcGenCtrl = uvm_reg_field::type_id::create("PpgcGenCtrl",,get_full_name());
      this.PpgcGenCtrl.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenCtrl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenCtrl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiCtrl extends uvm_reg;
	rand uvm_reg_field PpgcGenDbiCtrl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PpgcGenDbiCtrl: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiCtrl");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PpgcGenDbiCtrl = uvm_reg_field::type_id::create("PpgcGenDbiCtrl",,get_full_name());
      this.PpgcGenDbiCtrl.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiCtrl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiCtrl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiConfig extends uvm_reg;
	rand uvm_reg_field PpgcGenDbiConfig;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PpgcGenDbiConfig: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiConfig");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PpgcGenDbiConfig = uvm_reg_field::type_id::create("PpgcGenDbiConfig",,get_full_name());
      this.PpgcGenDbiConfig.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiConfig)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiConfig


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel0 extends uvm_reg;
	rand uvm_reg_field PpgcGenLaneMuxSel0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PpgcGenLaneMuxSel0: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PpgcGenLaneMuxSel0 = uvm_reg_field::type_id::create("PpgcGenLaneMuxSel0",,get_full_name());
      this.PpgcGenLaneMuxSel0.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel1 extends uvm_reg;
	rand uvm_reg_field PpgcGenLaneMuxSel1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PpgcGenLaneMuxSel1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PpgcGenLaneMuxSel1 = uvm_reg_field::type_id::create("PpgcGenLaneMuxSel1",,get_full_name());
      this.PpgcGenLaneMuxSel1.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_EnPhyUpdZQCalUpdate extends uvm_reg;
	rand uvm_reg_field EnPhyUpdZQCalUpdate;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   EnPhyUpdZQCalUpdate: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_EnPhyUpdZQCalUpdate");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.EnPhyUpdZQCalUpdate = uvm_reg_field::type_id::create("EnPhyUpdZQCalUpdate",,get_full_name());
      this.EnPhyUpdZQCalUpdate.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_EnPhyUpdZQCalUpdate)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_EnPhyUpdZQCalUpdate


class ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterface extends uvm_reg;
	rand uvm_reg_field BlockDfiInterfaceEn;
	rand uvm_reg_field BlockDfiInterfaceStatusReset;
	rand uvm_reg_field PmuBusy;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   BlockDfiInterfaceEn: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   BlockDfiInterfaceStatusReset: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PmuBusy: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_BlockDfiInterface");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.BlockDfiInterfaceEn = uvm_reg_field::type_id::create("BlockDfiInterfaceEn",,get_full_name());
      this.BlockDfiInterfaceEn.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.BlockDfiInterfaceStatusReset = uvm_reg_field::type_id::create("BlockDfiInterfaceStatusReset",,get_full_name());
      this.BlockDfiInterfaceStatusReset.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.PmuBusy = uvm_reg_field::type_id::create("PmuBusy",,get_full_name());
      this.PmuBusy.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterface)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterface


class ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterfaceStatus extends uvm_reg;
	uvm_reg_field BlockDfiInterfaceStatus;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   BlockDfiInterfaceStatus: coverpoint {m_data[7:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd = {9'b????????1};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd = {9'b????????1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd = {9'b????????1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd = {9'b????????1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd = {9'b????????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd = {9'b????????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd = {9'b????????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd = {9'b????????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_BlockDfiInterfaceStatus");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.BlockDfiInterfaceStatus = uvm_reg_field::type_id::create("BlockDfiInterfaceStatus",,get_full_name());
      this.BlockDfiInterfaceStatus.configure(this, 8, 0, "RO", 1, 8'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterfaceStatus)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterfaceStatus


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiCustMode_p0 extends uvm_reg;
	rand uvm_reg_field DfiCustMode_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DfiCustMode_p0: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiCustMode_p0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DfiCustMode_p0 = uvm_reg_field::type_id::create("DfiCustMode_p0",,get_full_name());
      this.DfiCustMode_p0.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiCustMode_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiCustMode_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtMRL_p0 extends uvm_reg;
	rand uvm_reg_field HwtMRL_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   HwtMRL_p0: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_HwtMRL_p0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.HwtMRL_p0 = uvm_reg_field::type_id::create("HwtMRL_p0",,get_full_name());
      this.HwtMRL_p0.configure(this, 6, 0, "RW", 0, 6'h6, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtMRL_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtMRL_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_RegRet extends uvm_reg;
	rand uvm_reg_field RegRet;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RegRet: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_RegRet");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RegRet = uvm_reg_field::type_id::create("RegRet",,get_full_name());
      this.RegRet.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_RegRet)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_RegRet


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DisableZQupdateOnSnoop extends uvm_reg;
	rand uvm_reg_field DisableZQupdateOnSnoop;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DisableZQupdateOnSnoop: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DisableZQupdateOnSnoop");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DisableZQupdateOnSnoop = uvm_reg_field::type_id::create("DisableZQupdateOnSnoop",,get_full_name());
      this.DisableZQupdateOnSnoop.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DisableZQupdateOnSnoop)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DisableZQupdateOnSnoop


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenModeSel extends uvm_reg;
	rand uvm_reg_field Prbs0GenModeSel;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenModeSel: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenModeSel");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenModeSel = uvm_reg_field::type_id::create("Prbs0GenModeSel",,get_full_name());
      this.Prbs0GenModeSel.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenModeSel)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenModeSel


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenUiMuxSel extends uvm_reg;
	rand uvm_reg_field Prbs0GenUiMuxSel;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenUiMuxSel: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenUiMuxSel");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenUiMuxSel = uvm_reg_field::type_id::create("Prbs0GenUiMuxSel",,get_full_name());
      this.Prbs0GenUiMuxSel.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenUiMuxSel)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenUiMuxSel


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly0 extends uvm_reg;
	rand uvm_reg_field Prbs0GenTapDly0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenTapDly0: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenTapDly0 = uvm_reg_field::type_id::create("Prbs0GenTapDly0",,get_full_name());
      this.Prbs0GenTapDly0.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly1 extends uvm_reg;
	rand uvm_reg_field Prbs0GenTapDly1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenTapDly1: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenTapDly1 = uvm_reg_field::type_id::create("Prbs0GenTapDly1",,get_full_name());
      this.Prbs0GenTapDly1.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly2 extends uvm_reg;
	rand uvm_reg_field Prbs0GenTapDly2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenTapDly2: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly2");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenTapDly2 = uvm_reg_field::type_id::create("Prbs0GenTapDly2",,get_full_name());
      this.Prbs0GenTapDly2.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly2)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly2


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly3 extends uvm_reg;
	rand uvm_reg_field Prbs0GenTapDly3;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenTapDly3: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly3");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenTapDly3 = uvm_reg_field::type_id::create("Prbs0GenTapDly3",,get_full_name());
      this.Prbs0GenTapDly3.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly3)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly3


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly4 extends uvm_reg;
	rand uvm_reg_field Prbs0GenTapDly4;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenTapDly4: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly4");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenTapDly4 = uvm_reg_field::type_id::create("Prbs0GenTapDly4",,get_full_name());
      this.Prbs0GenTapDly4.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly4)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly4


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly5 extends uvm_reg;
	rand uvm_reg_field Prbs0GenTapDly5;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenTapDly5: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly5");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenTapDly5 = uvm_reg_field::type_id::create("Prbs0GenTapDly5",,get_full_name());
      this.Prbs0GenTapDly5.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly5)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly5


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly6 extends uvm_reg;
	rand uvm_reg_field Prbs0GenTapDly6;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenTapDly6: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly6");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenTapDly6 = uvm_reg_field::type_id::create("Prbs0GenTapDly6",,get_full_name());
      this.Prbs0GenTapDly6.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly6)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly6


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly7 extends uvm_reg;
	rand uvm_reg_field Prbs0GenTapDly7;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenTapDly7: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly7");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenTapDly7 = uvm_reg_field::type_id::create("Prbs0GenTapDly7",,get_full_name());
      this.Prbs0GenTapDly7.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly7)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly7


class ral_reg_DWC_DDRPHYA_PPGC0_p0_MtestMuxSel extends uvm_reg;
	rand uvm_reg_field MtestMuxSel;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   MtestMuxSel: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_MtestMuxSel");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.MtestMuxSel = uvm_reg_field::type_id::create("MtestMuxSel",,get_full_name());
      this.MtestMuxSel.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_MtestMuxSel)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_MtestMuxSel


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateLo extends uvm_reg;
	rand uvm_reg_field Prbs0GenStateLo;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenStateLo: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateLo");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenStateLo = uvm_reg_field::type_id::create("Prbs0GenStateLo",,get_full_name());
      this.Prbs0GenStateLo.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateLo)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateLo


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateHi extends uvm_reg;
	rand uvm_reg_field Prbs0GenStateHi;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs0GenStateHi: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateHi");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs0GenStateHi = uvm_reg_field::type_id::create("Prbs0GenStateHi",,get_full_name());
      this.Prbs0GenStateHi.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateHi)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateHi


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenModeSel extends uvm_reg;
	rand uvm_reg_field Prbs1GenModeSel;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenModeSel: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenModeSel");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenModeSel = uvm_reg_field::type_id::create("Prbs1GenModeSel",,get_full_name());
      this.Prbs1GenModeSel.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenModeSel)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenModeSel


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenUiMuxSel extends uvm_reg;
	rand uvm_reg_field Prbs1GenUiMuxSel;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenUiMuxSel: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenUiMuxSel");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenUiMuxSel = uvm_reg_field::type_id::create("Prbs1GenUiMuxSel",,get_full_name());
      this.Prbs1GenUiMuxSel.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenUiMuxSel)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenUiMuxSel


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly0 extends uvm_reg;
	rand uvm_reg_field Prbs1GenTapDly0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenTapDly0: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenTapDly0 = uvm_reg_field::type_id::create("Prbs1GenTapDly0",,get_full_name());
      this.Prbs1GenTapDly0.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly1 extends uvm_reg;
	rand uvm_reg_field Prbs1GenTapDly1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenTapDly1: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenTapDly1 = uvm_reg_field::type_id::create("Prbs1GenTapDly1",,get_full_name());
      this.Prbs1GenTapDly1.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly2 extends uvm_reg;
	rand uvm_reg_field Prbs1GenTapDly2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenTapDly2: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly2");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenTapDly2 = uvm_reg_field::type_id::create("Prbs1GenTapDly2",,get_full_name());
      this.Prbs1GenTapDly2.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly2)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly2


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly3 extends uvm_reg;
	rand uvm_reg_field Prbs1GenTapDly3;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenTapDly3: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly3");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenTapDly3 = uvm_reg_field::type_id::create("Prbs1GenTapDly3",,get_full_name());
      this.Prbs1GenTapDly3.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly3)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly3


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly4 extends uvm_reg;
	rand uvm_reg_field Prbs1GenTapDly4;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenTapDly4: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly4");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenTapDly4 = uvm_reg_field::type_id::create("Prbs1GenTapDly4",,get_full_name());
      this.Prbs1GenTapDly4.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly4)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly4


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly5 extends uvm_reg;
	rand uvm_reg_field Prbs1GenTapDly5;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenTapDly5: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly5");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenTapDly5 = uvm_reg_field::type_id::create("Prbs1GenTapDly5",,get_full_name());
      this.Prbs1GenTapDly5.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly5)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly5


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly6 extends uvm_reg;
	rand uvm_reg_field Prbs1GenTapDly6;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenTapDly6: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly6");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenTapDly6 = uvm_reg_field::type_id::create("Prbs1GenTapDly6",,get_full_name());
      this.Prbs1GenTapDly6.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly6)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly6


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly7 extends uvm_reg;
	rand uvm_reg_field Prbs1GenTapDly7;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenTapDly7: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly7");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenTapDly7 = uvm_reg_field::type_id::create("Prbs1GenTapDly7",,get_full_name());
      this.Prbs1GenTapDly7.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly7)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly7


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateLo extends uvm_reg;
	rand uvm_reg_field Prbs1GenStateLo;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenStateLo: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateLo");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenStateLo = uvm_reg_field::type_id::create("Prbs1GenStateLo",,get_full_name());
      this.Prbs1GenStateLo.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateLo)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateLo


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateHi extends uvm_reg;
	rand uvm_reg_field Prbs1GenStateHi;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs1GenStateHi: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateHi");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs1GenStateHi = uvm_reg_field::type_id::create("Prbs1GenStateHi",,get_full_name());
      this.Prbs1GenStateHi.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateHi)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateHi


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenModeSel extends uvm_reg;
	rand uvm_reg_field Prbs2GenModeSel;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenModeSel: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenModeSel");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenModeSel = uvm_reg_field::type_id::create("Prbs2GenModeSel",,get_full_name());
      this.Prbs2GenModeSel.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenModeSel)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenModeSel


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenUiMuxSel extends uvm_reg;
	rand uvm_reg_field Prbs2GenUiMuxSel;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenUiMuxSel: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenUiMuxSel");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenUiMuxSel = uvm_reg_field::type_id::create("Prbs2GenUiMuxSel",,get_full_name());
      this.Prbs2GenUiMuxSel.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenUiMuxSel)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenUiMuxSel


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly0 extends uvm_reg;
	rand uvm_reg_field Prbs2GenTapDly0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenTapDly0: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenTapDly0 = uvm_reg_field::type_id::create("Prbs2GenTapDly0",,get_full_name());
      this.Prbs2GenTapDly0.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly1 extends uvm_reg;
	rand uvm_reg_field Prbs2GenTapDly1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenTapDly1: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenTapDly1 = uvm_reg_field::type_id::create("Prbs2GenTapDly1",,get_full_name());
      this.Prbs2GenTapDly1.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly2 extends uvm_reg;
	rand uvm_reg_field Prbs2GenTapDly2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenTapDly2: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly2");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenTapDly2 = uvm_reg_field::type_id::create("Prbs2GenTapDly2",,get_full_name());
      this.Prbs2GenTapDly2.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly2)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly2


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly3 extends uvm_reg;
	rand uvm_reg_field Prbs2GenTapDly3;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenTapDly3: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly3");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenTapDly3 = uvm_reg_field::type_id::create("Prbs2GenTapDly3",,get_full_name());
      this.Prbs2GenTapDly3.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly3)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly3


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly4 extends uvm_reg;
	rand uvm_reg_field Prbs2GenTapDly4;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenTapDly4: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly4");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenTapDly4 = uvm_reg_field::type_id::create("Prbs2GenTapDly4",,get_full_name());
      this.Prbs2GenTapDly4.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly4)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly4


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly5 extends uvm_reg;
	rand uvm_reg_field Prbs2GenTapDly5;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenTapDly5: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly5");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenTapDly5 = uvm_reg_field::type_id::create("Prbs2GenTapDly5",,get_full_name());
      this.Prbs2GenTapDly5.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly5)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly5


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly6 extends uvm_reg;
	rand uvm_reg_field Prbs2GenTapDly6;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenTapDly6: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly6");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenTapDly6 = uvm_reg_field::type_id::create("Prbs2GenTapDly6",,get_full_name());
      this.Prbs2GenTapDly6.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly6)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly6


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly7 extends uvm_reg;
	rand uvm_reg_field Prbs2GenTapDly7;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenTapDly7: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly7");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenTapDly7 = uvm_reg_field::type_id::create("Prbs2GenTapDly7",,get_full_name());
      this.Prbs2GenTapDly7.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly7)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly7


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateLo extends uvm_reg;
	rand uvm_reg_field Prbs2GenStateLo;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenStateLo: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateLo");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenStateLo = uvm_reg_field::type_id::create("Prbs2GenStateLo",,get_full_name());
      this.Prbs2GenStateLo.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateLo)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateLo


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateHi extends uvm_reg;
	rand uvm_reg_field Prbs2GenStateHi;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Prbs2GenStateHi: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateHi");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Prbs2GenStateHi = uvm_reg_field::type_id::create("Prbs2GenStateHi",,get_full_name());
      this.Prbs2GenStateHi.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateHi)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateHi


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PPTTrainSetup_p0 extends uvm_reg;
	rand uvm_reg_field PhyMstrTrainInterval;
	rand uvm_reg_field PhyMstrMaxReqToAck;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyMstrTrainInterval: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   PhyMstrMaxReqToAck: coverpoint {m_data[6:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PPTTrainSetup_p0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyMstrTrainInterval = uvm_reg_field::type_id::create("PhyMstrTrainInterval",,get_full_name());
      this.PhyMstrTrainInterval.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 0);
      this.PhyMstrMaxReqToAck = uvm_reg_field::type_id::create("PhyMstrMaxReqToAck",,get_full_name());
      this.PhyMstrMaxReqToAck.configure(this, 3, 4, "RW", 0, 3'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PPTTrainSetup_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PPTTrainSetup_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyMstrFreqOverride_p0 extends uvm_reg;
	rand uvm_reg_field PhyMstrFreqOverride_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyMstrFreqOverride_p0: coverpoint {m_data[4:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyMstrFreqOverride_p0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyMstrFreqOverride_p0 = uvm_reg_field::type_id::create("PhyMstrFreqOverride_p0",,get_full_name());
      this.PhyMstrFreqOverride_p0.configure(this, 5, 0, "RW", 0, 5'h2, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyMstrFreqOverride_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyMstrFreqOverride_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiInitComplete extends uvm_reg;
	rand uvm_reg_field DfiInitComplete;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DfiInitComplete: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiInitComplete");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DfiInitComplete = uvm_reg_field::type_id::create("DfiInitComplete",,get_full_name());
      this.DfiInitComplete.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiInitComplete)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiInitComplete


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCParityInvert extends uvm_reg;
	rand uvm_reg_field PPGCParityInvert;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PPGCParityInvert: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PPGCParityInvert");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PPGCParityInvert = uvm_reg_field::type_id::create("PPGCParityInvert",,get_full_name());
      this.PPGCParityInvert.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCParityInvert)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCParityInvert


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PMIEnable extends uvm_reg;
	rand uvm_reg_field PMIEnable;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PMIEnable: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PMIEnable");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PMIEnable = uvm_reg_field::type_id::create("PMIEnable",,get_full_name());
      this.PMIEnable.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PMIEnable)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PMIEnable


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi0Status extends uvm_reg;
	uvm_reg_field Dfi0Status;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Dfi0Status: coverpoint {m_data[12:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {14'b????????????00};
	      wildcard bins bit_0_wr_as_1 = {14'b????????????10};
	      wildcard bins bit_0_rd = {14'b?????????????1};
	      wildcard bins bit_1_wr_as_0 = {14'b???????????0?0};
	      wildcard bins bit_1_wr_as_1 = {14'b???????????1?0};
	      wildcard bins bit_1_rd = {14'b?????????????1};
	      wildcard bins bit_2_wr_as_0 = {14'b??????????0??0};
	      wildcard bins bit_2_wr_as_1 = {14'b??????????1??0};
	      wildcard bins bit_2_rd = {14'b?????????????1};
	      wildcard bins bit_3_wr_as_0 = {14'b?????????0???0};
	      wildcard bins bit_3_wr_as_1 = {14'b?????????1???0};
	      wildcard bins bit_3_rd = {14'b?????????????1};
	      wildcard bins bit_4_wr_as_0 = {14'b????????0????0};
	      wildcard bins bit_4_wr_as_1 = {14'b????????1????0};
	      wildcard bins bit_4_rd = {14'b?????????????1};
	      wildcard bins bit_5_wr_as_0 = {14'b???????0?????0};
	      wildcard bins bit_5_wr_as_1 = {14'b???????1?????0};
	      wildcard bins bit_5_rd = {14'b?????????????1};
	      wildcard bins bit_6_wr_as_0 = {14'b??????0??????0};
	      wildcard bins bit_6_wr_as_1 = {14'b??????1??????0};
	      wildcard bins bit_6_rd = {14'b?????????????1};
	      wildcard bins bit_7_wr_as_0 = {14'b?????0???????0};
	      wildcard bins bit_7_wr_as_1 = {14'b?????1???????0};
	      wildcard bins bit_7_rd = {14'b?????????????1};
	      wildcard bins bit_8_wr_as_0 = {14'b????0????????0};
	      wildcard bins bit_8_wr_as_1 = {14'b????1????????0};
	      wildcard bins bit_8_rd = {14'b?????????????1};
	      wildcard bins bit_9_wr_as_0 = {14'b???0?????????0};
	      wildcard bins bit_9_wr_as_1 = {14'b???1?????????0};
	      wildcard bins bit_9_rd = {14'b?????????????1};
	      wildcard bins bit_10_wr_as_0 = {14'b??0??????????0};
	      wildcard bins bit_10_wr_as_1 = {14'b??1??????????0};
	      wildcard bins bit_10_rd = {14'b?????????????1};
	      wildcard bins bit_11_wr_as_0 = {14'b?0???????????0};
	      wildcard bins bit_11_wr_as_1 = {14'b?1???????????0};
	      wildcard bins bit_11_rd = {14'b?????????????1};
	      wildcard bins bit_12_wr_as_0 = {14'b0????????????0};
	      wildcard bins bit_12_wr_as_1 = {14'b1????????????0};
	      wildcard bins bit_12_rd = {14'b?????????????1};
	      option.weight = 39;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Dfi0Status");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Dfi0Status = uvm_reg_field::type_id::create("Dfi0Status",,get_full_name());
      this.Dfi0Status.configure(this, 13, 0, "RO", 1, 13'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi0Status)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi0Status


class ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi1Status extends uvm_reg;
	uvm_reg_field Dfi1Status;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Dfi1Status: coverpoint {m_data[12:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {14'b????????????00};
	      wildcard bins bit_0_wr_as_1 = {14'b????????????10};
	      wildcard bins bit_0_rd = {14'b?????????????1};
	      wildcard bins bit_1_wr_as_0 = {14'b???????????0?0};
	      wildcard bins bit_1_wr_as_1 = {14'b???????????1?0};
	      wildcard bins bit_1_rd = {14'b?????????????1};
	      wildcard bins bit_2_wr_as_0 = {14'b??????????0??0};
	      wildcard bins bit_2_wr_as_1 = {14'b??????????1??0};
	      wildcard bins bit_2_rd = {14'b?????????????1};
	      wildcard bins bit_3_wr_as_0 = {14'b?????????0???0};
	      wildcard bins bit_3_wr_as_1 = {14'b?????????1???0};
	      wildcard bins bit_3_rd = {14'b?????????????1};
	      wildcard bins bit_4_wr_as_0 = {14'b????????0????0};
	      wildcard bins bit_4_wr_as_1 = {14'b????????1????0};
	      wildcard bins bit_4_rd = {14'b?????????????1};
	      wildcard bins bit_5_wr_as_0 = {14'b???????0?????0};
	      wildcard bins bit_5_wr_as_1 = {14'b???????1?????0};
	      wildcard bins bit_5_rd = {14'b?????????????1};
	      wildcard bins bit_6_wr_as_0 = {14'b??????0??????0};
	      wildcard bins bit_6_wr_as_1 = {14'b??????1??????0};
	      wildcard bins bit_6_rd = {14'b?????????????1};
	      wildcard bins bit_7_wr_as_0 = {14'b?????0???????0};
	      wildcard bins bit_7_wr_as_1 = {14'b?????1???????0};
	      wildcard bins bit_7_rd = {14'b?????????????1};
	      wildcard bins bit_8_wr_as_0 = {14'b????0????????0};
	      wildcard bins bit_8_wr_as_1 = {14'b????1????????0};
	      wildcard bins bit_8_rd = {14'b?????????????1};
	      wildcard bins bit_9_wr_as_0 = {14'b???0?????????0};
	      wildcard bins bit_9_wr_as_1 = {14'b???1?????????0};
	      wildcard bins bit_9_rd = {14'b?????????????1};
	      wildcard bins bit_10_wr_as_0 = {14'b??0??????????0};
	      wildcard bins bit_10_wr_as_1 = {14'b??1??????????0};
	      wildcard bins bit_10_rd = {14'b?????????????1};
	      wildcard bins bit_11_wr_as_0 = {14'b?0???????????0};
	      wildcard bins bit_11_wr_as_1 = {14'b?1???????????0};
	      wildcard bins bit_11_rd = {14'b?????????????1};
	      wildcard bins bit_12_wr_as_0 = {14'b0????????????0};
	      wildcard bins bit_12_wr_as_1 = {14'b1????????????0};
	      wildcard bins bit_12_rd = {14'b?????????????1};
	      option.weight = 39;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_Dfi1Status");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Dfi1Status = uvm_reg_field::type_id::create("Dfi1Status",,get_full_name());
      this.Dfi1Status.configure(this, 13, 0, "RO", 1, 13'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi1Status)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi1Status


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays0_p0 extends uvm_reg;
	rand uvm_reg_field PhyUpdAckDelay0;
	rand uvm_reg_field PhyUpdReqDelay0;
	rand uvm_reg_field CtrlUpdReqDelay0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyUpdAckDelay0: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   PhyUpdReqDelay0: coverpoint {m_data[7:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   CtrlUpdReqDelay0: coverpoint {m_data[11:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays0_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyUpdAckDelay0 = uvm_reg_field::type_id::create("PhyUpdAckDelay0",,get_full_name());
      this.PhyUpdAckDelay0.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 0);
      this.PhyUpdReqDelay0 = uvm_reg_field::type_id::create("PhyUpdReqDelay0",,get_full_name());
      this.PhyUpdReqDelay0.configure(this, 4, 4, "RW", 0, 4'h0, 1, 0, 0);
      this.CtrlUpdReqDelay0 = uvm_reg_field::type_id::create("CtrlUpdReqDelay0",,get_full_name());
      this.CtrlUpdReqDelay0.configure(this, 4, 8, "RW", 0, 4'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays0_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays0_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD0 extends uvm_reg;
	rand uvm_reg_field DFIPHYUPDCNT0;
	rand uvm_reg_field DFIPHYUPDRESP0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DFIPHYUPDCNT0: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   DFIPHYUPDRESP0: coverpoint {m_data[6:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DFIPHYUPDCNT0 = uvm_reg_field::type_id::create("DFIPHYUPDCNT0",,get_full_name());
      this.DFIPHYUPDCNT0.configure(this, 4, 0, "RW", 0, 4'h7, 1, 0, 0);
      this.DFIPHYUPDRESP0 = uvm_reg_field::type_id::create("DFIPHYUPDRESP0",,get_full_name());
      this.DFIPHYUPDRESP0.configure(this, 3, 4, "RW", 0, 3'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn0 extends uvm_reg;
	rand uvm_reg_field DfiLpCtrlEn0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DfiLpCtrlEn0: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DfiLpCtrlEn0 = uvm_reg_field::type_id::create("DfiLpCtrlEn0",,get_full_name());
      this.DfiLpCtrlEn0.configure(this, 1, 0, "RW", 0, 1'h1, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn0 extends uvm_reg;
	rand uvm_reg_field DfiLpDataEn0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DfiLpDataEn0: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DfiLpDataEn0 = uvm_reg_field::type_id::create("DfiLpDataEn0",,get_full_name());
      this.DfiLpDataEn0.configure(this, 1, 0, "RW", 0, 1'h1, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl0 extends uvm_reg;
	rand uvm_reg_field DbyteDynOdtEn0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DbyteDynOdtEn0: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DbyteDynOdtEn0 = uvm_reg_field::type_id::create("DbyteDynOdtEn0",,get_full_name());
      this.DbyteDynOdtEn0.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays0_p0 extends uvm_reg;
	rand uvm_reg_field LpCtrlAckDelay0;
	rand uvm_reg_field LpDataAckDelay0;
	rand uvm_reg_field CtrlUpdAckDelay0;
	rand uvm_reg_field LpAssertAckDelay0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   LpCtrlAckDelay0: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   LpDataAckDelay0: coverpoint {m_data[7:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   CtrlUpdAckDelay0: coverpoint {m_data[11:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   LpAssertAckDelay0: coverpoint {m_data[15:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays0_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.LpCtrlAckDelay0 = uvm_reg_field::type_id::create("LpCtrlAckDelay0",,get_full_name());
      this.LpCtrlAckDelay0.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 0);
      this.LpDataAckDelay0 = uvm_reg_field::type_id::create("LpDataAckDelay0",,get_full_name());
      this.LpDataAckDelay0.configure(this, 4, 4, "RW", 0, 4'h0, 1, 0, 0);
      this.CtrlUpdAckDelay0 = uvm_reg_field::type_id::create("CtrlUpdAckDelay0",,get_full_name());
      this.CtrlUpdAckDelay0.configure(this, 4, 8, "RW", 0, 4'h0, 1, 0, 0);
      this.LpAssertAckDelay0 = uvm_reg_field::type_id::create("LpAssertAckDelay0",,get_full_name());
      this.LpAssertAckDelay0.configure(this, 4, 12, "RW", 0, 4'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays0_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays0_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnA extends uvm_reg;
	rand uvm_reg_field HwtLpCsEnA;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   HwtLpCsEnA: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnA");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.HwtLpCsEnA = uvm_reg_field::type_id::create("HwtLpCsEnA",,get_full_name());
      this.HwtLpCsEnA.configure(this, 2, 0, "RW", 0, 2'h3, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnA)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnA


class ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnB extends uvm_reg;
	rand uvm_reg_field HwtLpCsEnB;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   HwtLpCsEnB: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnB");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.HwtLpCsEnB = uvm_reg_field::type_id::create("HwtLpCsEnB",,get_full_name());
      this.HwtLpCsEnB.configure(this, 2, 0, "RW", 0, 2'h3, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnB)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnB


class ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtCtrl extends uvm_reg;
	rand uvm_reg_field HwtCtrl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   HwtCtrl: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_HwtCtrl");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.HwtCtrl = uvm_reg_field::type_id::create("HwtCtrl",,get_full_name());
      this.HwtCtrl.configure(this, 1, 0, "RW", 0, 1'h1, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtCtrl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtCtrl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlOvr extends uvm_reg;
	rand uvm_reg_field HwtControlOvr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   HwtControlOvr: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_HwtControlOvr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.HwtControlOvr = uvm_reg_field::type_id::create("HwtControlOvr",,get_full_name());
      this.HwtControlOvr.configure(this, 12, 0, "RW", 0, 12'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlOvr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlOvr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ScratchPadPPGC extends uvm_reg;
	rand uvm_reg_field ScratchPadPPGC;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ScratchPadPPGC: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ScratchPadPPGC");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ScratchPadPPGC = uvm_reg_field::type_id::create("ScratchPadPPGC",,get_full_name());
      this.ScratchPadPPGC.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ScratchPadPPGC)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ScratchPadPPGC


class ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlVal extends uvm_reg;
	rand uvm_reg_field HwtControlVal;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   HwtControlVal: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_HwtControlVal");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.HwtControlVal = uvm_reg_field::type_id::create("HwtControlVal",,get_full_name());
      this.HwtControlVal.configure(this, 12, 0, "RW", 0, 12'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlVal)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlVal


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ForceHWTClkGaterEnables extends uvm_reg;
	rand uvm_reg_field ForceACSMClkEnHigh;
	rand uvm_reg_field ForceACSMClkEnLow;
	rand uvm_reg_field ForcePIEClkEnHigh;
	rand uvm_reg_field ForcePIEClkEnLow;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ForceACSMClkEnHigh: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ForceACSMClkEnLow: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ForcePIEClkEnHigh: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ForcePIEClkEnLow: coverpoint {m_data[3:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ForceHWTClkGaterEnables");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ForceACSMClkEnHigh = uvm_reg_field::type_id::create("ForceACSMClkEnHigh",,get_full_name());
      this.ForceACSMClkEnHigh.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.ForceACSMClkEnLow = uvm_reg_field::type_id::create("ForceACSMClkEnLow",,get_full_name());
      this.ForceACSMClkEnLow.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.ForcePIEClkEnHigh = uvm_reg_field::type_id::create("ForcePIEClkEnHigh",,get_full_name());
      this.ForcePIEClkEnHigh.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
      this.ForcePIEClkEnLow = uvm_reg_field::type_id::create("ForcePIEClkEnLow",,get_full_name());
      this.ForcePIEClkEnLow.configure(this, 1, 3, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ForceHWTClkGaterEnables)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ForceHWTClkGaterEnables


class ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdGoodCtr extends uvm_reg;
	uvm_reg_field MasUpdGoodCtr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   MasUpdGoodCtr: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd = {17'b????????????????1};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd = {17'b????????????????1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd = {17'b????????????????1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd = {17'b????????????????1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd = {17'b????????????????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd = {17'b????????????????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd = {17'b????????????????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd = {17'b????????????????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd = {17'b????????????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd = {17'b????????????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd = {17'b????????????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd = {17'b????????????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd = {17'b????????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd = {17'b????????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd = {17'b????????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd = {17'b????????????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_MasUpdGoodCtr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.MasUpdGoodCtr = uvm_reg_field::type_id::create("MasUpdGoodCtr",,get_full_name());
      this.MasUpdGoodCtr.configure(this, 16, 0, "RO", 1, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdGoodCtr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdGoodCtr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0GoodCtr extends uvm_reg;
	uvm_reg_field PhyUpd0GoodCtr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyUpd0GoodCtr: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd = {17'b????????????????1};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd = {17'b????????????????1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd = {17'b????????????????1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd = {17'b????????????????1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd = {17'b????????????????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd = {17'b????????????????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd = {17'b????????????????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd = {17'b????????????????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd = {17'b????????????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd = {17'b????????????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd = {17'b????????????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd = {17'b????????????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd = {17'b????????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd = {17'b????????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd = {17'b????????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd = {17'b????????????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyUpd0GoodCtr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyUpd0GoodCtr = uvm_reg_field::type_id::create("PhyUpd0GoodCtr",,get_full_name());
      this.PhyUpd0GoodCtr.configure(this, 16, 0, "RO", 1, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0GoodCtr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0GoodCtr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1GoodCtr extends uvm_reg;
	uvm_reg_field PhyUpd1GoodCtr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyUpd1GoodCtr: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd = {17'b????????????????1};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd = {17'b????????????????1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd = {17'b????????????????1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd = {17'b????????????????1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd = {17'b????????????????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd = {17'b????????????????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd = {17'b????????????????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd = {17'b????????????????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd = {17'b????????????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd = {17'b????????????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd = {17'b????????????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd = {17'b????????????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd = {17'b????????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd = {17'b????????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd = {17'b????????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd = {17'b????????????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyUpd1GoodCtr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyUpd1GoodCtr = uvm_reg_field::type_id::create("PhyUpd1GoodCtr",,get_full_name());
      this.PhyUpd1GoodCtr.configure(this, 16, 0, "RO", 1, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1GoodCtr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1GoodCtr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd0GoodCtr extends uvm_reg;
	uvm_reg_field CtlUpd0GoodCtr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   CtlUpd0GoodCtr: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd = {17'b????????????????1};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd = {17'b????????????????1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd = {17'b????????????????1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd = {17'b????????????????1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd = {17'b????????????????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd = {17'b????????????????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd = {17'b????????????????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd = {17'b????????????????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd = {17'b????????????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd = {17'b????????????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd = {17'b????????????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd = {17'b????????????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd = {17'b????????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd = {17'b????????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd = {17'b????????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd = {17'b????????????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_CtlUpd0GoodCtr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.CtlUpd0GoodCtr = uvm_reg_field::type_id::create("CtlUpd0GoodCtr",,get_full_name());
      this.CtlUpd0GoodCtr.configure(this, 16, 0, "RO", 1, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd0GoodCtr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd0GoodCtr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd1GoodCtr extends uvm_reg;
	uvm_reg_field CtlUpd1GoodCtr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   CtlUpd1GoodCtr: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd = {17'b????????????????1};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd = {17'b????????????????1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd = {17'b????????????????1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd = {17'b????????????????1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd = {17'b????????????????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd = {17'b????????????????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd = {17'b????????????????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd = {17'b????????????????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd = {17'b????????????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd = {17'b????????????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd = {17'b????????????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd = {17'b????????????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd = {17'b????????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd = {17'b????????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd = {17'b????????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd = {17'b????????????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_CtlUpd1GoodCtr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.CtlUpd1GoodCtr = uvm_reg_field::type_id::create("CtlUpd1GoodCtr",,get_full_name());
      this.CtlUpd1GoodCtr.configure(this, 16, 0, "RO", 1, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd1GoodCtr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd1GoodCtr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdFailCtr extends uvm_reg;
	uvm_reg_field MasUpdFailCtr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   MasUpdFailCtr: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd = {17'b????????????????1};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd = {17'b????????????????1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd = {17'b????????????????1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd = {17'b????????????????1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd = {17'b????????????????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd = {17'b????????????????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd = {17'b????????????????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd = {17'b????????????????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd = {17'b????????????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd = {17'b????????????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd = {17'b????????????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd = {17'b????????????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd = {17'b????????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd = {17'b????????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd = {17'b????????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd = {17'b????????????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_MasUpdFailCtr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.MasUpdFailCtr = uvm_reg_field::type_id::create("MasUpdFailCtr",,get_full_name());
      this.MasUpdFailCtr.configure(this, 16, 0, "RO", 1, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdFailCtr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdFailCtr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0FailCtr extends uvm_reg;
	uvm_reg_field PhyUpd0FailCtr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyUpd0FailCtr: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd = {17'b????????????????1};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd = {17'b????????????????1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd = {17'b????????????????1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd = {17'b????????????????1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd = {17'b????????????????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd = {17'b????????????????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd = {17'b????????????????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd = {17'b????????????????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd = {17'b????????????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd = {17'b????????????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd = {17'b????????????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd = {17'b????????????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd = {17'b????????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd = {17'b????????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd = {17'b????????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd = {17'b????????????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyUpd0FailCtr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyUpd0FailCtr = uvm_reg_field::type_id::create("PhyUpd0FailCtr",,get_full_name());
      this.PhyUpd0FailCtr.configure(this, 16, 0, "RO", 1, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0FailCtr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0FailCtr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1FailCtr extends uvm_reg;
	uvm_reg_field PhyUpd1FailCtr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyUpd1FailCtr: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd = {17'b????????????????1};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd = {17'b????????????????1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd = {17'b????????????????1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd = {17'b????????????????1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd = {17'b????????????????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd = {17'b????????????????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd = {17'b????????????????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd = {17'b????????????????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd = {17'b????????????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd = {17'b????????????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd = {17'b????????????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd = {17'b????????????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd = {17'b????????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd = {17'b????????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd = {17'b????????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd = {17'b????????????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyUpd1FailCtr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyUpd1FailCtr = uvm_reg_field::type_id::create("PhyUpd1FailCtr",,get_full_name());
      this.PhyUpd1FailCtr.configure(this, 16, 0, "RO", 1, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1FailCtr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1FailCtr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyPerfCtrEnable extends uvm_reg;
	rand uvm_reg_field MasUpdGoodCtl;
	rand uvm_reg_field PhyUpd0GoodCtl;
	rand uvm_reg_field PhyUpd1GoodCtl;
	rand uvm_reg_field CtlUpd0GoodCtl;
	rand uvm_reg_field CtlUpd1GoodCtl;
	rand uvm_reg_field MasUpdFailCtl;
	rand uvm_reg_field PhyUpd0FailCtl;
	rand uvm_reg_field PhyUpd1FailCtl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   MasUpdGoodCtl: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyUpd0GoodCtl: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyUpd1GoodCtl: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   CtlUpd0GoodCtl: coverpoint {m_data[3:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   CtlUpd1GoodCtl: coverpoint {m_data[4:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   MasUpdFailCtl: coverpoint {m_data[5:5], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyUpd0FailCtl: coverpoint {m_data[6:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyUpd1FailCtl: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyPerfCtrEnable");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.MasUpdGoodCtl = uvm_reg_field::type_id::create("MasUpdGoodCtl",,get_full_name());
      this.MasUpdGoodCtl.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyUpd0GoodCtl = uvm_reg_field::type_id::create("PhyUpd0GoodCtl",,get_full_name());
      this.PhyUpd0GoodCtl.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyUpd1GoodCtl = uvm_reg_field::type_id::create("PhyUpd1GoodCtl",,get_full_name());
      this.PhyUpd1GoodCtl.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
      this.CtlUpd0GoodCtl = uvm_reg_field::type_id::create("CtlUpd0GoodCtl",,get_full_name());
      this.CtlUpd0GoodCtl.configure(this, 1, 3, "RW", 0, 1'h0, 1, 0, 0);
      this.CtlUpd1GoodCtl = uvm_reg_field::type_id::create("CtlUpd1GoodCtl",,get_full_name());
      this.CtlUpd1GoodCtl.configure(this, 1, 4, "RW", 0, 1'h0, 1, 0, 0);
      this.MasUpdFailCtl = uvm_reg_field::type_id::create("MasUpdFailCtl",,get_full_name());
      this.MasUpdFailCtl.configure(this, 1, 5, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyUpd0FailCtl = uvm_reg_field::type_id::create("PhyUpd0FailCtl",,get_full_name());
      this.PhyUpd0FailCtl.configure(this, 1, 6, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyUpd1FailCtl = uvm_reg_field::type_id::create("PhyUpd1FailCtl",,get_full_name());
      this.PhyUpd1FailCtl.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyPerfCtrEnable)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyPerfCtrEnable


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays1_p0 extends uvm_reg;
	rand uvm_reg_field PhyUpdAckDelay1;
	rand uvm_reg_field PhyUpdReqDelay1;
	rand uvm_reg_field CtrlUpdReqDelay1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyUpdAckDelay1: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   PhyUpdReqDelay1: coverpoint {m_data[7:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   CtrlUpdReqDelay1: coverpoint {m_data[11:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays1_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyUpdAckDelay1 = uvm_reg_field::type_id::create("PhyUpdAckDelay1",,get_full_name());
      this.PhyUpdAckDelay1.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 0);
      this.PhyUpdReqDelay1 = uvm_reg_field::type_id::create("PhyUpdReqDelay1",,get_full_name());
      this.PhyUpdReqDelay1.configure(this, 4, 4, "RW", 0, 4'h0, 1, 0, 0);
      this.CtrlUpdReqDelay1 = uvm_reg_field::type_id::create("CtrlUpdReqDelay1",,get_full_name());
      this.CtrlUpdReqDelay1.configure(this, 4, 8, "RW", 0, 4'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays1_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays1_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD1 extends uvm_reg;
	rand uvm_reg_field DFIPHYUPDCNT1;
	rand uvm_reg_field DFIPHYUPDRESP1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DFIPHYUPDCNT1: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   DFIPHYUPDRESP1: coverpoint {m_data[6:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DFIPHYUPDCNT1 = uvm_reg_field::type_id::create("DFIPHYUPDCNT1",,get_full_name());
      this.DFIPHYUPDCNT1.configure(this, 4, 0, "RW", 0, 4'h7, 1, 0, 0);
      this.DFIPHYUPDRESP1 = uvm_reg_field::type_id::create("DFIPHYUPDRESP1",,get_full_name());
      this.DFIPHYUPDRESP1.configure(this, 3, 4, "RW", 0, 3'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn1 extends uvm_reg;
	rand uvm_reg_field DfiLpCtrlEn1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DfiLpCtrlEn1: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DfiLpCtrlEn1 = uvm_reg_field::type_id::create("DfiLpCtrlEn1",,get_full_name());
      this.DfiLpCtrlEn1.configure(this, 1, 0, "RW", 0, 1'h1, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn1 extends uvm_reg;
	rand uvm_reg_field DfiLpDataEn1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DfiLpDataEn1: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DfiLpDataEn1 = uvm_reg_field::type_id::create("DfiLpDataEn1",,get_full_name());
      this.DfiLpDataEn1.configure(this, 1, 0, "RW", 0, 1'h1, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl1 extends uvm_reg;
	rand uvm_reg_field DbyteDynOdtEn1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DbyteDynOdtEn1: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DbyteDynOdtEn1 = uvm_reg_field::type_id::create("DbyteDynOdtEn1",,get_full_name());
      this.DbyteDynOdtEn1.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays1_p0 extends uvm_reg;
	rand uvm_reg_field LpCtrlAckDelay1;
	rand uvm_reg_field LpDataAckDelay1;
	rand uvm_reg_field CtrlUpdAckDelay1;
	rand uvm_reg_field LpAssertAckDelay1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   LpCtrlAckDelay1: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   LpDataAckDelay1: coverpoint {m_data[7:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   CtrlUpdAckDelay1: coverpoint {m_data[11:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   LpAssertAckDelay1: coverpoint {m_data[15:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays1_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.LpCtrlAckDelay1 = uvm_reg_field::type_id::create("LpCtrlAckDelay1",,get_full_name());
      this.LpCtrlAckDelay1.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 0);
      this.LpDataAckDelay1 = uvm_reg_field::type_id::create("LpDataAckDelay1",,get_full_name());
      this.LpDataAckDelay1.configure(this, 4, 4, "RW", 0, 4'h0, 1, 0, 0);
      this.CtrlUpdAckDelay1 = uvm_reg_field::type_id::create("CtrlUpdAckDelay1",,get_full_name());
      this.CtrlUpdAckDelay1.configure(this, 4, 8, "RW", 0, 4'h0, 1, 0, 0);
      this.LpAssertAckDelay1 = uvm_reg_field::type_id::create("LpAssertAckDelay1",,get_full_name());
      this.LpAssertAckDelay1.configure(this, 4, 12, "RW", 0, 4'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays1_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays1_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_FspSkipList extends uvm_reg;
	rand uvm_reg_field FspPStateSkip0;
	rand uvm_reg_field FspPStateSkip1;
	rand uvm_reg_field FspPStateSkip2;
	rand uvm_reg_field FspPStateSkip3;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   FspPStateSkip0: coverpoint {m_data[2:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	   FspPStateSkip1: coverpoint {m_data[5:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	   FspPStateSkip2: coverpoint {m_data[8:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	   FspPStateSkip3: coverpoint {m_data[11:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_FspSkipList");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.FspPStateSkip0 = uvm_reg_field::type_id::create("FspPStateSkip0",,get_full_name());
      this.FspPStateSkip0.configure(this, 3, 0, "RW", 0, 3'h0, 1, 0, 0);
      this.FspPStateSkip1 = uvm_reg_field::type_id::create("FspPStateSkip1",,get_full_name());
      this.FspPStateSkip1.configure(this, 3, 3, "RW", 0, 3'h0, 1, 0, 0);
      this.FspPStateSkip2 = uvm_reg_field::type_id::create("FspPStateSkip2",,get_full_name());
      this.FspPStateSkip2.configure(this, 3, 6, "RW", 0, 3'h0, 1, 0, 0);
      this.FspPStateSkip3 = uvm_reg_field::type_id::create("FspPStateSkip3",,get_full_name());
      this.FspPStateSkip3.configure(this, 3, 9, "RW", 0, 3'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_FspSkipList)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_FspSkipList


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCReserved0 extends uvm_reg;
	rand uvm_reg_field PPGCReserved0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PPGCReserved0: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PPGCReserved0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PPGCReserved0 = uvm_reg_field::type_id::create("PPGCReserved0",,get_full_name());
      this.PPGCReserved0.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCReserved0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCReserved0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PUBReservedP1_p0 extends uvm_reg;
	rand uvm_reg_field PUBReservedP1_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PUBReservedP1_p0: coverpoint {m_data[7:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd_as_0 = {9'b???????01};
	      wildcard bins bit_0_rd_as_1 = {9'b???????11};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd_as_0 = {9'b??????0?1};
	      wildcard bins bit_1_rd_as_1 = {9'b??????1?1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd_as_0 = {9'b?????0??1};
	      wildcard bins bit_2_rd_as_1 = {9'b?????1??1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd_as_0 = {9'b????0???1};
	      wildcard bins bit_3_rd_as_1 = {9'b????1???1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd_as_0 = {9'b???0????1};
	      wildcard bins bit_4_rd_as_1 = {9'b???1????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd_as_0 = {9'b??0?????1};
	      wildcard bins bit_5_rd_as_1 = {9'b??1?????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd_as_0 = {9'b?0??????1};
	      wildcard bins bit_6_rd_as_1 = {9'b?1??????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd_as_0 = {9'b0???????1};
	      wildcard bins bit_7_rd_as_1 = {9'b1???????1};
	      option.weight = 32;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PUBReservedP1_p0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PUBReservedP1_p0 = uvm_reg_field::type_id::create("PUBReservedP1_p0",,get_full_name());
      this.PUBReservedP1_p0.configure(this, 8, 0, "RW", 0, 8'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PUBReservedP1_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PUBReservedP1_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptOverride extends uvm_reg;
	rand uvm_reg_field PhyInterruptOverride;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyInterruptOverride: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyInterruptOverride");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyInterruptOverride = uvm_reg_field::type_id::create("PhyInterruptOverride",,get_full_name());
      this.PhyInterruptOverride.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptOverride)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptOverride


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptEnable extends uvm_reg;
	rand uvm_reg_field PhyTrngCmpltEn;
	rand uvm_reg_field PhyInitCmpltEn;
	rand uvm_reg_field PhyTrngFailEn;
	rand uvm_reg_field PhyFWReservedEn;
	rand uvm_reg_field PhyAcsmParityErrEn;
	rand uvm_reg_field PhyPIEParityErrEn;
	rand uvm_reg_field PhyRdfPtrChkErrEn;
	rand uvm_reg_field PhyEccEn;
	rand uvm_reg_field PhyPIEProgErrEn;
	rand uvm_reg_field PhyHWReservedEn;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyTrngCmpltEn: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyInitCmpltEn: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyTrngFailEn: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyFWReservedEn: coverpoint {m_data[7:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	   PhyAcsmParityErrEn: coverpoint {m_data[8:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyPIEParityErrEn: coverpoint {m_data[9:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyRdfPtrChkErrEn: coverpoint {m_data[10:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyEccEn: coverpoint {m_data[11:11], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyPIEProgErrEn: coverpoint {m_data[12:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyHWReservedEn: coverpoint {m_data[15:13], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyInterruptEnable");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyTrngCmpltEn = uvm_reg_field::type_id::create("PhyTrngCmpltEn",,get_full_name());
      this.PhyTrngCmpltEn.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyInitCmpltEn = uvm_reg_field::type_id::create("PhyInitCmpltEn",,get_full_name());
      this.PhyInitCmpltEn.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyTrngFailEn = uvm_reg_field::type_id::create("PhyTrngFailEn",,get_full_name());
      this.PhyTrngFailEn.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyFWReservedEn = uvm_reg_field::type_id::create("PhyFWReservedEn",,get_full_name());
      this.PhyFWReservedEn.configure(this, 5, 3, "RW", 0, 5'h0, 1, 0, 0);
      this.PhyAcsmParityErrEn = uvm_reg_field::type_id::create("PhyAcsmParityErrEn",,get_full_name());
      this.PhyAcsmParityErrEn.configure(this, 1, 8, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyPIEParityErrEn = uvm_reg_field::type_id::create("PhyPIEParityErrEn",,get_full_name());
      this.PhyPIEParityErrEn.configure(this, 1, 9, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyRdfPtrChkErrEn = uvm_reg_field::type_id::create("PhyRdfPtrChkErrEn",,get_full_name());
      this.PhyRdfPtrChkErrEn.configure(this, 1, 10, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyEccEn = uvm_reg_field::type_id::create("PhyEccEn",,get_full_name());
      this.PhyEccEn.configure(this, 1, 11, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyPIEProgErrEn = uvm_reg_field::type_id::create("PhyPIEProgErrEn",,get_full_name());
      this.PhyPIEProgErrEn.configure(this, 1, 12, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyHWReservedEn = uvm_reg_field::type_id::create("PhyHWReservedEn",,get_full_name());
      this.PhyHWReservedEn.configure(this, 3, 13, "RW", 0, 3'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptEnable)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptEnable


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptFWControl extends uvm_reg;
	rand uvm_reg_field PhyTrngCmpltFW;
	rand uvm_reg_field PhyInitCmpltFW;
	rand uvm_reg_field PhyTrngFailFW;
	rand uvm_reg_field PhyFWReservedFW;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyTrngCmpltFW: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyInitCmpltFW: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyTrngFailFW: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyFWReservedFW: coverpoint {m_data[7:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyInterruptFWControl");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyTrngCmpltFW = uvm_reg_field::type_id::create("PhyTrngCmpltFW",,get_full_name());
      this.PhyTrngCmpltFW.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyInitCmpltFW = uvm_reg_field::type_id::create("PhyInitCmpltFW",,get_full_name());
      this.PhyInitCmpltFW.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyTrngFailFW = uvm_reg_field::type_id::create("PhyTrngFailFW",,get_full_name());
      this.PhyTrngFailFW.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyFWReservedFW = uvm_reg_field::type_id::create("PhyFWReservedFW",,get_full_name());
      this.PhyFWReservedFW.configure(this, 5, 3, "RW", 0, 5'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptFWControl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptFWControl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptMask extends uvm_reg;
	rand uvm_reg_field PhyTrngCmpltMsk;
	rand uvm_reg_field PhyInitCmpltMsk;
	rand uvm_reg_field PhyTrngFailMsk;
	rand uvm_reg_field PhyFWReservedMsk;
	rand uvm_reg_field PhyAcsmParityErrMsk;
	rand uvm_reg_field PhyPIEParityErrMsk;
	rand uvm_reg_field PhyRdfPtrChkErrMsk;
	rand uvm_reg_field PhyEccMsk;
	rand uvm_reg_field PhyPIEProgErrMsk;
	rand uvm_reg_field PhyHWReservedMsk;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyTrngCmpltMsk: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyInitCmpltMsk: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyTrngFailMsk: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyFWReservedMsk: coverpoint {m_data[7:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	   PhyAcsmParityErrMsk: coverpoint {m_data[8:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyPIEParityErrMsk: coverpoint {m_data[9:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyRdfPtrChkErrMsk: coverpoint {m_data[10:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyEccMsk: coverpoint {m_data[11:11], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyPIEProgErrMsk: coverpoint {m_data[12:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyHWReservedMsk: coverpoint {m_data[15:13], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyInterruptMask");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyTrngCmpltMsk = uvm_reg_field::type_id::create("PhyTrngCmpltMsk",,get_full_name());
      this.PhyTrngCmpltMsk.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyInitCmpltMsk = uvm_reg_field::type_id::create("PhyInitCmpltMsk",,get_full_name());
      this.PhyInitCmpltMsk.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyTrngFailMsk = uvm_reg_field::type_id::create("PhyTrngFailMsk",,get_full_name());
      this.PhyTrngFailMsk.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyFWReservedMsk = uvm_reg_field::type_id::create("PhyFWReservedMsk",,get_full_name());
      this.PhyFWReservedMsk.configure(this, 5, 3, "RW", 0, 5'h0, 1, 0, 0);
      this.PhyAcsmParityErrMsk = uvm_reg_field::type_id::create("PhyAcsmParityErrMsk",,get_full_name());
      this.PhyAcsmParityErrMsk.configure(this, 1, 8, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyPIEParityErrMsk = uvm_reg_field::type_id::create("PhyPIEParityErrMsk",,get_full_name());
      this.PhyPIEParityErrMsk.configure(this, 1, 9, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyRdfPtrChkErrMsk = uvm_reg_field::type_id::create("PhyRdfPtrChkErrMsk",,get_full_name());
      this.PhyRdfPtrChkErrMsk.configure(this, 1, 10, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyEccMsk = uvm_reg_field::type_id::create("PhyEccMsk",,get_full_name());
      this.PhyEccMsk.configure(this, 1, 11, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyPIEProgErrMsk = uvm_reg_field::type_id::create("PhyPIEProgErrMsk",,get_full_name());
      this.PhyPIEProgErrMsk.configure(this, 1, 12, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyHWReservedMsk = uvm_reg_field::type_id::create("PhyHWReservedMsk",,get_full_name());
      this.PhyHWReservedMsk.configure(this, 3, 13, "RW", 0, 3'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptMask)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptMask


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptClear extends uvm_reg;
	rand uvm_reg_field PhyTrngCmpltClr;
	rand uvm_reg_field PhyInitCmpltClr;
	rand uvm_reg_field PhyTrngFailClr;
	rand uvm_reg_field PhyFWReservedClr;
	rand uvm_reg_field PhyAcsmParityErrClr;
	rand uvm_reg_field PhyPIEParityErrClr;
	rand uvm_reg_field PhyRdfPtrChkErrClr;
	rand uvm_reg_field PhyEccClr;
	rand uvm_reg_field PhyPIEProgErrClr;
	rand uvm_reg_field PhyHWReservedClr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyTrngCmpltClr: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyInitCmpltClr: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyTrngFailClr: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyFWReservedClr: coverpoint {m_data[7:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	   PhyAcsmParityErrClr: coverpoint {m_data[8:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyPIEParityErrClr: coverpoint {m_data[9:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyRdfPtrChkErrClr: coverpoint {m_data[10:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyEccClr: coverpoint {m_data[11:11], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyPIEProgErrClr: coverpoint {m_data[12:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PhyHWReservedClr: coverpoint {m_data[15:13], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyInterruptClear");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyTrngCmpltClr = uvm_reg_field::type_id::create("PhyTrngCmpltClr",,get_full_name());
      this.PhyTrngCmpltClr.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyInitCmpltClr = uvm_reg_field::type_id::create("PhyInitCmpltClr",,get_full_name());
      this.PhyInitCmpltClr.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyTrngFailClr = uvm_reg_field::type_id::create("PhyTrngFailClr",,get_full_name());
      this.PhyTrngFailClr.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyFWReservedClr = uvm_reg_field::type_id::create("PhyFWReservedClr",,get_full_name());
      this.PhyFWReservedClr.configure(this, 5, 3, "RW", 0, 5'h0, 1, 0, 0);
      this.PhyAcsmParityErrClr = uvm_reg_field::type_id::create("PhyAcsmParityErrClr",,get_full_name());
      this.PhyAcsmParityErrClr.configure(this, 1, 8, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyPIEParityErrClr = uvm_reg_field::type_id::create("PhyPIEParityErrClr",,get_full_name());
      this.PhyPIEParityErrClr.configure(this, 1, 9, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyRdfPtrChkErrClr = uvm_reg_field::type_id::create("PhyRdfPtrChkErrClr",,get_full_name());
      this.PhyRdfPtrChkErrClr.configure(this, 1, 10, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyEccClr = uvm_reg_field::type_id::create("PhyEccClr",,get_full_name());
      this.PhyEccClr.configure(this, 1, 11, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyPIEProgErrClr = uvm_reg_field::type_id::create("PhyPIEProgErrClr",,get_full_name());
      this.PhyPIEProgErrClr.configure(this, 1, 12, "RW", 0, 1'h0, 1, 0, 0);
      this.PhyHWReservedClr = uvm_reg_field::type_id::create("PhyHWReservedClr",,get_full_name());
      this.PhyHWReservedClr.configure(this, 3, 13, "RW", 0, 3'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptClear)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptClear


class ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptStatus extends uvm_reg;
	uvm_reg_field PhyTrngCmplt;
	uvm_reg_field PhyInitCmplt;
	uvm_reg_field PhyTrngFail;
	uvm_reg_field PhyFWReserved;
	uvm_reg_field PhyAcsmParityErr;
	uvm_reg_field PhyPIEParityErr;
	uvm_reg_field PhyRdfPtrChkErr;
	uvm_reg_field PhyEccErr;
	uvm_reg_field PhyPIEProgErr;
	uvm_reg_field PhyHWReserved;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PhyTrngCmplt: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   PhyInitCmplt: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   PhyTrngFail: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   PhyFWReserved: coverpoint {m_data[7:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd = {6'b?????1};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd = {6'b?????1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd = {6'b?????1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd = {6'b?????1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd = {6'b?????1};
	      option.weight = 15;
	   }
	   PhyAcsmParityErr: coverpoint {m_data[8:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   PhyPIEParityErr: coverpoint {m_data[9:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   PhyRdfPtrChkErr: coverpoint {m_data[10:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   PhyEccErr: coverpoint {m_data[11:11], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   PhyPIEProgErr: coverpoint {m_data[12:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   PhyHWReserved: coverpoint {m_data[15:13], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd = {4'b???1};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd = {4'b???1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd = {4'b???1};
	      option.weight = 9;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_PhyInterruptStatus");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PhyTrngCmplt = uvm_reg_field::type_id::create("PhyTrngCmplt",,get_full_name());
      this.PhyTrngCmplt.configure(this, 1, 0, "RO", 1, 1'h0, 1, 0, 0);
      this.PhyInitCmplt = uvm_reg_field::type_id::create("PhyInitCmplt",,get_full_name());
      this.PhyInitCmplt.configure(this, 1, 1, "RO", 1, 1'h0, 1, 0, 0);
      this.PhyTrngFail = uvm_reg_field::type_id::create("PhyTrngFail",,get_full_name());
      this.PhyTrngFail.configure(this, 1, 2, "RO", 1, 1'h0, 1, 0, 0);
      this.PhyFWReserved = uvm_reg_field::type_id::create("PhyFWReserved",,get_full_name());
      this.PhyFWReserved.configure(this, 5, 3, "RO", 1, 5'h0, 1, 0, 0);
      this.PhyAcsmParityErr = uvm_reg_field::type_id::create("PhyAcsmParityErr",,get_full_name());
      this.PhyAcsmParityErr.configure(this, 1, 8, "RO", 1, 1'h0, 1, 0, 0);
      this.PhyPIEParityErr = uvm_reg_field::type_id::create("PhyPIEParityErr",,get_full_name());
      this.PhyPIEParityErr.configure(this, 1, 9, "RO", 1, 1'h0, 1, 0, 0);
      this.PhyRdfPtrChkErr = uvm_reg_field::type_id::create("PhyRdfPtrChkErr",,get_full_name());
      this.PhyRdfPtrChkErr.configure(this, 1, 10, "RO", 1, 1'h0, 1, 0, 0);
      this.PhyEccErr = uvm_reg_field::type_id::create("PhyEccErr",,get_full_name());
      this.PhyEccErr.configure(this, 1, 11, "RO", 1, 1'h0, 1, 0, 0);
      this.PhyPIEProgErr = uvm_reg_field::type_id::create("PhyPIEProgErr",,get_full_name());
      this.PhyPIEProgErr.configure(this, 1, 12, "RO", 1, 1'h0, 1, 0, 0);
      this.PhyHWReserved = uvm_reg_field::type_id::create("PhyHWReserved",,get_full_name());
      this.PhyHWReserved.configure(this, 3, 13, "RO", 1, 3'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptStatus)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptStatus


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRunCtrl extends uvm_reg;
	rand uvm_reg_field ACSMRun;
	rand uvm_reg_field AcsmProgPtr;
	rand uvm_reg_field ACSMXlatEn;
	rand uvm_reg_field ACSMNopFlag;
	rand uvm_reg_field ACSMRptCntOverrideEn;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMRun: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   AcsmProgPtr: coverpoint {m_data[5:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	   ACSMXlatEn: coverpoint {m_data[6:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMNopFlag: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMRptCntOverrideEn: coverpoint {m_data[8:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMRunCtrl");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMRun = uvm_reg_field::type_id::create("ACSMRun",,get_full_name());
      this.ACSMRun.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.AcsmProgPtr = uvm_reg_field::type_id::create("AcsmProgPtr",,get_full_name());
      this.AcsmProgPtr.configure(this, 5, 1, "RW", 0, 5'h0, 1, 0, 0);
      this.ACSMXlatEn = uvm_reg_field::type_id::create("ACSMXlatEn",,get_full_name());
      this.ACSMXlatEn.configure(this, 1, 6, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMNopFlag = uvm_reg_field::type_id::create("ACSMNopFlag",,get_full_name());
      this.ACSMNopFlag.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMRptCntOverrideEn = uvm_reg_field::type_id::create("ACSMRptCntOverrideEn",,get_full_name());
      this.ACSMRptCntOverrideEn.configure(this, 1, 8, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRunCtrl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRunCtrl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDone extends uvm_reg;
	uvm_reg_field ACSMDone;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMDone: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMDone");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMDone = uvm_reg_field::type_id::create("ACSMDone",,get_full_name());
      this.ACSMDone.configure(this, 1, 0, "RO", 1, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDone)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDone


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStartAddr_p0 extends uvm_reg;
	rand uvm_reg_field ACSMStartAddr_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMStartAddr_p0: coverpoint {m_data[10:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {12'b??????????00};
	      wildcard bins bit_0_wr_as_1 = {12'b??????????10};
	      wildcard bins bit_0_rd_as_0 = {12'b??????????01};
	      wildcard bins bit_0_rd_as_1 = {12'b??????????11};
	      wildcard bins bit_1_wr_as_0 = {12'b?????????0?0};
	      wildcard bins bit_1_wr_as_1 = {12'b?????????1?0};
	      wildcard bins bit_1_rd_as_0 = {12'b?????????0?1};
	      wildcard bins bit_1_rd_as_1 = {12'b?????????1?1};
	      wildcard bins bit_2_wr_as_0 = {12'b????????0??0};
	      wildcard bins bit_2_wr_as_1 = {12'b????????1??0};
	      wildcard bins bit_2_rd_as_0 = {12'b????????0??1};
	      wildcard bins bit_2_rd_as_1 = {12'b????????1??1};
	      wildcard bins bit_3_wr_as_0 = {12'b???????0???0};
	      wildcard bins bit_3_wr_as_1 = {12'b???????1???0};
	      wildcard bins bit_3_rd_as_0 = {12'b???????0???1};
	      wildcard bins bit_3_rd_as_1 = {12'b???????1???1};
	      wildcard bins bit_4_wr_as_0 = {12'b??????0????0};
	      wildcard bins bit_4_wr_as_1 = {12'b??????1????0};
	      wildcard bins bit_4_rd_as_0 = {12'b??????0????1};
	      wildcard bins bit_4_rd_as_1 = {12'b??????1????1};
	      wildcard bins bit_5_wr_as_0 = {12'b?????0?????0};
	      wildcard bins bit_5_wr_as_1 = {12'b?????1?????0};
	      wildcard bins bit_5_rd_as_0 = {12'b?????0?????1};
	      wildcard bins bit_5_rd_as_1 = {12'b?????1?????1};
	      wildcard bins bit_6_wr_as_0 = {12'b????0??????0};
	      wildcard bins bit_6_wr_as_1 = {12'b????1??????0};
	      wildcard bins bit_6_rd_as_0 = {12'b????0??????1};
	      wildcard bins bit_6_rd_as_1 = {12'b????1??????1};
	      wildcard bins bit_7_wr_as_0 = {12'b???0???????0};
	      wildcard bins bit_7_wr_as_1 = {12'b???1???????0};
	      wildcard bins bit_7_rd_as_0 = {12'b???0???????1};
	      wildcard bins bit_7_rd_as_1 = {12'b???1???????1};
	      wildcard bins bit_8_wr_as_0 = {12'b??0????????0};
	      wildcard bins bit_8_wr_as_1 = {12'b??1????????0};
	      wildcard bins bit_8_rd_as_0 = {12'b??0????????1};
	      wildcard bins bit_8_rd_as_1 = {12'b??1????????1};
	      wildcard bins bit_9_wr_as_0 = {12'b?0?????????0};
	      wildcard bins bit_9_wr_as_1 = {12'b?1?????????0};
	      wildcard bins bit_9_rd_as_0 = {12'b?0?????????1};
	      wildcard bins bit_9_rd_as_1 = {12'b?1?????????1};
	      wildcard bins bit_10_wr_as_0 = {12'b0??????????0};
	      wildcard bins bit_10_wr_as_1 = {12'b1??????????0};
	      wildcard bins bit_10_rd_as_0 = {12'b0??????????1};
	      wildcard bins bit_10_rd_as_1 = {12'b1??????????1};
	      option.weight = 44;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMStartAddr_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMStartAddr_p0 = uvm_reg_field::type_id::create("ACSMStartAddr_p0",,get_full_name());
      this.ACSMStartAddr_p0.configure(this, 11, 0, "RW", 0, 11'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStartAddr_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStartAddr_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStopAddr_p0 extends uvm_reg;
	rand uvm_reg_field ACSMStopAddr_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMStopAddr_p0: coverpoint {m_data[10:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {12'b??????????00};
	      wildcard bins bit_0_wr_as_1 = {12'b??????????10};
	      wildcard bins bit_0_rd_as_0 = {12'b??????????01};
	      wildcard bins bit_0_rd_as_1 = {12'b??????????11};
	      wildcard bins bit_1_wr_as_0 = {12'b?????????0?0};
	      wildcard bins bit_1_wr_as_1 = {12'b?????????1?0};
	      wildcard bins bit_1_rd_as_0 = {12'b?????????0?1};
	      wildcard bins bit_1_rd_as_1 = {12'b?????????1?1};
	      wildcard bins bit_2_wr_as_0 = {12'b????????0??0};
	      wildcard bins bit_2_wr_as_1 = {12'b????????1??0};
	      wildcard bins bit_2_rd_as_0 = {12'b????????0??1};
	      wildcard bins bit_2_rd_as_1 = {12'b????????1??1};
	      wildcard bins bit_3_wr_as_0 = {12'b???????0???0};
	      wildcard bins bit_3_wr_as_1 = {12'b???????1???0};
	      wildcard bins bit_3_rd_as_0 = {12'b???????0???1};
	      wildcard bins bit_3_rd_as_1 = {12'b???????1???1};
	      wildcard bins bit_4_wr_as_0 = {12'b??????0????0};
	      wildcard bins bit_4_wr_as_1 = {12'b??????1????0};
	      wildcard bins bit_4_rd_as_0 = {12'b??????0????1};
	      wildcard bins bit_4_rd_as_1 = {12'b??????1????1};
	      wildcard bins bit_5_wr_as_0 = {12'b?????0?????0};
	      wildcard bins bit_5_wr_as_1 = {12'b?????1?????0};
	      wildcard bins bit_5_rd_as_0 = {12'b?????0?????1};
	      wildcard bins bit_5_rd_as_1 = {12'b?????1?????1};
	      wildcard bins bit_6_wr_as_0 = {12'b????0??????0};
	      wildcard bins bit_6_wr_as_1 = {12'b????1??????0};
	      wildcard bins bit_6_rd_as_0 = {12'b????0??????1};
	      wildcard bins bit_6_rd_as_1 = {12'b????1??????1};
	      wildcard bins bit_7_wr_as_0 = {12'b???0???????0};
	      wildcard bins bit_7_wr_as_1 = {12'b???1???????0};
	      wildcard bins bit_7_rd_as_0 = {12'b???0???????1};
	      wildcard bins bit_7_rd_as_1 = {12'b???1???????1};
	      wildcard bins bit_8_wr_as_0 = {12'b??0????????0};
	      wildcard bins bit_8_wr_as_1 = {12'b??1????????0};
	      wildcard bins bit_8_rd_as_0 = {12'b??0????????1};
	      wildcard bins bit_8_rd_as_1 = {12'b??1????????1};
	      wildcard bins bit_9_wr_as_0 = {12'b?0?????????0};
	      wildcard bins bit_9_wr_as_1 = {12'b?1?????????0};
	      wildcard bins bit_9_rd_as_0 = {12'b?0?????????1};
	      wildcard bins bit_9_rd_as_1 = {12'b?1?????????1};
	      wildcard bins bit_10_wr_as_0 = {12'b0??????????0};
	      wildcard bins bit_10_wr_as_1 = {12'b1??????????0};
	      wildcard bins bit_10_rd_as_0 = {12'b0??????????1};
	      wildcard bins bit_10_rd_as_1 = {12'b1??????????1};
	      option.weight = 44;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMStopAddr_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMStopAddr_p0 = uvm_reg_field::type_id::create("ACSMStopAddr_p0",,get_full_name());
      this.ACSMStopAddr_p0.configure(this, 11, 0, "RW", 0, 11'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStopAddr_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStopAddr_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLastAddr extends uvm_reg;
	uvm_reg_field ACSMLastAddr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMLastAddr: coverpoint {m_data[10:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {12'b??????????00};
	      wildcard bins bit_0_wr_as_1 = {12'b??????????10};
	      wildcard bins bit_0_rd = {12'b???????????1};
	      wildcard bins bit_1_wr_as_0 = {12'b?????????0?0};
	      wildcard bins bit_1_wr_as_1 = {12'b?????????1?0};
	      wildcard bins bit_1_rd = {12'b???????????1};
	      wildcard bins bit_2_wr_as_0 = {12'b????????0??0};
	      wildcard bins bit_2_wr_as_1 = {12'b????????1??0};
	      wildcard bins bit_2_rd = {12'b???????????1};
	      wildcard bins bit_3_wr_as_0 = {12'b???????0???0};
	      wildcard bins bit_3_wr_as_1 = {12'b???????1???0};
	      wildcard bins bit_3_rd = {12'b???????????1};
	      wildcard bins bit_4_wr_as_0 = {12'b??????0????0};
	      wildcard bins bit_4_wr_as_1 = {12'b??????1????0};
	      wildcard bins bit_4_rd = {12'b???????????1};
	      wildcard bins bit_5_wr_as_0 = {12'b?????0?????0};
	      wildcard bins bit_5_wr_as_1 = {12'b?????1?????0};
	      wildcard bins bit_5_rd = {12'b???????????1};
	      wildcard bins bit_6_wr_as_0 = {12'b????0??????0};
	      wildcard bins bit_6_wr_as_1 = {12'b????1??????0};
	      wildcard bins bit_6_rd = {12'b???????????1};
	      wildcard bins bit_7_wr_as_0 = {12'b???0???????0};
	      wildcard bins bit_7_wr_as_1 = {12'b???1???????0};
	      wildcard bins bit_7_rd = {12'b???????????1};
	      wildcard bins bit_8_wr_as_0 = {12'b??0????????0};
	      wildcard bins bit_8_wr_as_1 = {12'b??1????????0};
	      wildcard bins bit_8_rd = {12'b???????????1};
	      wildcard bins bit_9_wr_as_0 = {12'b?0?????????0};
	      wildcard bins bit_9_wr_as_1 = {12'b?1?????????0};
	      wildcard bins bit_9_rd = {12'b???????????1};
	      wildcard bins bit_10_wr_as_0 = {12'b0??????????0};
	      wildcard bins bit_10_wr_as_1 = {12'b1??????????0};
	      wildcard bins bit_10_rd = {12'b???????????1};
	      option.weight = 33;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMLastAddr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMLastAddr = uvm_reg_field::type_id::create("ACSMLastAddr",,get_full_name());
      this.ACSMLastAddr.configure(this, 11, 0, "RO", 1, 11'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLastAddr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLastAddr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAlgaIncVal extends uvm_reg;
	rand uvm_reg_field ACSMAlgaIncVal;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMAlgaIncVal: coverpoint {m_data[13:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {15'b?????????????00};
	      wildcard bins bit_0_wr_as_1 = {15'b?????????????10};
	      wildcard bins bit_0_rd_as_0 = {15'b?????????????01};
	      wildcard bins bit_0_rd_as_1 = {15'b?????????????11};
	      wildcard bins bit_1_wr_as_0 = {15'b????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {15'b????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {15'b????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {15'b????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {15'b???????????0??0};
	      wildcard bins bit_2_wr_as_1 = {15'b???????????1??0};
	      wildcard bins bit_2_rd_as_0 = {15'b???????????0??1};
	      wildcard bins bit_2_rd_as_1 = {15'b???????????1??1};
	      wildcard bins bit_3_wr_as_0 = {15'b??????????0???0};
	      wildcard bins bit_3_wr_as_1 = {15'b??????????1???0};
	      wildcard bins bit_3_rd_as_0 = {15'b??????????0???1};
	      wildcard bins bit_3_rd_as_1 = {15'b??????????1???1};
	      wildcard bins bit_4_wr_as_0 = {15'b?????????0????0};
	      wildcard bins bit_4_wr_as_1 = {15'b?????????1????0};
	      wildcard bins bit_4_rd_as_0 = {15'b?????????0????1};
	      wildcard bins bit_4_rd_as_1 = {15'b?????????1????1};
	      wildcard bins bit_5_wr_as_0 = {15'b????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {15'b????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {15'b????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {15'b????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {15'b???????0??????0};
	      wildcard bins bit_6_wr_as_1 = {15'b???????1??????0};
	      wildcard bins bit_6_rd_as_0 = {15'b???????0??????1};
	      wildcard bins bit_6_rd_as_1 = {15'b???????1??????1};
	      wildcard bins bit_7_wr_as_0 = {15'b??????0???????0};
	      wildcard bins bit_7_wr_as_1 = {15'b??????1???????0};
	      wildcard bins bit_7_rd_as_0 = {15'b??????0???????1};
	      wildcard bins bit_7_rd_as_1 = {15'b??????1???????1};
	      wildcard bins bit_8_wr_as_0 = {15'b?????0????????0};
	      wildcard bins bit_8_wr_as_1 = {15'b?????1????????0};
	      wildcard bins bit_8_rd_as_0 = {15'b?????0????????1};
	      wildcard bins bit_8_rd_as_1 = {15'b?????1????????1};
	      wildcard bins bit_9_wr_as_0 = {15'b????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {15'b????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {15'b????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {15'b????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {15'b???0??????????0};
	      wildcard bins bit_10_wr_as_1 = {15'b???1??????????0};
	      wildcard bins bit_10_rd_as_0 = {15'b???0??????????1};
	      wildcard bins bit_10_rd_as_1 = {15'b???1??????????1};
	      wildcard bins bit_11_wr_as_0 = {15'b??0???????????0};
	      wildcard bins bit_11_wr_as_1 = {15'b??1???????????0};
	      wildcard bins bit_11_rd_as_0 = {15'b??0???????????1};
	      wildcard bins bit_11_rd_as_1 = {15'b??1???????????1};
	      wildcard bins bit_12_wr_as_0 = {15'b?0????????????0};
	      wildcard bins bit_12_wr_as_1 = {15'b?1????????????0};
	      wildcard bins bit_12_rd_as_0 = {15'b?0????????????1};
	      wildcard bins bit_12_rd_as_1 = {15'b?1????????????1};
	      wildcard bins bit_13_wr_as_0 = {15'b0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {15'b1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {15'b0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {15'b1?????????????1};
	      option.weight = 56;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMAlgaIncVal");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMAlgaIncVal = uvm_reg_field::type_id::create("ACSMAlgaIncVal",,get_full_name());
      this.ACSMAlgaIncVal.configure(this, 14, 0, "RW", 0, 14'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAlgaIncVal)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAlgaIncVal


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAddressMask extends uvm_reg;
	rand uvm_reg_field ACSMAddressMask;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMAddressMask: coverpoint {m_data[13:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {15'b?????????????00};
	      wildcard bins bit_0_wr_as_1 = {15'b?????????????10};
	      wildcard bins bit_0_rd_as_0 = {15'b?????????????01};
	      wildcard bins bit_0_rd_as_1 = {15'b?????????????11};
	      wildcard bins bit_1_wr_as_0 = {15'b????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {15'b????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {15'b????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {15'b????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {15'b???????????0??0};
	      wildcard bins bit_2_wr_as_1 = {15'b???????????1??0};
	      wildcard bins bit_2_rd_as_0 = {15'b???????????0??1};
	      wildcard bins bit_2_rd_as_1 = {15'b???????????1??1};
	      wildcard bins bit_3_wr_as_0 = {15'b??????????0???0};
	      wildcard bins bit_3_wr_as_1 = {15'b??????????1???0};
	      wildcard bins bit_3_rd_as_0 = {15'b??????????0???1};
	      wildcard bins bit_3_rd_as_1 = {15'b??????????1???1};
	      wildcard bins bit_4_wr_as_0 = {15'b?????????0????0};
	      wildcard bins bit_4_wr_as_1 = {15'b?????????1????0};
	      wildcard bins bit_4_rd_as_0 = {15'b?????????0????1};
	      wildcard bins bit_4_rd_as_1 = {15'b?????????1????1};
	      wildcard bins bit_5_wr_as_0 = {15'b????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {15'b????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {15'b????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {15'b????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {15'b???????0??????0};
	      wildcard bins bit_6_wr_as_1 = {15'b???????1??????0};
	      wildcard bins bit_6_rd_as_0 = {15'b???????0??????1};
	      wildcard bins bit_6_rd_as_1 = {15'b???????1??????1};
	      wildcard bins bit_7_wr_as_0 = {15'b??????0???????0};
	      wildcard bins bit_7_wr_as_1 = {15'b??????1???????0};
	      wildcard bins bit_7_rd_as_0 = {15'b??????0???????1};
	      wildcard bins bit_7_rd_as_1 = {15'b??????1???????1};
	      wildcard bins bit_8_wr_as_0 = {15'b?????0????????0};
	      wildcard bins bit_8_wr_as_1 = {15'b?????1????????0};
	      wildcard bins bit_8_rd_as_0 = {15'b?????0????????1};
	      wildcard bins bit_8_rd_as_1 = {15'b?????1????????1};
	      wildcard bins bit_9_wr_as_0 = {15'b????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {15'b????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {15'b????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {15'b????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {15'b???0??????????0};
	      wildcard bins bit_10_wr_as_1 = {15'b???1??????????0};
	      wildcard bins bit_10_rd_as_0 = {15'b???0??????????1};
	      wildcard bins bit_10_rd_as_1 = {15'b???1??????????1};
	      wildcard bins bit_11_wr_as_0 = {15'b??0???????????0};
	      wildcard bins bit_11_wr_as_1 = {15'b??1???????????0};
	      wildcard bins bit_11_rd_as_0 = {15'b??0???????????1};
	      wildcard bins bit_11_rd_as_1 = {15'b??1???????????1};
	      wildcard bins bit_12_wr_as_0 = {15'b?0????????????0};
	      wildcard bins bit_12_wr_as_1 = {15'b?1????????????0};
	      wildcard bins bit_12_rd_as_0 = {15'b?0????????????1};
	      wildcard bins bit_12_rd_as_1 = {15'b?1????????????1};
	      wildcard bins bit_13_wr_as_0 = {15'b0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {15'b1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {15'b0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {15'b1?????????????1};
	      option.weight = 56;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMAddressMask");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMAddressMask = uvm_reg_field::type_id::create("ACSMAddressMask",,get_full_name());
      this.ACSMAddressMask.configure(this, 14, 0, "RW", 0, 14'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAddressMask)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAddressMask


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMOuterLoopRepeatCnt extends uvm_reg;
	rand uvm_reg_field ACSMOuterLoopRepeatCnt;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMOuterLoopRepeatCnt: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMOuterLoopRepeatCnt");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMOuterLoopRepeatCnt = uvm_reg_field::type_id::create("ACSMOuterLoopRepeatCnt",,get_full_name());
      this.ACSMOuterLoopRepeatCnt.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMOuterLoopRepeatCnt)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMOuterLoopRepeatCnt


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeControl extends uvm_reg;
	rand uvm_reg_field ACSMCkeControl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMCkeControl: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMCkeControl");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMCkeControl = uvm_reg_field::type_id::create("ACSMCkeControl",,get_full_name());
      this.ACSMCkeControl.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeControl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeControl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeStatus extends uvm_reg;
	uvm_reg_field ACSMCkeStatus;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMCkeStatus: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMCkeStatus");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMCkeStatus = uvm_reg_field::type_id::create("ACSMCkeStatus",,get_full_name());
      this.ACSMCkeStatus.configure(this, 1, 0, "RO", 1, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeStatus)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeStatus


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnControl extends uvm_reg;
	rand uvm_reg_field ACSMWckEnControl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckEnControl: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckEnControl");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckEnControl = uvm_reg_field::type_id::create("ACSMWckEnControl",,get_full_name());
      this.ACSMWckEnControl.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnControl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnControl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnStatus extends uvm_reg;
	uvm_reg_field ACSMWckEnStatus;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckEnStatus: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckEnStatus");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckEnStatus = uvm_reg_field::type_id::create("ACSMWckEnStatus",,get_full_name());
      this.ACSMWckEnStatus.configure(this, 1, 0, "RO", 1, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnStatus)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnStatus


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxEnPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMRxEnDelay;
	rand uvm_reg_field ACSMRxEnDelayReserved;
	rand uvm_reg_field ACSMRxEnWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMRxEnDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMRxEnDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMRxEnWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMRxEnPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMRxEnDelay = uvm_reg_field::type_id::create("ACSMRxEnDelay",,get_full_name());
      this.ACSMRxEnDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMRxEnDelayReserved = uvm_reg_field::type_id::create("ACSMRxEnDelayReserved",,get_full_name());
      this.ACSMRxEnDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMRxEnWidth = uvm_reg_field::type_id::create("ACSMRxEnWidth",,get_full_name());
      this.ACSMRxEnWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxEnPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxEnPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxValPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMRxValDelay;
	rand uvm_reg_field ACSMRxValDelayReserved;
	rand uvm_reg_field ACSMRxValWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMRxValDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMRxValDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMRxValWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMRxValPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMRxValDelay = uvm_reg_field::type_id::create("ACSMRxValDelay",,get_full_name());
      this.ACSMRxValDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMRxValDelayReserved = uvm_reg_field::type_id::create("ACSMRxValDelayReserved",,get_full_name());
      this.ACSMRxValDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMRxValWidth = uvm_reg_field::type_id::create("ACSMRxValWidth",,get_full_name());
      this.ACSMRxValWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxValPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxValPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMTxEnPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMTxEnDelay;
	rand uvm_reg_field ACSMTxEnDelayReserved;
	rand uvm_reg_field ACSMTxEnWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMTxEnDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMTxEnDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMTxEnWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMTxEnPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMTxEnDelay = uvm_reg_field::type_id::create("ACSMTxEnDelay",,get_full_name());
      this.ACSMTxEnDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMTxEnDelayReserved = uvm_reg_field::type_id::create("ACSMTxEnDelayReserved",,get_full_name());
      this.ACSMTxEnDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMTxEnWidth = uvm_reg_field::type_id::create("ACSMTxEnWidth",,get_full_name());
      this.ACSMTxEnWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMTxEnPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMTxEnPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWrcsPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWrcsDelay;
	rand uvm_reg_field ACSMWrcsDelayReserved;
	rand uvm_reg_field ACSMWrcsWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWrcsDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWrcsDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWrcsWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWrcsPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWrcsDelay = uvm_reg_field::type_id::create("ACSMWrcsDelay",,get_full_name());
      this.ACSMWrcsDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWrcsDelayReserved = uvm_reg_field::type_id::create("ACSMWrcsDelayReserved",,get_full_name());
      this.ACSMWrcsDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWrcsWidth = uvm_reg_field::type_id::create("ACSMWrcsWidth",,get_full_name());
      this.ACSMWrcsWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWrcsPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWrcsPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRdcsPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMRdcsDelay;
	rand uvm_reg_field ACSMRdcsDelayReserved;
	rand uvm_reg_field ACSMRdcsWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMRdcsDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMRdcsDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMRdcsWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMRdcsPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMRdcsDelay = uvm_reg_field::type_id::create("ACSMRdcsDelay",,get_full_name());
      this.ACSMRdcsDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMRdcsDelayReserved = uvm_reg_field::type_id::create("ACSMRdcsDelayReserved",,get_full_name());
      this.ACSMRdcsDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMRdcsWidth = uvm_reg_field::type_id::create("ACSMRdcsWidth",,get_full_name());
      this.ACSMRdcsWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRdcsPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRdcsPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMInfiniteOLRC extends uvm_reg;
	rand uvm_reg_field ACSMInfiniteOLRC;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMInfiniteOLRC: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMInfiniteOLRC");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMInfiniteOLRC = uvm_reg_field::type_id::create("ACSMInfiniteOLRC",,get_full_name());
      this.ACSMInfiniteOLRC.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMInfiniteOLRC)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMInfiniteOLRC


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultAddr extends uvm_reg;
	rand uvm_reg_field ACSMDefaultAddr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMDefaultAddr: coverpoint {m_data[13:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {15'b?????????????00};
	      wildcard bins bit_0_wr_as_1 = {15'b?????????????10};
	      wildcard bins bit_0_rd_as_0 = {15'b?????????????01};
	      wildcard bins bit_0_rd_as_1 = {15'b?????????????11};
	      wildcard bins bit_1_wr_as_0 = {15'b????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {15'b????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {15'b????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {15'b????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {15'b???????????0??0};
	      wildcard bins bit_2_wr_as_1 = {15'b???????????1??0};
	      wildcard bins bit_2_rd_as_0 = {15'b???????????0??1};
	      wildcard bins bit_2_rd_as_1 = {15'b???????????1??1};
	      wildcard bins bit_3_wr_as_0 = {15'b??????????0???0};
	      wildcard bins bit_3_wr_as_1 = {15'b??????????1???0};
	      wildcard bins bit_3_rd_as_0 = {15'b??????????0???1};
	      wildcard bins bit_3_rd_as_1 = {15'b??????????1???1};
	      wildcard bins bit_4_wr_as_0 = {15'b?????????0????0};
	      wildcard bins bit_4_wr_as_1 = {15'b?????????1????0};
	      wildcard bins bit_4_rd_as_0 = {15'b?????????0????1};
	      wildcard bins bit_4_rd_as_1 = {15'b?????????1????1};
	      wildcard bins bit_5_wr_as_0 = {15'b????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {15'b????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {15'b????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {15'b????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {15'b???????0??????0};
	      wildcard bins bit_6_wr_as_1 = {15'b???????1??????0};
	      wildcard bins bit_6_rd_as_0 = {15'b???????0??????1};
	      wildcard bins bit_6_rd_as_1 = {15'b???????1??????1};
	      wildcard bins bit_7_wr_as_0 = {15'b??????0???????0};
	      wildcard bins bit_7_wr_as_1 = {15'b??????1???????0};
	      wildcard bins bit_7_rd_as_0 = {15'b??????0???????1};
	      wildcard bins bit_7_rd_as_1 = {15'b??????1???????1};
	      wildcard bins bit_8_wr_as_0 = {15'b?????0????????0};
	      wildcard bins bit_8_wr_as_1 = {15'b?????1????????0};
	      wildcard bins bit_8_rd_as_0 = {15'b?????0????????1};
	      wildcard bins bit_8_rd_as_1 = {15'b?????1????????1};
	      wildcard bins bit_9_wr_as_0 = {15'b????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {15'b????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {15'b????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {15'b????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {15'b???0??????????0};
	      wildcard bins bit_10_wr_as_1 = {15'b???1??????????0};
	      wildcard bins bit_10_rd_as_0 = {15'b???0??????????1};
	      wildcard bins bit_10_rd_as_1 = {15'b???1??????????1};
	      wildcard bins bit_11_wr_as_0 = {15'b??0???????????0};
	      wildcard bins bit_11_wr_as_1 = {15'b??1???????????0};
	      wildcard bins bit_11_rd_as_0 = {15'b??0???????????1};
	      wildcard bins bit_11_rd_as_1 = {15'b??1???????????1};
	      wildcard bins bit_12_wr_as_0 = {15'b?0????????????0};
	      wildcard bins bit_12_wr_as_1 = {15'b?1????????????0};
	      wildcard bins bit_12_rd_as_0 = {15'b?0????????????1};
	      wildcard bins bit_12_rd_as_1 = {15'b?1????????????1};
	      wildcard bins bit_13_wr_as_0 = {15'b0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {15'b1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {15'b0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {15'b1?????????????1};
	      option.weight = 56;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMDefaultAddr");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMDefaultAddr = uvm_reg_field::type_id::create("ACSMDefaultAddr",,get_full_name());
      this.ACSMDefaultAddr.configure(this, 14, 0, "RW", 0, 14'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultAddr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultAddr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultCs extends uvm_reg;
	rand uvm_reg_field ACSMDefaultCs;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMDefaultCs: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMDefaultCs");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMDefaultCs = uvm_reg_field::type_id::create("ACSMDefaultCs",,get_full_name());
      this.ACSMDefaultCs.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultCs)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultCs


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStaticCtrl extends uvm_reg;
	rand uvm_reg_field ACSMPhaseControl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMPhaseControl: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMStaticCtrl");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMPhaseControl = uvm_reg_field::type_id::create("ACSMPhaseControl",,get_full_name());
      this.ACSMPhaseControl.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStaticCtrl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStaticCtrl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticLoPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckWriteStaticLoDelay;
	rand uvm_reg_field ACSMWckWriteStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckWriteStaticLoWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckWriteStaticLoDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckWriteStaticLoDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckWriteStaticLoWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticLoPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckWriteStaticLoDelay = uvm_reg_field::type_id::create("ACSMWckWriteStaticLoDelay",,get_full_name());
      this.ACSMWckWriteStaticLoDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckWriteStaticLoDelayReserved = uvm_reg_field::type_id::create("ACSMWckWriteStaticLoDelayReserved",,get_full_name());
      this.ACSMWckWriteStaticLoDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckWriteStaticLoWidth = uvm_reg_field::type_id::create("ACSMWckWriteStaticLoWidth",,get_full_name());
      this.ACSMWckWriteStaticLoWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticLoPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticLoPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticHiPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckWriteStaticHiDelay;
	rand uvm_reg_field ACSMWckWriteStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckWriteStaticHiWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckWriteStaticHiDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckWriteStaticHiDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckWriteStaticHiWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticHiPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckWriteStaticHiDelay = uvm_reg_field::type_id::create("ACSMWckWriteStaticHiDelay",,get_full_name());
      this.ACSMWckWriteStaticHiDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckWriteStaticHiDelayReserved = uvm_reg_field::type_id::create("ACSMWckWriteStaticHiDelayReserved",,get_full_name());
      this.ACSMWckWriteStaticHiDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckWriteStaticHiWidth = uvm_reg_field::type_id::create("ACSMWckWriteStaticHiWidth",,get_full_name());
      this.ACSMWckWriteStaticHiWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticHiPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticHiPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteTogglePulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckWriteToggleDelay;
	rand uvm_reg_field ACSMWckWriteToggleDelayReserved;
	rand uvm_reg_field ACSMWckWriteToggleWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckWriteToggleDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckWriteToggleDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckWriteToggleWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteTogglePulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckWriteToggleDelay = uvm_reg_field::type_id::create("ACSMWckWriteToggleDelay",,get_full_name());
      this.ACSMWckWriteToggleDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckWriteToggleDelayReserved = uvm_reg_field::type_id::create("ACSMWckWriteToggleDelayReserved",,get_full_name());
      this.ACSMWckWriteToggleDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckWriteToggleWidth = uvm_reg_field::type_id::create("ACSMWckWriteToggleWidth",,get_full_name());
      this.ACSMWckWriteToggleWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteTogglePulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteTogglePulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteFastTogglePulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckWriteFastToggleDelay;
	rand uvm_reg_field ACSMWckWriteFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckWriteFastToggleWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckWriteFastToggleDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckWriteFastToggleDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckWriteFastToggleWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteFastTogglePulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckWriteFastToggleDelay = uvm_reg_field::type_id::create("ACSMWckWriteFastToggleDelay",,get_full_name());
      this.ACSMWckWriteFastToggleDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckWriteFastToggleDelayReserved = uvm_reg_field::type_id::create("ACSMWckWriteFastToggleDelayReserved",,get_full_name());
      this.ACSMWckWriteFastToggleDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckWriteFastToggleWidth = uvm_reg_field::type_id::create("ACSMWckWriteFastToggleWidth",,get_full_name());
      this.ACSMWckWriteFastToggleWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteFastTogglePulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteFastTogglePulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticLoPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckReadStaticLoDelay;
	rand uvm_reg_field ACSMWckReadStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckReadStaticLoWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckReadStaticLoDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckReadStaticLoDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckReadStaticLoWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticLoPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckReadStaticLoDelay = uvm_reg_field::type_id::create("ACSMWckReadStaticLoDelay",,get_full_name());
      this.ACSMWckReadStaticLoDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckReadStaticLoDelayReserved = uvm_reg_field::type_id::create("ACSMWckReadStaticLoDelayReserved",,get_full_name());
      this.ACSMWckReadStaticLoDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckReadStaticLoWidth = uvm_reg_field::type_id::create("ACSMWckReadStaticLoWidth",,get_full_name());
      this.ACSMWckReadStaticLoWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticLoPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticLoPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticHiPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckReadStaticHiDelay;
	rand uvm_reg_field ACSMWckReadStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckReadStaticHiWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckReadStaticHiDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckReadStaticHiDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckReadStaticHiWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticHiPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckReadStaticHiDelay = uvm_reg_field::type_id::create("ACSMWckReadStaticHiDelay",,get_full_name());
      this.ACSMWckReadStaticHiDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckReadStaticHiDelayReserved = uvm_reg_field::type_id::create("ACSMWckReadStaticHiDelayReserved",,get_full_name());
      this.ACSMWckReadStaticHiDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckReadStaticHiWidth = uvm_reg_field::type_id::create("ACSMWckReadStaticHiWidth",,get_full_name());
      this.ACSMWckReadStaticHiWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticHiPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticHiPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadTogglePulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckReadToggleDelay;
	rand uvm_reg_field ACSMWckReadToggleDelayReserved;
	rand uvm_reg_field ACSMWckReadToggleWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckReadToggleDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckReadToggleDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckReadToggleWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckReadTogglePulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckReadToggleDelay = uvm_reg_field::type_id::create("ACSMWckReadToggleDelay",,get_full_name());
      this.ACSMWckReadToggleDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckReadToggleDelayReserved = uvm_reg_field::type_id::create("ACSMWckReadToggleDelayReserved",,get_full_name());
      this.ACSMWckReadToggleDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckReadToggleWidth = uvm_reg_field::type_id::create("ACSMWckReadToggleWidth",,get_full_name());
      this.ACSMWckReadToggleWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadTogglePulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadTogglePulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadFastTogglePulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckReadFastToggleDelay;
	rand uvm_reg_field ACSMWckReadFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckReadFastToggleWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckReadFastToggleDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckReadFastToggleDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckReadFastToggleWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckReadFastTogglePulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckReadFastToggleDelay = uvm_reg_field::type_id::create("ACSMWckReadFastToggleDelay",,get_full_name());
      this.ACSMWckReadFastToggleDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckReadFastToggleDelayReserved = uvm_reg_field::type_id::create("ACSMWckReadFastToggleDelayReserved",,get_full_name());
      this.ACSMWckReadFastToggleDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckReadFastToggleWidth = uvm_reg_field::type_id::create("ACSMWckReadFastToggleWidth",,get_full_name());
      this.ACSMWckReadFastToggleWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadFastTogglePulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadFastTogglePulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticLoPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckFreqSwStaticLoDelay;
	rand uvm_reg_field ACSMWckFreqSwStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwStaticLoWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckFreqSwStaticLoDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckFreqSwStaticLoDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckFreqSwStaticLoWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticLoPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckFreqSwStaticLoDelay = uvm_reg_field::type_id::create("ACSMWckFreqSwStaticLoDelay",,get_full_name());
      this.ACSMWckFreqSwStaticLoDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckFreqSwStaticLoDelayReserved = uvm_reg_field::type_id::create("ACSMWckFreqSwStaticLoDelayReserved",,get_full_name());
      this.ACSMWckFreqSwStaticLoDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckFreqSwStaticLoWidth = uvm_reg_field::type_id::create("ACSMWckFreqSwStaticLoWidth",,get_full_name());
      this.ACSMWckFreqSwStaticLoWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticLoPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticLoPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticHiPulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckFreqSwStaticHiDelay;
	rand uvm_reg_field ACSMWckFreqSwStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwStaticHiWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckFreqSwStaticHiDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckFreqSwStaticHiDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckFreqSwStaticHiWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticHiPulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckFreqSwStaticHiDelay = uvm_reg_field::type_id::create("ACSMWckFreqSwStaticHiDelay",,get_full_name());
      this.ACSMWckFreqSwStaticHiDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckFreqSwStaticHiDelayReserved = uvm_reg_field::type_id::create("ACSMWckFreqSwStaticHiDelayReserved",,get_full_name());
      this.ACSMWckFreqSwStaticHiDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckFreqSwStaticHiWidth = uvm_reg_field::type_id::create("ACSMWckFreqSwStaticHiWidth",,get_full_name());
      this.ACSMWckFreqSwStaticHiWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticHiPulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticHiPulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwTogglePulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckFreqSwToggleDelay;
	rand uvm_reg_field ACSMWckFreqSwToggleDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwToggleWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckFreqSwToggleDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckFreqSwToggleDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckFreqSwToggleWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwTogglePulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckFreqSwToggleDelay = uvm_reg_field::type_id::create("ACSMWckFreqSwToggleDelay",,get_full_name());
      this.ACSMWckFreqSwToggleDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckFreqSwToggleDelayReserved = uvm_reg_field::type_id::create("ACSMWckFreqSwToggleDelayReserved",,get_full_name());
      this.ACSMWckFreqSwToggleDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckFreqSwToggleWidth = uvm_reg_field::type_id::create("ACSMWckFreqSwToggleWidth",,get_full_name());
      this.ACSMWckFreqSwToggleWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwTogglePulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwTogglePulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwFastTogglePulse_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckFreqSwFastToggleDelay;
	rand uvm_reg_field ACSMWckFreqSwFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwFastToggleWidth;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckFreqSwFastToggleDelay: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   ACSMWckFreqSwFastToggleDelayReserved: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   ACSMWckFreqSwFastToggleWidth: coverpoint {m_data[13:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwFastTogglePulse_p0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckFreqSwFastToggleDelay = uvm_reg_field::type_id::create("ACSMWckFreqSwFastToggleDelay",,get_full_name());
      this.ACSMWckFreqSwFastToggleDelay.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 0);
      this.ACSMWckFreqSwFastToggleDelayReserved = uvm_reg_field::type_id::create("ACSMWckFreqSwFastToggleDelayReserved",,get_full_name());
      this.ACSMWckFreqSwFastToggleDelayReserved.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.ACSMWckFreqSwFastToggleWidth = uvm_reg_field::type_id::create("ACSMWckFreqSwFastToggleWidth",,get_full_name());
      this.ACSMWckFreqSwFastToggleWidth.configure(this, 6, 8, "RW", 0, 6'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwFastTogglePulse_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwFastTogglePulse_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreeRunMode_p0 extends uvm_reg;
	rand uvm_reg_field ACSMWckFreeRunMode_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMWckFreeRunMode_p0: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMWckFreeRunMode_p0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMWckFreeRunMode_p0 = uvm_reg_field::type_id::create("ACSMWckFreeRunMode_p0",,get_full_name());
      this.ACSMWckFreeRunMode_p0.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreeRunMode_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreeRunMode_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockEnable extends uvm_reg;
	rand uvm_reg_field ACSMLowSpeedClockEnable;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMLowSpeedClockEnable: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockEnable");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMLowSpeedClockEnable = uvm_reg_field::type_id::create("ACSMLowSpeedClockEnable",,get_full_name());
      this.ACSMLowSpeedClockEnable.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockEnable)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockEnable


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockDelay extends uvm_reg;
	rand uvm_reg_field ACSMLowSpeedClockDelay;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMLowSpeedClockDelay: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockDelay");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMLowSpeedClockDelay = uvm_reg_field::type_id::create("ACSMLowSpeedClockDelay",,get_full_name());
      this.ACSMLowSpeedClockDelay.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockDelay)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockDelay


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntOverride_p0 extends uvm_reg;
	rand uvm_reg_field ACSMRptCntOverride_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMRptCntOverride_p0: coverpoint {m_data[7:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd_as_0 = {9'b???????01};
	      wildcard bins bit_0_rd_as_1 = {9'b???????11};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd_as_0 = {9'b??????0?1};
	      wildcard bins bit_1_rd_as_1 = {9'b??????1?1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd_as_0 = {9'b?????0??1};
	      wildcard bins bit_2_rd_as_1 = {9'b?????1??1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd_as_0 = {9'b????0???1};
	      wildcard bins bit_3_rd_as_1 = {9'b????1???1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd_as_0 = {9'b???0????1};
	      wildcard bins bit_4_rd_as_1 = {9'b???1????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd_as_0 = {9'b??0?????1};
	      wildcard bins bit_5_rd_as_1 = {9'b??1?????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd_as_0 = {9'b?0??????1};
	      wildcard bins bit_6_rd_as_1 = {9'b?1??????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd_as_0 = {9'b0???????1};
	      wildcard bins bit_7_rd_as_1 = {9'b1???????1};
	      option.weight = 32;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMRptCntOverride_p0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMRptCntOverride_p0 = uvm_reg_field::type_id::create("ACSMRptCntOverride_p0",,get_full_name());
      this.ACSMRptCntOverride_p0.configure(this, 8, 0, "RW", 0, 8'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntOverride_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntOverride_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntDbl_p0 extends uvm_reg;
	rand uvm_reg_field ACSMRptCntDbl_p0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMRptCntDbl_p0: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMRptCntDbl_p0");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMRptCntDbl_p0 = uvm_reg_field::type_id::create("ACSMRptCntDbl_p0",,get_full_name());
      this.ACSMRptCntDbl_p0.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntDbl_p0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntDbl_p0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityStatus extends uvm_reg;
	uvm_reg_field ACSMParityStatus;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMParityStatus: coverpoint {m_data[7:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd = {9'b????????1};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd = {9'b????????1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd = {9'b????????1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd = {9'b????????1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd = {9'b????????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd = {9'b????????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd = {9'b????????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd = {9'b????????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMParityStatus");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMParityStatus = uvm_reg_field::type_id::create("ACSMParityStatus",,get_full_name());
      this.ACSMParityStatus.configure(this, 8, 0, "RO", 1, 8'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityStatus)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityStatus


class ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnBypass extends uvm_reg;
	rand uvm_reg_field HwtLpCsEnBypass;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   HwtLpCsEnBypass: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnBypass");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.HwtLpCsEnBypass = uvm_reg_field::type_id::create("HwtLpCsEnBypass",,get_full_name());
      this.HwtLpCsEnBypass.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnBypass)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnBypass


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMNopAddr extends uvm_reg;
	rand uvm_reg_field ACSMNopAddr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMNopAddr: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMNopAddr");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMNopAddr = uvm_reg_field::type_id::create("ACSMNopAddr",,get_full_name());
      this.ACSMNopAddr.configure(this, 7, 0, "RW", 0, 7'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMNopAddr)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMNopAddr


class ral_reg_DWC_DDRPHYA_PPGC0_p0_SnoopCntrl extends uvm_reg;
	rand uvm_reg_field SnoopCntrl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   SnoopCntrl: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_SnoopCntrl");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.SnoopCntrl = uvm_reg_field::type_id::create("SnoopCntrl",,get_full_name());
      this.SnoopCntrl.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_SnoopCntrl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_SnoopCntrl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityInvert extends uvm_reg;
	rand uvm_reg_field ACSMParityInvert;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   ACSMParityInvert: coverpoint {m_data[7:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd_as_0 = {9'b???????01};
	      wildcard bins bit_0_rd_as_1 = {9'b???????11};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd_as_0 = {9'b??????0?1};
	      wildcard bins bit_1_rd_as_1 = {9'b??????1?1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd_as_0 = {9'b?????0??1};
	      wildcard bins bit_2_rd_as_1 = {9'b?????1??1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd_as_0 = {9'b????0???1};
	      wildcard bins bit_3_rd_as_1 = {9'b????1???1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd_as_0 = {9'b???0????1};
	      wildcard bins bit_4_rd_as_1 = {9'b???1????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd_as_0 = {9'b??0?????1};
	      wildcard bins bit_5_rd_as_1 = {9'b??1?????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd_as_0 = {9'b?0??????1};
	      wildcard bins bit_6_rd_as_1 = {9'b?1??????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd_as_0 = {9'b0???????1};
	      wildcard bins bit_7_rd_as_1 = {9'b1???????1};
	      option.weight = 32;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_ACSMParityInvert");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.ACSMParityInvert = uvm_reg_field::type_id::create("ACSMParityInvert",,get_full_name());
      this.ACSMParityInvert.configure(this, 8, 0, "RW", 0, 8'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityInvert)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityInvert


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmPsIndx extends uvm_reg;
	rand uvm_reg_field AcsmPsIndx;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmPsIndx: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmPsIndx");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmPsIndx = uvm_reg_field::type_id::create("AcsmPsIndx",,get_full_name());
      this.AcsmPsIndx.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmPsIndx)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmPsIndx


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmDynPtrCtrl extends uvm_reg;
	rand uvm_reg_field AcsmDynPtrCtrl;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmDynPtrCtrl: coverpoint {m_data[2:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmDynPtrCtrl");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmDynPtrCtrl = uvm_reg_field::type_id::create("AcsmDynPtrCtrl",,get_full_name());
      this.AcsmDynPtrCtrl.configure(this, 3, 0, "RW", 0, 3'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmDynPtrCtrl)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmDynPtrCtrl


class ral_reg_DWC_DDRPHYA_PPGC0_p0_FspState extends uvm_reg;
	rand uvm_reg_field DramFsp0xPhyPs;
	rand uvm_reg_field DramFsp1xPhyPs;
	rand uvm_reg_field DramFsp2xPhyPs;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DramFsp0xPhyPs: coverpoint {m_data[4:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	   DramFsp1xPhyPs: coverpoint {m_data[9:5], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	   DramFsp2xPhyPs: coverpoint {m_data[14:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {6'b????00};
	      wildcard bins bit_0_wr_as_1 = {6'b????10};
	      wildcard bins bit_0_rd_as_0 = {6'b????01};
	      wildcard bins bit_0_rd_as_1 = {6'b????11};
	      wildcard bins bit_1_wr_as_0 = {6'b???0?0};
	      wildcard bins bit_1_wr_as_1 = {6'b???1?0};
	      wildcard bins bit_1_rd_as_0 = {6'b???0?1};
	      wildcard bins bit_1_rd_as_1 = {6'b???1?1};
	      wildcard bins bit_2_wr_as_0 = {6'b??0??0};
	      wildcard bins bit_2_wr_as_1 = {6'b??1??0};
	      wildcard bins bit_2_rd_as_0 = {6'b??0??1};
	      wildcard bins bit_2_rd_as_1 = {6'b??1??1};
	      wildcard bins bit_3_wr_as_0 = {6'b?0???0};
	      wildcard bins bit_3_wr_as_1 = {6'b?1???0};
	      wildcard bins bit_3_rd_as_0 = {6'b?0???1};
	      wildcard bins bit_3_rd_as_1 = {6'b?1???1};
	      wildcard bins bit_4_wr_as_0 = {6'b0????0};
	      wildcard bins bit_4_wr_as_1 = {6'b1????0};
	      wildcard bins bit_4_rd_as_0 = {6'b0????1};
	      wildcard bins bit_4_rd_as_1 = {6'b1????1};
	      option.weight = 20;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_FspState");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DramFsp0xPhyPs = uvm_reg_field::type_id::create("DramFsp0xPhyPs",,get_full_name());
      this.DramFsp0xPhyPs.configure(this, 5, 0, "RW", 0, 5'h0, 1, 0, 0);
      this.DramFsp1xPhyPs = uvm_reg_field::type_id::create("DramFsp1xPhyPs",,get_full_name());
      this.DramFsp1xPhyPs.configure(this, 5, 5, "RW", 0, 5'h0, 1, 0, 0);
      this.DramFsp2xPhyPs = uvm_reg_field::type_id::create("DramFsp2xPhyPs",,get_full_name());
      this.DramFsp2xPhyPs.configure(this, 5, 10, "RW", 0, 5'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_FspState)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_FspState


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable0 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal0;
	rand uvm_reg_field AcsmMapTableVal1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal0: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal1: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal0 = uvm_reg_field::type_id::create("AcsmMapTableVal0",,get_full_name());
      this.AcsmMapTableVal0.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal1 = uvm_reg_field::type_id::create("AcsmMapTableVal1",,get_full_name());
      this.AcsmMapTableVal1.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable1 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal2;
	rand uvm_reg_field AcsmMapTableVal3;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal2: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal3: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal2 = uvm_reg_field::type_id::create("AcsmMapTableVal2",,get_full_name());
      this.AcsmMapTableVal2.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal3 = uvm_reg_field::type_id::create("AcsmMapTableVal3",,get_full_name());
      this.AcsmMapTableVal3.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable2 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal4;
	rand uvm_reg_field AcsmMapTableVal5;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal4: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal5: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable2");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal4 = uvm_reg_field::type_id::create("AcsmMapTableVal4",,get_full_name());
      this.AcsmMapTableVal4.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal5 = uvm_reg_field::type_id::create("AcsmMapTableVal5",,get_full_name());
      this.AcsmMapTableVal5.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable2)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable2


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable3 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal6;
	rand uvm_reg_field AcsmMapTableVal7;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal6: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal7: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable3");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal6 = uvm_reg_field::type_id::create("AcsmMapTableVal6",,get_full_name());
      this.AcsmMapTableVal6.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal7 = uvm_reg_field::type_id::create("AcsmMapTableVal7",,get_full_name());
      this.AcsmMapTableVal7.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable3)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable3


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable4 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal8;
	rand uvm_reg_field AcsmMapTableVal9;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal8: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal9: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable4");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal8 = uvm_reg_field::type_id::create("AcsmMapTableVal8",,get_full_name());
      this.AcsmMapTableVal8.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal9 = uvm_reg_field::type_id::create("AcsmMapTableVal9",,get_full_name());
      this.AcsmMapTableVal9.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable4)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable4


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable5 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal10;
	rand uvm_reg_field AcsmMapTableVal11;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal10: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal11: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable5");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal10 = uvm_reg_field::type_id::create("AcsmMapTableVal10",,get_full_name());
      this.AcsmMapTableVal10.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal11 = uvm_reg_field::type_id::create("AcsmMapTableVal11",,get_full_name());
      this.AcsmMapTableVal11.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable5)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable5


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable6 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal12;
	rand uvm_reg_field AcsmMapTableVal13;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal12: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal13: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable6");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal12 = uvm_reg_field::type_id::create("AcsmMapTableVal12",,get_full_name());
      this.AcsmMapTableVal12.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal13 = uvm_reg_field::type_id::create("AcsmMapTableVal13",,get_full_name());
      this.AcsmMapTableVal13.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable6)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable6


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable7 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal14;
	rand uvm_reg_field AcsmMapTableVal15;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal14: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal15: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable7");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal14 = uvm_reg_field::type_id::create("AcsmMapTableVal14",,get_full_name());
      this.AcsmMapTableVal14.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal15 = uvm_reg_field::type_id::create("AcsmMapTableVal15",,get_full_name());
      this.AcsmMapTableVal15.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable7)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable7


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable8 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal16;
	rand uvm_reg_field AcsmMapTableVal17;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal16: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal17: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable8");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal16 = uvm_reg_field::type_id::create("AcsmMapTableVal16",,get_full_name());
      this.AcsmMapTableVal16.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal17 = uvm_reg_field::type_id::create("AcsmMapTableVal17",,get_full_name());
      this.AcsmMapTableVal17.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable8)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable8


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable9 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal18;
	rand uvm_reg_field AcsmMapTableVal19;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal18: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal19: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable9");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal18 = uvm_reg_field::type_id::create("AcsmMapTableVal18",,get_full_name());
      this.AcsmMapTableVal18.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal19 = uvm_reg_field::type_id::create("AcsmMapTableVal19",,get_full_name());
      this.AcsmMapTableVal19.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable9)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable9


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable10 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal20;
	rand uvm_reg_field AcsmMapTableVal21;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal20: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal21: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable10");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal20 = uvm_reg_field::type_id::create("AcsmMapTableVal20",,get_full_name());
      this.AcsmMapTableVal20.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal21 = uvm_reg_field::type_id::create("AcsmMapTableVal21",,get_full_name());
      this.AcsmMapTableVal21.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable10)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable10


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable11 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal22;
	rand uvm_reg_field AcsmMapTableVal23;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal22: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal23: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable11");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal22 = uvm_reg_field::type_id::create("AcsmMapTableVal22",,get_full_name());
      this.AcsmMapTableVal22.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal23 = uvm_reg_field::type_id::create("AcsmMapTableVal23",,get_full_name());
      this.AcsmMapTableVal23.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable11)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable11


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable12 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal24;
	rand uvm_reg_field AcsmMapTableVal25;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal24: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal25: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable12");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal24 = uvm_reg_field::type_id::create("AcsmMapTableVal24",,get_full_name());
      this.AcsmMapTableVal24.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal25 = uvm_reg_field::type_id::create("AcsmMapTableVal25",,get_full_name());
      this.AcsmMapTableVal25.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable12)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable12


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable13 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal26;
	rand uvm_reg_field AcsmMapTableVal27;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal26: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal27: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable13");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal26 = uvm_reg_field::type_id::create("AcsmMapTableVal26",,get_full_name());
      this.AcsmMapTableVal26.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal27 = uvm_reg_field::type_id::create("AcsmMapTableVal27",,get_full_name());
      this.AcsmMapTableVal27.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable13)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable13


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable14 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal28;
	rand uvm_reg_field AcsmMapTableVal29;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal28: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal29: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable14");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal28 = uvm_reg_field::type_id::create("AcsmMapTableVal28",,get_full_name());
      this.AcsmMapTableVal28.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal29 = uvm_reg_field::type_id::create("AcsmMapTableVal29",,get_full_name());
      this.AcsmMapTableVal29.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable14)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable14


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable15 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal30;
	rand uvm_reg_field AcsmMapTableVal31;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal30: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal31: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable15");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal30 = uvm_reg_field::type_id::create("AcsmMapTableVal30",,get_full_name());
      this.AcsmMapTableVal30.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal31 = uvm_reg_field::type_id::create("AcsmMapTableVal31",,get_full_name());
      this.AcsmMapTableVal31.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable15)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable15


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable16 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal32;
	rand uvm_reg_field AcsmMapTableVal33;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal32: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal33: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable16");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal32 = uvm_reg_field::type_id::create("AcsmMapTableVal32",,get_full_name());
      this.AcsmMapTableVal32.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal33 = uvm_reg_field::type_id::create("AcsmMapTableVal33",,get_full_name());
      this.AcsmMapTableVal33.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable16)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable16


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable17 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal34;
	rand uvm_reg_field AcsmMapTableVal35;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal34: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal35: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable17");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal34 = uvm_reg_field::type_id::create("AcsmMapTableVal34",,get_full_name());
      this.AcsmMapTableVal34.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal35 = uvm_reg_field::type_id::create("AcsmMapTableVal35",,get_full_name());
      this.AcsmMapTableVal35.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable17)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable17


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable18 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal36;
	rand uvm_reg_field AcsmMapTableVal37;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal36: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal37: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable18");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal36 = uvm_reg_field::type_id::create("AcsmMapTableVal36",,get_full_name());
      this.AcsmMapTableVal36.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal37 = uvm_reg_field::type_id::create("AcsmMapTableVal37",,get_full_name());
      this.AcsmMapTableVal37.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable18)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable18


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable19 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal38;
	rand uvm_reg_field AcsmMapTableVal39;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal38: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal39: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable19");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal38 = uvm_reg_field::type_id::create("AcsmMapTableVal38",,get_full_name());
      this.AcsmMapTableVal38.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal39 = uvm_reg_field::type_id::create("AcsmMapTableVal39",,get_full_name());
      this.AcsmMapTableVal39.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable19)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable19


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable20 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal40;
	rand uvm_reg_field AcsmMapTableVal41;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal40: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal41: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable20");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal40 = uvm_reg_field::type_id::create("AcsmMapTableVal40",,get_full_name());
      this.AcsmMapTableVal40.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal41 = uvm_reg_field::type_id::create("AcsmMapTableVal41",,get_full_name());
      this.AcsmMapTableVal41.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable20)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable20


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable21 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal42;
	rand uvm_reg_field AcsmMapTableVal43;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal42: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal43: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable21");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal42 = uvm_reg_field::type_id::create("AcsmMapTableVal42",,get_full_name());
      this.AcsmMapTableVal42.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal43 = uvm_reg_field::type_id::create("AcsmMapTableVal43",,get_full_name());
      this.AcsmMapTableVal43.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable21)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable21


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable22 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal44;
	rand uvm_reg_field AcsmMapTableVal45;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal44: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal45: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable22");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal44 = uvm_reg_field::type_id::create("AcsmMapTableVal44",,get_full_name());
      this.AcsmMapTableVal44.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal45 = uvm_reg_field::type_id::create("AcsmMapTableVal45",,get_full_name());
      this.AcsmMapTableVal45.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable22)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable22


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable23 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal46;
	rand uvm_reg_field AcsmMapTableVal47;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal46: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal47: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable23");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal46 = uvm_reg_field::type_id::create("AcsmMapTableVal46",,get_full_name());
      this.AcsmMapTableVal46.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal47 = uvm_reg_field::type_id::create("AcsmMapTableVal47",,get_full_name());
      this.AcsmMapTableVal47.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable23)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable23


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable24 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal48;
	rand uvm_reg_field AcsmMapTableVal49;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal48: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal49: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable24");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal48 = uvm_reg_field::type_id::create("AcsmMapTableVal48",,get_full_name());
      this.AcsmMapTableVal48.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal49 = uvm_reg_field::type_id::create("AcsmMapTableVal49",,get_full_name());
      this.AcsmMapTableVal49.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable24)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable24


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable25 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal50;
	rand uvm_reg_field AcsmMapTableVal51;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal50: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal51: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable25");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal50 = uvm_reg_field::type_id::create("AcsmMapTableVal50",,get_full_name());
      this.AcsmMapTableVal50.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal51 = uvm_reg_field::type_id::create("AcsmMapTableVal51",,get_full_name());
      this.AcsmMapTableVal51.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable25)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable25


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable26 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal52;
	rand uvm_reg_field AcsmMapTableVal53;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal52: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal53: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable26");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal52 = uvm_reg_field::type_id::create("AcsmMapTableVal52",,get_full_name());
      this.AcsmMapTableVal52.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal53 = uvm_reg_field::type_id::create("AcsmMapTableVal53",,get_full_name());
      this.AcsmMapTableVal53.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable26)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable26


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable27 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal54;
	rand uvm_reg_field AcsmMapTableVal55;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal54: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal55: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable27");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal54 = uvm_reg_field::type_id::create("AcsmMapTableVal54",,get_full_name());
      this.AcsmMapTableVal54.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal55 = uvm_reg_field::type_id::create("AcsmMapTableVal55",,get_full_name());
      this.AcsmMapTableVal55.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable27)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable27


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable28 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal56;
	rand uvm_reg_field AcsmMapTableVal57;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal56: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal57: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable28");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal56 = uvm_reg_field::type_id::create("AcsmMapTableVal56",,get_full_name());
      this.AcsmMapTableVal56.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal57 = uvm_reg_field::type_id::create("AcsmMapTableVal57",,get_full_name());
      this.AcsmMapTableVal57.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable28)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable28


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable29 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal58;
	rand uvm_reg_field AcsmMapTableVal59;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal58: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal59: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable29");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal58 = uvm_reg_field::type_id::create("AcsmMapTableVal58",,get_full_name());
      this.AcsmMapTableVal58.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal59 = uvm_reg_field::type_id::create("AcsmMapTableVal59",,get_full_name());
      this.AcsmMapTableVal59.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable29)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable29


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable30 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal60;
	rand uvm_reg_field AcsmMapTableVal61;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal60: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal61: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable30");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal60 = uvm_reg_field::type_id::create("AcsmMapTableVal60",,get_full_name());
      this.AcsmMapTableVal60.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal61 = uvm_reg_field::type_id::create("AcsmMapTableVal61",,get_full_name());
      this.AcsmMapTableVal61.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable30)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable30


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable31 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal62;
	rand uvm_reg_field AcsmMapTableVal63;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal62: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal63: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable31");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal62 = uvm_reg_field::type_id::create("AcsmMapTableVal62",,get_full_name());
      this.AcsmMapTableVal62.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal63 = uvm_reg_field::type_id::create("AcsmMapTableVal63",,get_full_name());
      this.AcsmMapTableVal63.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable31)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable31


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable32 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal64;
	rand uvm_reg_field AcsmMapTableVal65;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal64: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal65: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable32");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal64 = uvm_reg_field::type_id::create("AcsmMapTableVal64",,get_full_name());
      this.AcsmMapTableVal64.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal65 = uvm_reg_field::type_id::create("AcsmMapTableVal65",,get_full_name());
      this.AcsmMapTableVal65.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable32)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable32


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable33 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal66;
	rand uvm_reg_field AcsmMapTableVal67;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal66: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal67: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable33");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal66 = uvm_reg_field::type_id::create("AcsmMapTableVal66",,get_full_name());
      this.AcsmMapTableVal66.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal67 = uvm_reg_field::type_id::create("AcsmMapTableVal67",,get_full_name());
      this.AcsmMapTableVal67.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable33)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable33


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable34 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal68;
	rand uvm_reg_field AcsmMapTableVal69;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal68: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal69: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable34");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal68 = uvm_reg_field::type_id::create("AcsmMapTableVal68",,get_full_name());
      this.AcsmMapTableVal68.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal69 = uvm_reg_field::type_id::create("AcsmMapTableVal69",,get_full_name());
      this.AcsmMapTableVal69.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable34)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable34


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable35 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal70;
	rand uvm_reg_field AcsmMapTableVal71;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal70: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal71: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable35");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal70 = uvm_reg_field::type_id::create("AcsmMapTableVal70",,get_full_name());
      this.AcsmMapTableVal70.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal71 = uvm_reg_field::type_id::create("AcsmMapTableVal71",,get_full_name());
      this.AcsmMapTableVal71.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable35)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable35


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable36 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal72;
	rand uvm_reg_field AcsmMapTableVal73;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal72: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal73: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable36");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal72 = uvm_reg_field::type_id::create("AcsmMapTableVal72",,get_full_name());
      this.AcsmMapTableVal72.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal73 = uvm_reg_field::type_id::create("AcsmMapTableVal73",,get_full_name());
      this.AcsmMapTableVal73.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable36)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable36


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable37 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal74;
	rand uvm_reg_field AcsmMapTableVal75;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal74: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal75: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable37");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal74 = uvm_reg_field::type_id::create("AcsmMapTableVal74",,get_full_name());
      this.AcsmMapTableVal74.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal75 = uvm_reg_field::type_id::create("AcsmMapTableVal75",,get_full_name());
      this.AcsmMapTableVal75.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable37)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable37


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable38 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal76;
	rand uvm_reg_field AcsmMapTableVal77;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal76: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal77: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable38");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal76 = uvm_reg_field::type_id::create("AcsmMapTableVal76",,get_full_name());
      this.AcsmMapTableVal76.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal77 = uvm_reg_field::type_id::create("AcsmMapTableVal77",,get_full_name());
      this.AcsmMapTableVal77.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable38)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable38


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable39 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal78;
	rand uvm_reg_field AcsmMapTableVal79;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal78: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal79: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable39");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal78 = uvm_reg_field::type_id::create("AcsmMapTableVal78",,get_full_name());
      this.AcsmMapTableVal78.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal79 = uvm_reg_field::type_id::create("AcsmMapTableVal79",,get_full_name());
      this.AcsmMapTableVal79.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable39)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable39


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable40 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal80;
	rand uvm_reg_field AcsmMapTableVal81;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal80: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal81: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable40");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal80 = uvm_reg_field::type_id::create("AcsmMapTableVal80",,get_full_name());
      this.AcsmMapTableVal80.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal81 = uvm_reg_field::type_id::create("AcsmMapTableVal81",,get_full_name());
      this.AcsmMapTableVal81.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable40)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable40


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable41 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal82;
	rand uvm_reg_field AcsmMapTableVal83;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal82: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal83: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable41");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal82 = uvm_reg_field::type_id::create("AcsmMapTableVal82",,get_full_name());
      this.AcsmMapTableVal82.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal83 = uvm_reg_field::type_id::create("AcsmMapTableVal83",,get_full_name());
      this.AcsmMapTableVal83.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable41)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable41


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable42 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal84;
	rand uvm_reg_field AcsmMapTableVal85;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal84: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal85: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable42");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal84 = uvm_reg_field::type_id::create("AcsmMapTableVal84",,get_full_name());
      this.AcsmMapTableVal84.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal85 = uvm_reg_field::type_id::create("AcsmMapTableVal85",,get_full_name());
      this.AcsmMapTableVal85.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable42)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable42


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable43 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal86;
	rand uvm_reg_field AcsmMapTableVal87;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal86: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal87: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable43");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal86 = uvm_reg_field::type_id::create("AcsmMapTableVal86",,get_full_name());
      this.AcsmMapTableVal86.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal87 = uvm_reg_field::type_id::create("AcsmMapTableVal87",,get_full_name());
      this.AcsmMapTableVal87.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable43)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable43


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable44 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal88;
	rand uvm_reg_field AcsmMapTableVal89;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal88: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal89: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable44");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal88 = uvm_reg_field::type_id::create("AcsmMapTableVal88",,get_full_name());
      this.AcsmMapTableVal88.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal89 = uvm_reg_field::type_id::create("AcsmMapTableVal89",,get_full_name());
      this.AcsmMapTableVal89.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable44)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable44


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable45 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal90;
	rand uvm_reg_field AcsmMapTableVal91;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal90: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal91: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable45");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal90 = uvm_reg_field::type_id::create("AcsmMapTableVal90",,get_full_name());
      this.AcsmMapTableVal90.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal91 = uvm_reg_field::type_id::create("AcsmMapTableVal91",,get_full_name());
      this.AcsmMapTableVal91.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable45)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable45


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable46 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal92;
	rand uvm_reg_field AcsmMapTableVal93;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal92: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal93: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable46");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal92 = uvm_reg_field::type_id::create("AcsmMapTableVal92",,get_full_name());
      this.AcsmMapTableVal92.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal93 = uvm_reg_field::type_id::create("AcsmMapTableVal93",,get_full_name());
      this.AcsmMapTableVal93.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable46)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable46


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable47 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal94;
	rand uvm_reg_field AcsmMapTableVal95;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal94: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal95: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable47");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal94 = uvm_reg_field::type_id::create("AcsmMapTableVal94",,get_full_name());
      this.AcsmMapTableVal94.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal95 = uvm_reg_field::type_id::create("AcsmMapTableVal95",,get_full_name());
      this.AcsmMapTableVal95.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable47)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable47


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable48 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal96;
	rand uvm_reg_field AcsmMapTableVal97;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal96: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal97: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable48");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal96 = uvm_reg_field::type_id::create("AcsmMapTableVal96",,get_full_name());
      this.AcsmMapTableVal96.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal97 = uvm_reg_field::type_id::create("AcsmMapTableVal97",,get_full_name());
      this.AcsmMapTableVal97.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable48)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable48


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable49 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal98;
	rand uvm_reg_field AcsmMapTableVal99;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal98: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal99: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable49");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal98 = uvm_reg_field::type_id::create("AcsmMapTableVal98",,get_full_name());
      this.AcsmMapTableVal98.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal99 = uvm_reg_field::type_id::create("AcsmMapTableVal99",,get_full_name());
      this.AcsmMapTableVal99.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable49)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable49


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable50 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal100;
	rand uvm_reg_field AcsmMapTableVal101;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal100: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal101: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable50");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal100 = uvm_reg_field::type_id::create("AcsmMapTableVal100",,get_full_name());
      this.AcsmMapTableVal100.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal101 = uvm_reg_field::type_id::create("AcsmMapTableVal101",,get_full_name());
      this.AcsmMapTableVal101.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable50)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable50


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable51 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal102;
	rand uvm_reg_field AcsmMapTableVal103;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal102: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal103: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable51");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal102 = uvm_reg_field::type_id::create("AcsmMapTableVal102",,get_full_name());
      this.AcsmMapTableVal102.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal103 = uvm_reg_field::type_id::create("AcsmMapTableVal103",,get_full_name());
      this.AcsmMapTableVal103.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable51)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable51


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable52 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal104;
	rand uvm_reg_field AcsmMapTableVal105;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal104: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal105: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable52");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal104 = uvm_reg_field::type_id::create("AcsmMapTableVal104",,get_full_name());
      this.AcsmMapTableVal104.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal105 = uvm_reg_field::type_id::create("AcsmMapTableVal105",,get_full_name());
      this.AcsmMapTableVal105.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable52)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable52


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable53 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal106;
	rand uvm_reg_field AcsmMapTableVal107;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal106: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal107: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable53");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal106 = uvm_reg_field::type_id::create("AcsmMapTableVal106",,get_full_name());
      this.AcsmMapTableVal106.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal107 = uvm_reg_field::type_id::create("AcsmMapTableVal107",,get_full_name());
      this.AcsmMapTableVal107.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable53)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable53


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable54 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal108;
	rand uvm_reg_field AcsmMapTableVal109;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal108: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal109: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable54");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal108 = uvm_reg_field::type_id::create("AcsmMapTableVal108",,get_full_name());
      this.AcsmMapTableVal108.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal109 = uvm_reg_field::type_id::create("AcsmMapTableVal109",,get_full_name());
      this.AcsmMapTableVal109.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable54)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable54


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable55 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal110;
	rand uvm_reg_field AcsmMapTableVal111;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal110: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal111: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable55");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal110 = uvm_reg_field::type_id::create("AcsmMapTableVal110",,get_full_name());
      this.AcsmMapTableVal110.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal111 = uvm_reg_field::type_id::create("AcsmMapTableVal111",,get_full_name());
      this.AcsmMapTableVal111.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable55)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable55


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable56 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal112;
	rand uvm_reg_field AcsmMapTableVal113;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal112: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal113: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable56");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal112 = uvm_reg_field::type_id::create("AcsmMapTableVal112",,get_full_name());
      this.AcsmMapTableVal112.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal113 = uvm_reg_field::type_id::create("AcsmMapTableVal113",,get_full_name());
      this.AcsmMapTableVal113.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable56)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable56


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable57 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal114;
	rand uvm_reg_field AcsmMapTableVal115;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal114: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal115: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable57");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal114 = uvm_reg_field::type_id::create("AcsmMapTableVal114",,get_full_name());
      this.AcsmMapTableVal114.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal115 = uvm_reg_field::type_id::create("AcsmMapTableVal115",,get_full_name());
      this.AcsmMapTableVal115.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable57)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable57


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable58 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal116;
	rand uvm_reg_field AcsmMapTableVal117;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal116: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal117: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable58");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal116 = uvm_reg_field::type_id::create("AcsmMapTableVal116",,get_full_name());
      this.AcsmMapTableVal116.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal117 = uvm_reg_field::type_id::create("AcsmMapTableVal117",,get_full_name());
      this.AcsmMapTableVal117.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable58)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable58


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable59 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal118;
	rand uvm_reg_field AcsmMapTableVal119;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal118: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal119: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable59");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal118 = uvm_reg_field::type_id::create("AcsmMapTableVal118",,get_full_name());
      this.AcsmMapTableVal118.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal119 = uvm_reg_field::type_id::create("AcsmMapTableVal119",,get_full_name());
      this.AcsmMapTableVal119.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable59)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable59


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable60 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal120;
	rand uvm_reg_field AcsmMapTableVal121;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal120: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal121: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable60");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal120 = uvm_reg_field::type_id::create("AcsmMapTableVal120",,get_full_name());
      this.AcsmMapTableVal120.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal121 = uvm_reg_field::type_id::create("AcsmMapTableVal121",,get_full_name());
      this.AcsmMapTableVal121.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable60)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable60


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable61 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal122;
	rand uvm_reg_field AcsmMapTableVal123;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal122: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal123: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable61");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal122 = uvm_reg_field::type_id::create("AcsmMapTableVal122",,get_full_name());
      this.AcsmMapTableVal122.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal123 = uvm_reg_field::type_id::create("AcsmMapTableVal123",,get_full_name());
      this.AcsmMapTableVal123.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable61)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable61


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable62 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal124;
	rand uvm_reg_field AcsmMapTableVal125;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal124: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal125: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable62");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal124 = uvm_reg_field::type_id::create("AcsmMapTableVal124",,get_full_name());
      this.AcsmMapTableVal124.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal125 = uvm_reg_field::type_id::create("AcsmMapTableVal125",,get_full_name());
      this.AcsmMapTableVal125.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable62)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable62


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable63 extends uvm_reg;
	rand uvm_reg_field AcsmMapTableVal126;
	rand uvm_reg_field AcsmMapTableVal127;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmMapTableVal126: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	   AcsmMapTableVal127: coverpoint {m_data[11:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmMapTable63");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmMapTableVal126 = uvm_reg_field::type_id::create("AcsmMapTableVal126",,get_full_name());
      this.AcsmMapTableVal126.configure(this, 6, 0, "RW", 0, 6'h0, 1, 0, 0);
      this.AcsmMapTableVal127 = uvm_reg_field::type_id::create("AcsmMapTableVal127",,get_full_name());
      this.AcsmMapTableVal127.configure(this, 6, 6, "RW", 0, 6'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable63)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable63


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal0 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal0: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal0 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal0",,get_full_name());
      this.AcsmStartAddrXlatVal0.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal1 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal1 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal1",,get_full_name());
      this.AcsmStartAddrXlatVal1.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal2 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal2: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal2");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal2 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal2",,get_full_name());
      this.AcsmStartAddrXlatVal2.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal2)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal2


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal3 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal3;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal3: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal3");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal3 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal3",,get_full_name());
      this.AcsmStartAddrXlatVal3.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal3)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal3


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal4 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal4;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal4: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal4");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal4 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal4",,get_full_name());
      this.AcsmStartAddrXlatVal4.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal4)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal4


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal5 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal5;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal5: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal5");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal5 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal5",,get_full_name());
      this.AcsmStartAddrXlatVal5.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal5)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal5


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal6 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal6;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal6: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal6");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal6 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal6",,get_full_name());
      this.AcsmStartAddrXlatVal6.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal6)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal6


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal7 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal7;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal7: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal7");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal7 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal7",,get_full_name());
      this.AcsmStartAddrXlatVal7.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal7)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal7


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal8 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal8;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal8: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal8");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal8 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal8",,get_full_name());
      this.AcsmStartAddrXlatVal8.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal8)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal8


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal9 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal9;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal9: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal9");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal9 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal9",,get_full_name());
      this.AcsmStartAddrXlatVal9.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal9)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal9


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal10 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal10;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal10: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal10");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal10 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal10",,get_full_name());
      this.AcsmStartAddrXlatVal10.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal10)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal10


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal11 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal11;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal11: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal11");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal11 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal11",,get_full_name());
      this.AcsmStartAddrXlatVal11.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal11)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal11


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal12 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal12;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal12: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal12");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal12 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal12",,get_full_name());
      this.AcsmStartAddrXlatVal12.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal12)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal12


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal13 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal13;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal13: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal13");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal13 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal13",,get_full_name());
      this.AcsmStartAddrXlatVal13.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal13)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal13


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal14 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal14;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal14: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal14");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal14 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal14",,get_full_name());
      this.AcsmStartAddrXlatVal14.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal14)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal14


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal15 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal15;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal15: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal15");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal15 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal15",,get_full_name());
      this.AcsmStartAddrXlatVal15.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal15)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal15


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal16 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal16;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal16: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal16");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal16 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal16",,get_full_name());
      this.AcsmStartAddrXlatVal16.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal16)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal16


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal17 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal17;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal17: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal17");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal17 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal17",,get_full_name());
      this.AcsmStartAddrXlatVal17.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal17)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal17


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal18 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal18;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal18: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal18");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal18 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal18",,get_full_name());
      this.AcsmStartAddrXlatVal18.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal18)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal18


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal19 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal19;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal19: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal19");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal19 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal19",,get_full_name());
      this.AcsmStartAddrXlatVal19.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal19)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal19


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal20 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal20;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal20: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal20");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal20 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal20",,get_full_name());
      this.AcsmStartAddrXlatVal20.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal20)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal20


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal21 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal21;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal21: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal21");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal21 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal21",,get_full_name());
      this.AcsmStartAddrXlatVal21.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal21)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal21


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal22 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal22;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal22: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal22");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal22 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal22",,get_full_name());
      this.AcsmStartAddrXlatVal22.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal22)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal22


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal23 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal23;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal23: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal23");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal23 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal23",,get_full_name());
      this.AcsmStartAddrXlatVal23.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal23)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal23


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal24 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal24;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal24: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal24");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal24 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal24",,get_full_name());
      this.AcsmStartAddrXlatVal24.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal24)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal24


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal25 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal25;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal25: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal25");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal25 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal25",,get_full_name());
      this.AcsmStartAddrXlatVal25.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal25)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal25


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal26 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal26;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal26: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal26");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal26 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal26",,get_full_name());
      this.AcsmStartAddrXlatVal26.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal26)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal26


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal27 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal27;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal27: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal27");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal27 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal27",,get_full_name());
      this.AcsmStartAddrXlatVal27.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal27)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal27


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal28 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal28;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal28: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal28");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal28 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal28",,get_full_name());
      this.AcsmStartAddrXlatVal28.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal28)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal28


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal29 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal29;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal29: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal29");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal29 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal29",,get_full_name());
      this.AcsmStartAddrXlatVal29.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal29)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal29


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal30 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal30;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal30: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal30");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal30 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal30",,get_full_name());
      this.AcsmStartAddrXlatVal30.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal30)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal30


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal31 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal31;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal31: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal31");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal31 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal31",,get_full_name());
      this.AcsmStartAddrXlatVal31.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal31)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal31


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal32 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal32;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal32: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal32");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal32 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal32",,get_full_name());
      this.AcsmStartAddrXlatVal32.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal32)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal32


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal33 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal33;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal33: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal33");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal33 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal33",,get_full_name());
      this.AcsmStartAddrXlatVal33.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal33)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal33


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal34 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal34;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal34: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal34");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal34 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal34",,get_full_name());
      this.AcsmStartAddrXlatVal34.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal34)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal34


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal35 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal35;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal35: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal35");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal35 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal35",,get_full_name());
      this.AcsmStartAddrXlatVal35.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal35)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal35


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal36 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal36;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal36: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal36");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal36 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal36",,get_full_name());
      this.AcsmStartAddrXlatVal36.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal36)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal36


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal37 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal37;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal37: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal37");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal37 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal37",,get_full_name());
      this.AcsmStartAddrXlatVal37.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal37)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal37


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal38 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal38;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal38: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal38");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal38 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal38",,get_full_name());
      this.AcsmStartAddrXlatVal38.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal38)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal38


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal39 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal39;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal39: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal39");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal39 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal39",,get_full_name());
      this.AcsmStartAddrXlatVal39.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal39)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal39


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal40 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal40;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal40: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal40");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal40 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal40",,get_full_name());
      this.AcsmStartAddrXlatVal40.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal40)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal40


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal41 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal41;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal41: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal41");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal41 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal41",,get_full_name());
      this.AcsmStartAddrXlatVal41.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal41)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal41


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal42 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal42;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal42: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal42");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal42 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal42",,get_full_name());
      this.AcsmStartAddrXlatVal42.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal42)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal42


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal43 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal43;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal43: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal43");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal43 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal43",,get_full_name());
      this.AcsmStartAddrXlatVal43.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal43)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal43


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal44 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal44;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal44: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal44");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal44 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal44",,get_full_name());
      this.AcsmStartAddrXlatVal44.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal44)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal44


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal45 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal45;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal45: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal45");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal45 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal45",,get_full_name());
      this.AcsmStartAddrXlatVal45.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal45)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal45


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal46 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal46;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal46: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal46");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal46 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal46",,get_full_name());
      this.AcsmStartAddrXlatVal46.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal46)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal46


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal47 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal47;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal47: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal47");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal47 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal47",,get_full_name());
      this.AcsmStartAddrXlatVal47.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal47)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal47


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal48 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal48;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal48: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal48");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal48 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal48",,get_full_name());
      this.AcsmStartAddrXlatVal48.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal48)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal48


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal49 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal49;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal49: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal49");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal49 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal49",,get_full_name());
      this.AcsmStartAddrXlatVal49.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal49)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal49


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal50 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal50;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal50: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal50");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal50 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal50",,get_full_name());
      this.AcsmStartAddrXlatVal50.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal50)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal50


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal51 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal51;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal51: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal51");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal51 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal51",,get_full_name());
      this.AcsmStartAddrXlatVal51.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal51)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal51


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal52 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal52;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal52: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal52");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal52 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal52",,get_full_name());
      this.AcsmStartAddrXlatVal52.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal52)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal52


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal53 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal53;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal53: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal53");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal53 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal53",,get_full_name());
      this.AcsmStartAddrXlatVal53.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal53)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal53


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal54 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal54;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal54: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal54");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal54 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal54",,get_full_name());
      this.AcsmStartAddrXlatVal54.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal54)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal54


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal55 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal55;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal55: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal55");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal55 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal55",,get_full_name());
      this.AcsmStartAddrXlatVal55.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal55)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal55


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal56 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal56;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal56: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal56");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal56 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal56",,get_full_name());
      this.AcsmStartAddrXlatVal56.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal56)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal56


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal57 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal57;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal57: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal57");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal57 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal57",,get_full_name());
      this.AcsmStartAddrXlatVal57.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal57)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal57


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal58 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal58;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal58: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal58");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal58 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal58",,get_full_name());
      this.AcsmStartAddrXlatVal58.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal58)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal58


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal59 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal59;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal59: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal59");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal59 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal59",,get_full_name());
      this.AcsmStartAddrXlatVal59.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal59)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal59


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal60 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal60;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal60: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal60");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal60 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal60",,get_full_name());
      this.AcsmStartAddrXlatVal60.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal60)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal60


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal61 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal61;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal61: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal61");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal61 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal61",,get_full_name());
      this.AcsmStartAddrXlatVal61.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal61)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal61


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal62 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal62;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal62: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal62");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal62 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal62",,get_full_name());
      this.AcsmStartAddrXlatVal62.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal62)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal62


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal63 extends uvm_reg;
	rand uvm_reg_field AcsmStartAddrXlatVal63;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStartAddrXlatVal63: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal63");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStartAddrXlatVal63 = uvm_reg_field::type_id::create("AcsmStartAddrXlatVal63",,get_full_name());
      this.AcsmStartAddrXlatVal63.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal63)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal63


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal0 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal0: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal0");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal0 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal0",,get_full_name());
      this.AcsmStopAddrXlatVal0.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal0


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal1 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal1 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal1",,get_full_name());
      this.AcsmStopAddrXlatVal1.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal1


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal2 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal2: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal2");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal2 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal2",,get_full_name());
      this.AcsmStopAddrXlatVal2.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal2)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal2


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal3 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal3;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal3: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal3");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal3 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal3",,get_full_name());
      this.AcsmStopAddrXlatVal3.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal3)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal3


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal4 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal4;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal4: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal4");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal4 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal4",,get_full_name());
      this.AcsmStopAddrXlatVal4.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal4)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal4


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal5 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal5;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal5: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal5");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal5 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal5",,get_full_name());
      this.AcsmStopAddrXlatVal5.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal5)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal5


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal6 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal6;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal6: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal6");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal6 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal6",,get_full_name());
      this.AcsmStopAddrXlatVal6.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal6)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal6


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal7 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal7;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal7: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal7");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal7 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal7",,get_full_name());
      this.AcsmStopAddrXlatVal7.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal7)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal7


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal8 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal8;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal8: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal8");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal8 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal8",,get_full_name());
      this.AcsmStopAddrXlatVal8.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal8)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal8


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal9 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal9;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal9: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal9");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal9 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal9",,get_full_name());
      this.AcsmStopAddrXlatVal9.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal9)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal9


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal10 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal10;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal10: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal10");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal10 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal10",,get_full_name());
      this.AcsmStopAddrXlatVal10.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal10)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal10


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal11 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal11;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal11: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal11");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal11 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal11",,get_full_name());
      this.AcsmStopAddrXlatVal11.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal11)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal11


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal12 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal12;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal12: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal12");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal12 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal12",,get_full_name());
      this.AcsmStopAddrXlatVal12.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal12)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal12


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal13 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal13;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal13: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal13");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal13 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal13",,get_full_name());
      this.AcsmStopAddrXlatVal13.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal13)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal13


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal14 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal14;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal14: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal14");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal14 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal14",,get_full_name());
      this.AcsmStopAddrXlatVal14.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal14)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal14


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal15 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal15;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal15: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal15");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal15 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal15",,get_full_name());
      this.AcsmStopAddrXlatVal15.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal15)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal15


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal16 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal16;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal16: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal16");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal16 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal16",,get_full_name());
      this.AcsmStopAddrXlatVal16.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal16)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal16


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal17 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal17;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal17: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal17");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal17 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal17",,get_full_name());
      this.AcsmStopAddrXlatVal17.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal17)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal17


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal18 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal18;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal18: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal18");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal18 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal18",,get_full_name());
      this.AcsmStopAddrXlatVal18.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal18)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal18


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal19 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal19;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal19: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal19");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal19 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal19",,get_full_name());
      this.AcsmStopAddrXlatVal19.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal19)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal19


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal20 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal20;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal20: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal20");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal20 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal20",,get_full_name());
      this.AcsmStopAddrXlatVal20.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal20)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal20


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal21 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal21;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal21: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal21");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal21 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal21",,get_full_name());
      this.AcsmStopAddrXlatVal21.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal21)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal21


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal22 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal22;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal22: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal22");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal22 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal22",,get_full_name());
      this.AcsmStopAddrXlatVal22.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal22)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal22


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal23 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal23;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal23: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal23");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal23 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal23",,get_full_name());
      this.AcsmStopAddrXlatVal23.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal23)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal23


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal24 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal24;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal24: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal24");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal24 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal24",,get_full_name());
      this.AcsmStopAddrXlatVal24.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal24)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal24


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal25 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal25;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal25: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal25");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal25 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal25",,get_full_name());
      this.AcsmStopAddrXlatVal25.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal25)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal25


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal26 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal26;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal26: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal26");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal26 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal26",,get_full_name());
      this.AcsmStopAddrXlatVal26.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal26)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal26


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal27 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal27;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal27: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal27");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal27 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal27",,get_full_name());
      this.AcsmStopAddrXlatVal27.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal27)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal27


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal28 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal28;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal28: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal28");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal28 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal28",,get_full_name());
      this.AcsmStopAddrXlatVal28.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal28)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal28


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal29 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal29;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal29: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal29");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal29 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal29",,get_full_name());
      this.AcsmStopAddrXlatVal29.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal29)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal29


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal30 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal30;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal30: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal30");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal30 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal30",,get_full_name());
      this.AcsmStopAddrXlatVal30.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal30)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal30


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal31 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal31;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal31: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal31");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal31 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal31",,get_full_name());
      this.AcsmStopAddrXlatVal31.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal31)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal31


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal32 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal32;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal32: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal32");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal32 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal32",,get_full_name());
      this.AcsmStopAddrXlatVal32.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal32)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal32


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal33 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal33;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal33: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal33");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal33 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal33",,get_full_name());
      this.AcsmStopAddrXlatVal33.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal33)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal33


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal34 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal34;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal34: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal34");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal34 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal34",,get_full_name());
      this.AcsmStopAddrXlatVal34.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal34)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal34


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal35 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal35;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal35: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal35");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal35 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal35",,get_full_name());
      this.AcsmStopAddrXlatVal35.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal35)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal35


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal36 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal36;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal36: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal36");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal36 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal36",,get_full_name());
      this.AcsmStopAddrXlatVal36.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal36)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal36


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal37 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal37;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal37: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal37");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal37 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal37",,get_full_name());
      this.AcsmStopAddrXlatVal37.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal37)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal37


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal38 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal38;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal38: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal38");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal38 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal38",,get_full_name());
      this.AcsmStopAddrXlatVal38.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal38)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal38


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal39 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal39;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal39: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal39");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal39 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal39",,get_full_name());
      this.AcsmStopAddrXlatVal39.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal39)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal39


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal40 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal40;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal40: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal40");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal40 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal40",,get_full_name());
      this.AcsmStopAddrXlatVal40.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal40)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal40


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal41 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal41;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal41: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal41");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal41 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal41",,get_full_name());
      this.AcsmStopAddrXlatVal41.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal41)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal41


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal42 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal42;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal42: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal42");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal42 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal42",,get_full_name());
      this.AcsmStopAddrXlatVal42.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal42)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal42


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal43 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal43;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal43: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal43");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal43 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal43",,get_full_name());
      this.AcsmStopAddrXlatVal43.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal43)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal43


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal44 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal44;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal44: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal44");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal44 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal44",,get_full_name());
      this.AcsmStopAddrXlatVal44.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal44)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal44


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal45 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal45;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal45: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal45");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal45 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal45",,get_full_name());
      this.AcsmStopAddrXlatVal45.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal45)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal45


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal46 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal46;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal46: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal46");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal46 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal46",,get_full_name());
      this.AcsmStopAddrXlatVal46.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal46)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal46


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal47 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal47;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal47: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal47");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal47 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal47",,get_full_name());
      this.AcsmStopAddrXlatVal47.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal47)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal47


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal48 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal48;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal48: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal48");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal48 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal48",,get_full_name());
      this.AcsmStopAddrXlatVal48.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal48)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal48


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal49 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal49;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal49: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal49");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal49 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal49",,get_full_name());
      this.AcsmStopAddrXlatVal49.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal49)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal49


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal50 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal50;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal50: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal50");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal50 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal50",,get_full_name());
      this.AcsmStopAddrXlatVal50.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal50)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal50


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal51 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal51;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal51: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal51");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal51 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal51",,get_full_name());
      this.AcsmStopAddrXlatVal51.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal51)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal51


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal52 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal52;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal52: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal52");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal52 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal52",,get_full_name());
      this.AcsmStopAddrXlatVal52.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal52)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal52


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal53 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal53;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal53: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal53");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal53 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal53",,get_full_name());
      this.AcsmStopAddrXlatVal53.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal53)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal53


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal54 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal54;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal54: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal54");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal54 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal54",,get_full_name());
      this.AcsmStopAddrXlatVal54.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal54)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal54


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal55 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal55;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal55: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal55");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal55 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal55",,get_full_name());
      this.AcsmStopAddrXlatVal55.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal55)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal55


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal56 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal56;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal56: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal56");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal56 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal56",,get_full_name());
      this.AcsmStopAddrXlatVal56.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal56)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal56


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal57 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal57;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal57: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal57");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal57 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal57",,get_full_name());
      this.AcsmStopAddrXlatVal57.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal57)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal57


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal58 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal58;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal58: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal58");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal58 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal58",,get_full_name());
      this.AcsmStopAddrXlatVal58.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal58)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal58


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal59 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal59;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal59: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal59");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal59 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal59",,get_full_name());
      this.AcsmStopAddrXlatVal59.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal59)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal59


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal60 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal60;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal60: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal60");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal60 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal60",,get_full_name());
      this.AcsmStopAddrXlatVal60.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal60)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal60


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal61 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal61;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal61: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal61");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal61 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal61",,get_full_name());
      this.AcsmStopAddrXlatVal61.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal61)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal61


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal62 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal62;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal62: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal62");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal62 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal62",,get_full_name());
      this.AcsmStopAddrXlatVal62.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal62)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal62


class ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal63 extends uvm_reg;
	rand uvm_reg_field AcsmStopAddrXlatVal63;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   AcsmStopAddrXlatVal63: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal63");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.AcsmStopAddrXlatVal63 = uvm_reg_field::type_id::create("AcsmStopAddrXlatVal63",,get_full_name());
      this.AcsmStopAddrXlatVal63.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal63)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal63


class ral_block_DWC_DDRPHYA_PPGC0_p0 extends uvm_reg_block;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenCtrl PpgcGenCtrl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiCtrl PpgcGenDbiCtrl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiConfig PpgcGenDbiConfig;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel0 PpgcGenLaneMuxSel0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel1 PpgcGenLaneMuxSel1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_EnPhyUpdZQCalUpdate EnPhyUpdZQCalUpdate;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterface BlockDfiInterface;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterfaceStatus BlockDfiInterfaceStatus;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiCustMode_p0 DfiCustMode_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtMRL_p0 HwtMRL_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_RegRet RegRet;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DisableZQupdateOnSnoop DisableZQupdateOnSnoop;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenModeSel Prbs0GenModeSel;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenUiMuxSel Prbs0GenUiMuxSel;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly0 Prbs0GenTapDly0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly1 Prbs0GenTapDly1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly2 Prbs0GenTapDly2;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly3 Prbs0GenTapDly3;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly4 Prbs0GenTapDly4;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly5 Prbs0GenTapDly5;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly6 Prbs0GenTapDly6;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly7 Prbs0GenTapDly7;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_MtestMuxSel MtestMuxSel;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateLo Prbs0GenStateLo;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateHi Prbs0GenStateHi;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenModeSel Prbs1GenModeSel;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenUiMuxSel Prbs1GenUiMuxSel;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly0 Prbs1GenTapDly0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly1 Prbs1GenTapDly1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly2 Prbs1GenTapDly2;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly3 Prbs1GenTapDly3;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly4 Prbs1GenTapDly4;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly5 Prbs1GenTapDly5;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly6 Prbs1GenTapDly6;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly7 Prbs1GenTapDly7;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateLo Prbs1GenStateLo;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateHi Prbs1GenStateHi;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenModeSel Prbs2GenModeSel;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenUiMuxSel Prbs2GenUiMuxSel;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly0 Prbs2GenTapDly0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly1 Prbs2GenTapDly1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly2 Prbs2GenTapDly2;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly3 Prbs2GenTapDly3;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly4 Prbs2GenTapDly4;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly5 Prbs2GenTapDly5;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly6 Prbs2GenTapDly6;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly7 Prbs2GenTapDly7;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateLo Prbs2GenStateLo;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateHi Prbs2GenStateHi;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PPTTrainSetup_p0 PPTTrainSetup_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyMstrFreqOverride_p0 PhyMstrFreqOverride_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiInitComplete DfiInitComplete;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCParityInvert PPGCParityInvert;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PMIEnable PMIEnable;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi0Status Dfi0Status;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi1Status Dfi1Status;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays0_p0 DfiHandshakeDelays0_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD0 DFIPHYUPD0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn0 DfiLpCtrlEn0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn0 DfiLpDataEn0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl0 DynOdtEnCntrl0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays0_p0 DfiRespHandshakeDelays0_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnA HwtLpCsEnA;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnB HwtLpCsEnB;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtCtrl HwtCtrl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlOvr HwtControlOvr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ScratchPadPPGC ScratchPadPPGC;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlVal HwtControlVal;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ForceHWTClkGaterEnables ForceHWTClkGaterEnables;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdGoodCtr MasUpdGoodCtr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0GoodCtr PhyUpd0GoodCtr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1GoodCtr PhyUpd1GoodCtr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd0GoodCtr CtlUpd0GoodCtr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd1GoodCtr CtlUpd1GoodCtr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdFailCtr MasUpdFailCtr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0FailCtr PhyUpd0FailCtr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1FailCtr PhyUpd1FailCtr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyPerfCtrEnable PhyPerfCtrEnable;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays1_p0 DfiHandshakeDelays1_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD1 DFIPHYUPD1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn1 DfiLpCtrlEn1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn1 DfiLpDataEn1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl1 DynOdtEnCntrl1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays1_p0 DfiRespHandshakeDelays1_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_FspSkipList FspSkipList;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCReserved0 PPGCReserved0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PUBReservedP1_p0 PUBReservedP1_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptOverride PhyInterruptOverride;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptEnable PhyInterruptEnable;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptFWControl PhyInterruptFWControl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptMask PhyInterruptMask;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptClear PhyInterruptClear;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptStatus PhyInterruptStatus;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRunCtrl ACSMRunCtrl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDone ACSMDone;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStartAddr_p0 ACSMStartAddr_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStopAddr_p0 ACSMStopAddr_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLastAddr ACSMLastAddr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAlgaIncVal ACSMAlgaIncVal;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAddressMask ACSMAddressMask;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMOuterLoopRepeatCnt ACSMOuterLoopRepeatCnt;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeControl ACSMCkeControl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeStatus ACSMCkeStatus;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnControl ACSMWckEnControl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnStatus ACSMWckEnStatus;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxEnPulse_p0 ACSMRxEnPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxValPulse_p0 ACSMRxValPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMTxEnPulse_p0 ACSMTxEnPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWrcsPulse_p0 ACSMWrcsPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRdcsPulse_p0 ACSMRdcsPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMInfiniteOLRC ACSMInfiniteOLRC;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultAddr ACSMDefaultAddr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultCs ACSMDefaultCs;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStaticCtrl ACSMStaticCtrl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticLoPulse_p0 ACSMWckWriteStaticLoPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticHiPulse_p0 ACSMWckWriteStaticHiPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteTogglePulse_p0 ACSMWckWriteTogglePulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteFastTogglePulse_p0 ACSMWckWriteFastTogglePulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticLoPulse_p0 ACSMWckReadStaticLoPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticHiPulse_p0 ACSMWckReadStaticHiPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadTogglePulse_p0 ACSMWckReadTogglePulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadFastTogglePulse_p0 ACSMWckReadFastTogglePulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticLoPulse_p0 ACSMWckFreqSwStaticLoPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticHiPulse_p0 ACSMWckFreqSwStaticHiPulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwTogglePulse_p0 ACSMWckFreqSwTogglePulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwFastTogglePulse_p0 ACSMWckFreqSwFastTogglePulse_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreeRunMode_p0 ACSMWckFreeRunMode_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockEnable ACSMLowSpeedClockEnable;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockDelay ACSMLowSpeedClockDelay;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntOverride_p0 ACSMRptCntOverride_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntDbl_p0 ACSMRptCntDbl_p0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityStatus ACSMParityStatus;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnBypass HwtLpCsEnBypass;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMNopAddr ACSMNopAddr;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_SnoopCntrl SnoopCntrl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityInvert ACSMParityInvert;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmPsIndx AcsmPsIndx;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmDynPtrCtrl AcsmDynPtrCtrl;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_FspState FspState;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable0 AcsmMapTable0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable1 AcsmMapTable1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable2 AcsmMapTable2;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable3 AcsmMapTable3;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable4 AcsmMapTable4;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable5 AcsmMapTable5;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable6 AcsmMapTable6;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable7 AcsmMapTable7;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable8 AcsmMapTable8;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable9 AcsmMapTable9;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable10 AcsmMapTable10;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable11 AcsmMapTable11;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable12 AcsmMapTable12;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable13 AcsmMapTable13;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable14 AcsmMapTable14;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable15 AcsmMapTable15;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable16 AcsmMapTable16;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable17 AcsmMapTable17;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable18 AcsmMapTable18;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable19 AcsmMapTable19;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable20 AcsmMapTable20;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable21 AcsmMapTable21;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable22 AcsmMapTable22;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable23 AcsmMapTable23;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable24 AcsmMapTable24;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable25 AcsmMapTable25;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable26 AcsmMapTable26;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable27 AcsmMapTable27;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable28 AcsmMapTable28;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable29 AcsmMapTable29;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable30 AcsmMapTable30;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable31 AcsmMapTable31;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable32 AcsmMapTable32;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable33 AcsmMapTable33;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable34 AcsmMapTable34;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable35 AcsmMapTable35;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable36 AcsmMapTable36;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable37 AcsmMapTable37;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable38 AcsmMapTable38;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable39 AcsmMapTable39;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable40 AcsmMapTable40;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable41 AcsmMapTable41;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable42 AcsmMapTable42;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable43 AcsmMapTable43;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable44 AcsmMapTable44;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable45 AcsmMapTable45;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable46 AcsmMapTable46;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable47 AcsmMapTable47;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable48 AcsmMapTable48;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable49 AcsmMapTable49;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable50 AcsmMapTable50;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable51 AcsmMapTable51;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable52 AcsmMapTable52;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable53 AcsmMapTable53;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable54 AcsmMapTable54;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable55 AcsmMapTable55;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable56 AcsmMapTable56;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable57 AcsmMapTable57;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable58 AcsmMapTable58;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable59 AcsmMapTable59;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable60 AcsmMapTable60;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable61 AcsmMapTable61;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable62 AcsmMapTable62;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable63 AcsmMapTable63;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal0 AcsmStartAddrXlatVal0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal1 AcsmStartAddrXlatVal1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal2 AcsmStartAddrXlatVal2;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal3 AcsmStartAddrXlatVal3;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal4 AcsmStartAddrXlatVal4;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal5 AcsmStartAddrXlatVal5;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal6 AcsmStartAddrXlatVal6;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal7 AcsmStartAddrXlatVal7;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal8 AcsmStartAddrXlatVal8;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal9 AcsmStartAddrXlatVal9;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal10 AcsmStartAddrXlatVal10;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal11 AcsmStartAddrXlatVal11;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal12 AcsmStartAddrXlatVal12;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal13 AcsmStartAddrXlatVal13;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal14 AcsmStartAddrXlatVal14;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal15 AcsmStartAddrXlatVal15;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal16 AcsmStartAddrXlatVal16;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal17 AcsmStartAddrXlatVal17;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal18 AcsmStartAddrXlatVal18;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal19 AcsmStartAddrXlatVal19;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal20 AcsmStartAddrXlatVal20;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal21 AcsmStartAddrXlatVal21;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal22 AcsmStartAddrXlatVal22;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal23 AcsmStartAddrXlatVal23;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal24 AcsmStartAddrXlatVal24;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal25 AcsmStartAddrXlatVal25;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal26 AcsmStartAddrXlatVal26;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal27 AcsmStartAddrXlatVal27;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal28 AcsmStartAddrXlatVal28;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal29 AcsmStartAddrXlatVal29;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal30 AcsmStartAddrXlatVal30;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal31 AcsmStartAddrXlatVal31;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal32 AcsmStartAddrXlatVal32;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal33 AcsmStartAddrXlatVal33;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal34 AcsmStartAddrXlatVal34;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal35 AcsmStartAddrXlatVal35;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal36 AcsmStartAddrXlatVal36;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal37 AcsmStartAddrXlatVal37;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal38 AcsmStartAddrXlatVal38;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal39 AcsmStartAddrXlatVal39;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal40 AcsmStartAddrXlatVal40;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal41 AcsmStartAddrXlatVal41;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal42 AcsmStartAddrXlatVal42;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal43 AcsmStartAddrXlatVal43;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal44 AcsmStartAddrXlatVal44;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal45 AcsmStartAddrXlatVal45;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal46 AcsmStartAddrXlatVal46;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal47 AcsmStartAddrXlatVal47;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal48 AcsmStartAddrXlatVal48;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal49 AcsmStartAddrXlatVal49;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal50 AcsmStartAddrXlatVal50;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal51 AcsmStartAddrXlatVal51;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal52 AcsmStartAddrXlatVal52;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal53 AcsmStartAddrXlatVal53;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal54 AcsmStartAddrXlatVal54;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal55 AcsmStartAddrXlatVal55;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal56 AcsmStartAddrXlatVal56;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal57 AcsmStartAddrXlatVal57;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal58 AcsmStartAddrXlatVal58;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal59 AcsmStartAddrXlatVal59;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal60 AcsmStartAddrXlatVal60;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal61 AcsmStartAddrXlatVal61;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal62 AcsmStartAddrXlatVal62;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal63 AcsmStartAddrXlatVal63;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal0 AcsmStopAddrXlatVal0;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal1 AcsmStopAddrXlatVal1;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal2 AcsmStopAddrXlatVal2;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal3 AcsmStopAddrXlatVal3;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal4 AcsmStopAddrXlatVal4;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal5 AcsmStopAddrXlatVal5;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal6 AcsmStopAddrXlatVal6;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal7 AcsmStopAddrXlatVal7;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal8 AcsmStopAddrXlatVal8;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal9 AcsmStopAddrXlatVal9;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal10 AcsmStopAddrXlatVal10;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal11 AcsmStopAddrXlatVal11;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal12 AcsmStopAddrXlatVal12;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal13 AcsmStopAddrXlatVal13;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal14 AcsmStopAddrXlatVal14;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal15 AcsmStopAddrXlatVal15;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal16 AcsmStopAddrXlatVal16;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal17 AcsmStopAddrXlatVal17;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal18 AcsmStopAddrXlatVal18;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal19 AcsmStopAddrXlatVal19;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal20 AcsmStopAddrXlatVal20;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal21 AcsmStopAddrXlatVal21;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal22 AcsmStopAddrXlatVal22;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal23 AcsmStopAddrXlatVal23;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal24 AcsmStopAddrXlatVal24;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal25 AcsmStopAddrXlatVal25;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal26 AcsmStopAddrXlatVal26;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal27 AcsmStopAddrXlatVal27;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal28 AcsmStopAddrXlatVal28;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal29 AcsmStopAddrXlatVal29;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal30 AcsmStopAddrXlatVal30;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal31 AcsmStopAddrXlatVal31;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal32 AcsmStopAddrXlatVal32;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal33 AcsmStopAddrXlatVal33;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal34 AcsmStopAddrXlatVal34;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal35 AcsmStopAddrXlatVal35;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal36 AcsmStopAddrXlatVal36;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal37 AcsmStopAddrXlatVal37;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal38 AcsmStopAddrXlatVal38;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal39 AcsmStopAddrXlatVal39;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal40 AcsmStopAddrXlatVal40;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal41 AcsmStopAddrXlatVal41;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal42 AcsmStopAddrXlatVal42;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal43 AcsmStopAddrXlatVal43;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal44 AcsmStopAddrXlatVal44;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal45 AcsmStopAddrXlatVal45;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal46 AcsmStopAddrXlatVal46;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal47 AcsmStopAddrXlatVal47;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal48 AcsmStopAddrXlatVal48;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal49 AcsmStopAddrXlatVal49;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal50 AcsmStopAddrXlatVal50;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal51 AcsmStopAddrXlatVal51;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal52 AcsmStopAddrXlatVal52;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal53 AcsmStopAddrXlatVal53;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal54 AcsmStopAddrXlatVal54;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal55 AcsmStopAddrXlatVal55;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal56 AcsmStopAddrXlatVal56;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal57 AcsmStopAddrXlatVal57;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal58 AcsmStopAddrXlatVal58;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal59 AcsmStopAddrXlatVal59;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal60 AcsmStopAddrXlatVal60;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal61 AcsmStopAddrXlatVal61;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal62 AcsmStopAddrXlatVal62;
	rand ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal63 AcsmStopAddrXlatVal63;
   local uvm_reg_data_t m_offset;
	rand uvm_reg_field PpgcGenCtrl_PpgcGenCtrl;
	rand uvm_reg_field PpgcGenDbiCtrl_PpgcGenDbiCtrl;
	rand uvm_reg_field PpgcGenDbiConfig_PpgcGenDbiConfig;
	rand uvm_reg_field PpgcGenLaneMuxSel0_PpgcGenLaneMuxSel0;
	rand uvm_reg_field PpgcGenLaneMuxSel1_PpgcGenLaneMuxSel1;
	rand uvm_reg_field EnPhyUpdZQCalUpdate_EnPhyUpdZQCalUpdate;
	rand uvm_reg_field BlockDfiInterface_BlockDfiInterfaceEn;
	rand uvm_reg_field BlockDfiInterfaceEn;
	rand uvm_reg_field BlockDfiInterface_BlockDfiInterfaceStatusReset;
	rand uvm_reg_field BlockDfiInterfaceStatusReset;
	rand uvm_reg_field BlockDfiInterface_PmuBusy;
	rand uvm_reg_field PmuBusy;
	uvm_reg_field BlockDfiInterfaceStatus_BlockDfiInterfaceStatus;
	rand uvm_reg_field DfiCustMode_p0_DfiCustMode_p0;
	rand uvm_reg_field HwtMRL_p0_HwtMRL_p0;
	rand uvm_reg_field RegRet_RegRet;
	rand uvm_reg_field DisableZQupdateOnSnoop_DisableZQupdateOnSnoop;
	rand uvm_reg_field Prbs0GenModeSel_Prbs0GenModeSel;
	rand uvm_reg_field Prbs0GenUiMuxSel_Prbs0GenUiMuxSel;
	rand uvm_reg_field Prbs0GenTapDly0_Prbs0GenTapDly0;
	rand uvm_reg_field Prbs0GenTapDly1_Prbs0GenTapDly1;
	rand uvm_reg_field Prbs0GenTapDly2_Prbs0GenTapDly2;
	rand uvm_reg_field Prbs0GenTapDly3_Prbs0GenTapDly3;
	rand uvm_reg_field Prbs0GenTapDly4_Prbs0GenTapDly4;
	rand uvm_reg_field Prbs0GenTapDly5_Prbs0GenTapDly5;
	rand uvm_reg_field Prbs0GenTapDly6_Prbs0GenTapDly6;
	rand uvm_reg_field Prbs0GenTapDly7_Prbs0GenTapDly7;
	rand uvm_reg_field MtestMuxSel_MtestMuxSel;
	rand uvm_reg_field Prbs0GenStateLo_Prbs0GenStateLo;
	rand uvm_reg_field Prbs0GenStateHi_Prbs0GenStateHi;
	rand uvm_reg_field Prbs1GenModeSel_Prbs1GenModeSel;
	rand uvm_reg_field Prbs1GenUiMuxSel_Prbs1GenUiMuxSel;
	rand uvm_reg_field Prbs1GenTapDly0_Prbs1GenTapDly0;
	rand uvm_reg_field Prbs1GenTapDly1_Prbs1GenTapDly1;
	rand uvm_reg_field Prbs1GenTapDly2_Prbs1GenTapDly2;
	rand uvm_reg_field Prbs1GenTapDly3_Prbs1GenTapDly3;
	rand uvm_reg_field Prbs1GenTapDly4_Prbs1GenTapDly4;
	rand uvm_reg_field Prbs1GenTapDly5_Prbs1GenTapDly5;
	rand uvm_reg_field Prbs1GenTapDly6_Prbs1GenTapDly6;
	rand uvm_reg_field Prbs1GenTapDly7_Prbs1GenTapDly7;
	rand uvm_reg_field Prbs1GenStateLo_Prbs1GenStateLo;
	rand uvm_reg_field Prbs1GenStateHi_Prbs1GenStateHi;
	rand uvm_reg_field Prbs2GenModeSel_Prbs2GenModeSel;
	rand uvm_reg_field Prbs2GenUiMuxSel_Prbs2GenUiMuxSel;
	rand uvm_reg_field Prbs2GenTapDly0_Prbs2GenTapDly0;
	rand uvm_reg_field Prbs2GenTapDly1_Prbs2GenTapDly1;
	rand uvm_reg_field Prbs2GenTapDly2_Prbs2GenTapDly2;
	rand uvm_reg_field Prbs2GenTapDly3_Prbs2GenTapDly3;
	rand uvm_reg_field Prbs2GenTapDly4_Prbs2GenTapDly4;
	rand uvm_reg_field Prbs2GenTapDly5_Prbs2GenTapDly5;
	rand uvm_reg_field Prbs2GenTapDly6_Prbs2GenTapDly6;
	rand uvm_reg_field Prbs2GenTapDly7_Prbs2GenTapDly7;
	rand uvm_reg_field Prbs2GenStateLo_Prbs2GenStateLo;
	rand uvm_reg_field Prbs2GenStateHi_Prbs2GenStateHi;
	rand uvm_reg_field PPTTrainSetup_p0_PhyMstrTrainInterval;
	rand uvm_reg_field PhyMstrTrainInterval;
	rand uvm_reg_field PPTTrainSetup_p0_PhyMstrMaxReqToAck;
	rand uvm_reg_field PhyMstrMaxReqToAck;
	rand uvm_reg_field PhyMstrFreqOverride_p0_PhyMstrFreqOverride_p0;
	rand uvm_reg_field DfiInitComplete_DfiInitComplete;
	rand uvm_reg_field PPGCParityInvert_PPGCParityInvert;
	rand uvm_reg_field PMIEnable_PMIEnable;
	uvm_reg_field Dfi0Status_Dfi0Status;
	uvm_reg_field Dfi1Status_Dfi1Status;
	rand uvm_reg_field DfiHandshakeDelays0_p0_PhyUpdAckDelay0;
	rand uvm_reg_field PhyUpdAckDelay0;
	rand uvm_reg_field DfiHandshakeDelays0_p0_PhyUpdReqDelay0;
	rand uvm_reg_field PhyUpdReqDelay0;
	rand uvm_reg_field DfiHandshakeDelays0_p0_CtrlUpdReqDelay0;
	rand uvm_reg_field CtrlUpdReqDelay0;
	rand uvm_reg_field DFIPHYUPD0_DFIPHYUPDCNT0;
	rand uvm_reg_field DFIPHYUPDCNT0;
	rand uvm_reg_field DFIPHYUPD0_DFIPHYUPDRESP0;
	rand uvm_reg_field DFIPHYUPDRESP0;
	rand uvm_reg_field DfiLpCtrlEn0_DfiLpCtrlEn0;
	rand uvm_reg_field DfiLpDataEn0_DfiLpDataEn0;
	rand uvm_reg_field DynOdtEnCntrl0_DbyteDynOdtEn0;
	rand uvm_reg_field DbyteDynOdtEn0;
	rand uvm_reg_field DfiRespHandshakeDelays0_p0_LpCtrlAckDelay0;
	rand uvm_reg_field LpCtrlAckDelay0;
	rand uvm_reg_field DfiRespHandshakeDelays0_p0_LpDataAckDelay0;
	rand uvm_reg_field LpDataAckDelay0;
	rand uvm_reg_field DfiRespHandshakeDelays0_p0_CtrlUpdAckDelay0;
	rand uvm_reg_field CtrlUpdAckDelay0;
	rand uvm_reg_field DfiRespHandshakeDelays0_p0_LpAssertAckDelay0;
	rand uvm_reg_field LpAssertAckDelay0;
	rand uvm_reg_field HwtLpCsEnA_HwtLpCsEnA;
	rand uvm_reg_field HwtLpCsEnB_HwtLpCsEnB;
	rand uvm_reg_field HwtCtrl_HwtCtrl;
	rand uvm_reg_field HwtControlOvr_HwtControlOvr;
	rand uvm_reg_field ScratchPadPPGC_ScratchPadPPGC;
	rand uvm_reg_field HwtControlVal_HwtControlVal;
	rand uvm_reg_field ForceHWTClkGaterEnables_ForceACSMClkEnHigh;
	rand uvm_reg_field ForceACSMClkEnHigh;
	rand uvm_reg_field ForceHWTClkGaterEnables_ForceACSMClkEnLow;
	rand uvm_reg_field ForceACSMClkEnLow;
	rand uvm_reg_field ForceHWTClkGaterEnables_ForcePIEClkEnHigh;
	rand uvm_reg_field ForcePIEClkEnHigh;
	rand uvm_reg_field ForceHWTClkGaterEnables_ForcePIEClkEnLow;
	rand uvm_reg_field ForcePIEClkEnLow;
	uvm_reg_field MasUpdGoodCtr_MasUpdGoodCtr;
	uvm_reg_field PhyUpd0GoodCtr_PhyUpd0GoodCtr;
	uvm_reg_field PhyUpd1GoodCtr_PhyUpd1GoodCtr;
	uvm_reg_field CtlUpd0GoodCtr_CtlUpd0GoodCtr;
	uvm_reg_field CtlUpd1GoodCtr_CtlUpd1GoodCtr;
	uvm_reg_field MasUpdFailCtr_MasUpdFailCtr;
	uvm_reg_field PhyUpd0FailCtr_PhyUpd0FailCtr;
	uvm_reg_field PhyUpd1FailCtr_PhyUpd1FailCtr;
	rand uvm_reg_field PhyPerfCtrEnable_MasUpdGoodCtl;
	rand uvm_reg_field MasUpdGoodCtl;
	rand uvm_reg_field PhyPerfCtrEnable_PhyUpd0GoodCtl;
	rand uvm_reg_field PhyUpd0GoodCtl;
	rand uvm_reg_field PhyPerfCtrEnable_PhyUpd1GoodCtl;
	rand uvm_reg_field PhyUpd1GoodCtl;
	rand uvm_reg_field PhyPerfCtrEnable_CtlUpd0GoodCtl;
	rand uvm_reg_field CtlUpd0GoodCtl;
	rand uvm_reg_field PhyPerfCtrEnable_CtlUpd1GoodCtl;
	rand uvm_reg_field CtlUpd1GoodCtl;
	rand uvm_reg_field PhyPerfCtrEnable_MasUpdFailCtl;
	rand uvm_reg_field MasUpdFailCtl;
	rand uvm_reg_field PhyPerfCtrEnable_PhyUpd0FailCtl;
	rand uvm_reg_field PhyUpd0FailCtl;
	rand uvm_reg_field PhyPerfCtrEnable_PhyUpd1FailCtl;
	rand uvm_reg_field PhyUpd1FailCtl;
	rand uvm_reg_field DfiHandshakeDelays1_p0_PhyUpdAckDelay1;
	rand uvm_reg_field PhyUpdAckDelay1;
	rand uvm_reg_field DfiHandshakeDelays1_p0_PhyUpdReqDelay1;
	rand uvm_reg_field PhyUpdReqDelay1;
	rand uvm_reg_field DfiHandshakeDelays1_p0_CtrlUpdReqDelay1;
	rand uvm_reg_field CtrlUpdReqDelay1;
	rand uvm_reg_field DFIPHYUPD1_DFIPHYUPDCNT1;
	rand uvm_reg_field DFIPHYUPDCNT1;
	rand uvm_reg_field DFIPHYUPD1_DFIPHYUPDRESP1;
	rand uvm_reg_field DFIPHYUPDRESP1;
	rand uvm_reg_field DfiLpCtrlEn1_DfiLpCtrlEn1;
	rand uvm_reg_field DfiLpDataEn1_DfiLpDataEn1;
	rand uvm_reg_field DynOdtEnCntrl1_DbyteDynOdtEn1;
	rand uvm_reg_field DbyteDynOdtEn1;
	rand uvm_reg_field DfiRespHandshakeDelays1_p0_LpCtrlAckDelay1;
	rand uvm_reg_field LpCtrlAckDelay1;
	rand uvm_reg_field DfiRespHandshakeDelays1_p0_LpDataAckDelay1;
	rand uvm_reg_field LpDataAckDelay1;
	rand uvm_reg_field DfiRespHandshakeDelays1_p0_CtrlUpdAckDelay1;
	rand uvm_reg_field CtrlUpdAckDelay1;
	rand uvm_reg_field DfiRespHandshakeDelays1_p0_LpAssertAckDelay1;
	rand uvm_reg_field LpAssertAckDelay1;
	rand uvm_reg_field FspSkipList_FspPStateSkip0;
	rand uvm_reg_field FspPStateSkip0;
	rand uvm_reg_field FspSkipList_FspPStateSkip1;
	rand uvm_reg_field FspPStateSkip1;
	rand uvm_reg_field FspSkipList_FspPStateSkip2;
	rand uvm_reg_field FspPStateSkip2;
	rand uvm_reg_field FspSkipList_FspPStateSkip3;
	rand uvm_reg_field FspPStateSkip3;
	rand uvm_reg_field PPGCReserved0_PPGCReserved0;
	rand uvm_reg_field PUBReservedP1_p0_PUBReservedP1_p0;
	rand uvm_reg_field PhyInterruptOverride_PhyInterruptOverride;
	rand uvm_reg_field PhyInterruptEnable_PhyTrngCmpltEn;
	rand uvm_reg_field PhyTrngCmpltEn;
	rand uvm_reg_field PhyInterruptEnable_PhyInitCmpltEn;
	rand uvm_reg_field PhyInitCmpltEn;
	rand uvm_reg_field PhyInterruptEnable_PhyTrngFailEn;
	rand uvm_reg_field PhyTrngFailEn;
	rand uvm_reg_field PhyInterruptEnable_PhyFWReservedEn;
	rand uvm_reg_field PhyFWReservedEn;
	rand uvm_reg_field PhyInterruptEnable_PhyAcsmParityErrEn;
	rand uvm_reg_field PhyAcsmParityErrEn;
	rand uvm_reg_field PhyInterruptEnable_PhyPIEParityErrEn;
	rand uvm_reg_field PhyPIEParityErrEn;
	rand uvm_reg_field PhyInterruptEnable_PhyRdfPtrChkErrEn;
	rand uvm_reg_field PhyRdfPtrChkErrEn;
	rand uvm_reg_field PhyInterruptEnable_PhyEccEn;
	rand uvm_reg_field PhyEccEn;
	rand uvm_reg_field PhyInterruptEnable_PhyPIEProgErrEn;
	rand uvm_reg_field PhyPIEProgErrEn;
	rand uvm_reg_field PhyInterruptEnable_PhyHWReservedEn;
	rand uvm_reg_field PhyHWReservedEn;
	rand uvm_reg_field PhyInterruptFWControl_PhyTrngCmpltFW;
	rand uvm_reg_field PhyTrngCmpltFW;
	rand uvm_reg_field PhyInterruptFWControl_PhyInitCmpltFW;
	rand uvm_reg_field PhyInitCmpltFW;
	rand uvm_reg_field PhyInterruptFWControl_PhyTrngFailFW;
	rand uvm_reg_field PhyTrngFailFW;
	rand uvm_reg_field PhyInterruptFWControl_PhyFWReservedFW;
	rand uvm_reg_field PhyFWReservedFW;
	rand uvm_reg_field PhyInterruptMask_PhyTrngCmpltMsk;
	rand uvm_reg_field PhyTrngCmpltMsk;
	rand uvm_reg_field PhyInterruptMask_PhyInitCmpltMsk;
	rand uvm_reg_field PhyInitCmpltMsk;
	rand uvm_reg_field PhyInterruptMask_PhyTrngFailMsk;
	rand uvm_reg_field PhyTrngFailMsk;
	rand uvm_reg_field PhyInterruptMask_PhyFWReservedMsk;
	rand uvm_reg_field PhyFWReservedMsk;
	rand uvm_reg_field PhyInterruptMask_PhyAcsmParityErrMsk;
	rand uvm_reg_field PhyAcsmParityErrMsk;
	rand uvm_reg_field PhyInterruptMask_PhyPIEParityErrMsk;
	rand uvm_reg_field PhyPIEParityErrMsk;
	rand uvm_reg_field PhyInterruptMask_PhyRdfPtrChkErrMsk;
	rand uvm_reg_field PhyRdfPtrChkErrMsk;
	rand uvm_reg_field PhyInterruptMask_PhyEccMsk;
	rand uvm_reg_field PhyEccMsk;
	rand uvm_reg_field PhyInterruptMask_PhyPIEProgErrMsk;
	rand uvm_reg_field PhyPIEProgErrMsk;
	rand uvm_reg_field PhyInterruptMask_PhyHWReservedMsk;
	rand uvm_reg_field PhyHWReservedMsk;
	rand uvm_reg_field PhyInterruptClear_PhyTrngCmpltClr;
	rand uvm_reg_field PhyTrngCmpltClr;
	rand uvm_reg_field PhyInterruptClear_PhyInitCmpltClr;
	rand uvm_reg_field PhyInitCmpltClr;
	rand uvm_reg_field PhyInterruptClear_PhyTrngFailClr;
	rand uvm_reg_field PhyTrngFailClr;
	rand uvm_reg_field PhyInterruptClear_PhyFWReservedClr;
	rand uvm_reg_field PhyFWReservedClr;
	rand uvm_reg_field PhyInterruptClear_PhyAcsmParityErrClr;
	rand uvm_reg_field PhyAcsmParityErrClr;
	rand uvm_reg_field PhyInterruptClear_PhyPIEParityErrClr;
	rand uvm_reg_field PhyPIEParityErrClr;
	rand uvm_reg_field PhyInterruptClear_PhyRdfPtrChkErrClr;
	rand uvm_reg_field PhyRdfPtrChkErrClr;
	rand uvm_reg_field PhyInterruptClear_PhyEccClr;
	rand uvm_reg_field PhyEccClr;
	rand uvm_reg_field PhyInterruptClear_PhyPIEProgErrClr;
	rand uvm_reg_field PhyPIEProgErrClr;
	rand uvm_reg_field PhyInterruptClear_PhyHWReservedClr;
	rand uvm_reg_field PhyHWReservedClr;
	uvm_reg_field PhyInterruptStatus_PhyTrngCmplt;
	uvm_reg_field PhyTrngCmplt;
	uvm_reg_field PhyInterruptStatus_PhyInitCmplt;
	uvm_reg_field PhyInitCmplt;
	uvm_reg_field PhyInterruptStatus_PhyTrngFail;
	uvm_reg_field PhyTrngFail;
	uvm_reg_field PhyInterruptStatus_PhyFWReserved;
	uvm_reg_field PhyFWReserved;
	uvm_reg_field PhyInterruptStatus_PhyAcsmParityErr;
	uvm_reg_field PhyAcsmParityErr;
	uvm_reg_field PhyInterruptStatus_PhyPIEParityErr;
	uvm_reg_field PhyPIEParityErr;
	uvm_reg_field PhyInterruptStatus_PhyRdfPtrChkErr;
	uvm_reg_field PhyRdfPtrChkErr;
	uvm_reg_field PhyInterruptStatus_PhyEccErr;
	uvm_reg_field PhyEccErr;
	uvm_reg_field PhyInterruptStatus_PhyPIEProgErr;
	uvm_reg_field PhyPIEProgErr;
	uvm_reg_field PhyInterruptStatus_PhyHWReserved;
	uvm_reg_field PhyHWReserved;
	rand uvm_reg_field ACSMRunCtrl_ACSMRun;
	rand uvm_reg_field ACSMRun;
	rand uvm_reg_field ACSMRunCtrl_AcsmProgPtr;
	rand uvm_reg_field AcsmProgPtr;
	rand uvm_reg_field ACSMRunCtrl_ACSMXlatEn;
	rand uvm_reg_field ACSMXlatEn;
	rand uvm_reg_field ACSMRunCtrl_ACSMNopFlag;
	rand uvm_reg_field ACSMNopFlag;
	rand uvm_reg_field ACSMRunCtrl_ACSMRptCntOverrideEn;
	rand uvm_reg_field ACSMRptCntOverrideEn;
	uvm_reg_field ACSMDone_ACSMDone;
	rand uvm_reg_field ACSMStartAddr_p0_ACSMStartAddr_p0;
	rand uvm_reg_field ACSMStopAddr_p0_ACSMStopAddr_p0;
	uvm_reg_field ACSMLastAddr_ACSMLastAddr;
	rand uvm_reg_field ACSMAlgaIncVal_ACSMAlgaIncVal;
	rand uvm_reg_field ACSMAddressMask_ACSMAddressMask;
	rand uvm_reg_field ACSMOuterLoopRepeatCnt_ACSMOuterLoopRepeatCnt;
	rand uvm_reg_field ACSMCkeControl_ACSMCkeControl;
	uvm_reg_field ACSMCkeStatus_ACSMCkeStatus;
	rand uvm_reg_field ACSMWckEnControl_ACSMWckEnControl;
	uvm_reg_field ACSMWckEnStatus_ACSMWckEnStatus;
	rand uvm_reg_field ACSMRxEnPulse_p0_ACSMRxEnDelay;
	rand uvm_reg_field ACSMRxEnDelay;
	rand uvm_reg_field ACSMRxEnPulse_p0_ACSMRxEnDelayReserved;
	rand uvm_reg_field ACSMRxEnDelayReserved;
	rand uvm_reg_field ACSMRxEnPulse_p0_ACSMRxEnWidth;
	rand uvm_reg_field ACSMRxEnWidth;
	rand uvm_reg_field ACSMRxValPulse_p0_ACSMRxValDelay;
	rand uvm_reg_field ACSMRxValDelay;
	rand uvm_reg_field ACSMRxValPulse_p0_ACSMRxValDelayReserved;
	rand uvm_reg_field ACSMRxValDelayReserved;
	rand uvm_reg_field ACSMRxValPulse_p0_ACSMRxValWidth;
	rand uvm_reg_field ACSMRxValWidth;
	rand uvm_reg_field ACSMTxEnPulse_p0_ACSMTxEnDelay;
	rand uvm_reg_field ACSMTxEnDelay;
	rand uvm_reg_field ACSMTxEnPulse_p0_ACSMTxEnDelayReserved;
	rand uvm_reg_field ACSMTxEnDelayReserved;
	rand uvm_reg_field ACSMTxEnPulse_p0_ACSMTxEnWidth;
	rand uvm_reg_field ACSMTxEnWidth;
	rand uvm_reg_field ACSMWrcsPulse_p0_ACSMWrcsDelay;
	rand uvm_reg_field ACSMWrcsDelay;
	rand uvm_reg_field ACSMWrcsPulse_p0_ACSMWrcsDelayReserved;
	rand uvm_reg_field ACSMWrcsDelayReserved;
	rand uvm_reg_field ACSMWrcsPulse_p0_ACSMWrcsWidth;
	rand uvm_reg_field ACSMWrcsWidth;
	rand uvm_reg_field ACSMRdcsPulse_p0_ACSMRdcsDelay;
	rand uvm_reg_field ACSMRdcsDelay;
	rand uvm_reg_field ACSMRdcsPulse_p0_ACSMRdcsDelayReserved;
	rand uvm_reg_field ACSMRdcsDelayReserved;
	rand uvm_reg_field ACSMRdcsPulse_p0_ACSMRdcsWidth;
	rand uvm_reg_field ACSMRdcsWidth;
	rand uvm_reg_field ACSMInfiniteOLRC_ACSMInfiniteOLRC;
	rand uvm_reg_field ACSMDefaultAddr_ACSMDefaultAddr;
	rand uvm_reg_field ACSMDefaultCs_ACSMDefaultCs;
	rand uvm_reg_field ACSMStaticCtrl_ACSMPhaseControl;
	rand uvm_reg_field ACSMPhaseControl;
	rand uvm_reg_field ACSMWckWriteStaticLoPulse_p0_ACSMWckWriteStaticLoDelay;
	rand uvm_reg_field ACSMWckWriteStaticLoDelay;
	rand uvm_reg_field ACSMWckWriteStaticLoPulse_p0_ACSMWckWriteStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckWriteStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckWriteStaticLoPulse_p0_ACSMWckWriteStaticLoWidth;
	rand uvm_reg_field ACSMWckWriteStaticLoWidth;
	rand uvm_reg_field ACSMWckWriteStaticHiPulse_p0_ACSMWckWriteStaticHiDelay;
	rand uvm_reg_field ACSMWckWriteStaticHiDelay;
	rand uvm_reg_field ACSMWckWriteStaticHiPulse_p0_ACSMWckWriteStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckWriteStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckWriteStaticHiPulse_p0_ACSMWckWriteStaticHiWidth;
	rand uvm_reg_field ACSMWckWriteStaticHiWidth;
	rand uvm_reg_field ACSMWckWriteTogglePulse_p0_ACSMWckWriteToggleDelay;
	rand uvm_reg_field ACSMWckWriteToggleDelay;
	rand uvm_reg_field ACSMWckWriteTogglePulse_p0_ACSMWckWriteToggleDelayReserved;
	rand uvm_reg_field ACSMWckWriteToggleDelayReserved;
	rand uvm_reg_field ACSMWckWriteTogglePulse_p0_ACSMWckWriteToggleWidth;
	rand uvm_reg_field ACSMWckWriteToggleWidth;
	rand uvm_reg_field ACSMWckWriteFastTogglePulse_p0_ACSMWckWriteFastToggleDelay;
	rand uvm_reg_field ACSMWckWriteFastToggleDelay;
	rand uvm_reg_field ACSMWckWriteFastTogglePulse_p0_ACSMWckWriteFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckWriteFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckWriteFastTogglePulse_p0_ACSMWckWriteFastToggleWidth;
	rand uvm_reg_field ACSMWckWriteFastToggleWidth;
	rand uvm_reg_field ACSMWckReadStaticLoPulse_p0_ACSMWckReadStaticLoDelay;
	rand uvm_reg_field ACSMWckReadStaticLoDelay;
	rand uvm_reg_field ACSMWckReadStaticLoPulse_p0_ACSMWckReadStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckReadStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckReadStaticLoPulse_p0_ACSMWckReadStaticLoWidth;
	rand uvm_reg_field ACSMWckReadStaticLoWidth;
	rand uvm_reg_field ACSMWckReadStaticHiPulse_p0_ACSMWckReadStaticHiDelay;
	rand uvm_reg_field ACSMWckReadStaticHiDelay;
	rand uvm_reg_field ACSMWckReadStaticHiPulse_p0_ACSMWckReadStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckReadStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckReadStaticHiPulse_p0_ACSMWckReadStaticHiWidth;
	rand uvm_reg_field ACSMWckReadStaticHiWidth;
	rand uvm_reg_field ACSMWckReadTogglePulse_p0_ACSMWckReadToggleDelay;
	rand uvm_reg_field ACSMWckReadToggleDelay;
	rand uvm_reg_field ACSMWckReadTogglePulse_p0_ACSMWckReadToggleDelayReserved;
	rand uvm_reg_field ACSMWckReadToggleDelayReserved;
	rand uvm_reg_field ACSMWckReadTogglePulse_p0_ACSMWckReadToggleWidth;
	rand uvm_reg_field ACSMWckReadToggleWidth;
	rand uvm_reg_field ACSMWckReadFastTogglePulse_p0_ACSMWckReadFastToggleDelay;
	rand uvm_reg_field ACSMWckReadFastToggleDelay;
	rand uvm_reg_field ACSMWckReadFastTogglePulse_p0_ACSMWckReadFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckReadFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckReadFastTogglePulse_p0_ACSMWckReadFastToggleWidth;
	rand uvm_reg_field ACSMWckReadFastToggleWidth;
	rand uvm_reg_field ACSMWckFreqSwStaticLoPulse_p0_ACSMWckFreqSwStaticLoDelay;
	rand uvm_reg_field ACSMWckFreqSwStaticLoDelay;
	rand uvm_reg_field ACSMWckFreqSwStaticLoPulse_p0_ACSMWckFreqSwStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwStaticLoDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwStaticLoPulse_p0_ACSMWckFreqSwStaticLoWidth;
	rand uvm_reg_field ACSMWckFreqSwStaticLoWidth;
	rand uvm_reg_field ACSMWckFreqSwStaticHiPulse_p0_ACSMWckFreqSwStaticHiDelay;
	rand uvm_reg_field ACSMWckFreqSwStaticHiDelay;
	rand uvm_reg_field ACSMWckFreqSwStaticHiPulse_p0_ACSMWckFreqSwStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwStaticHiDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwStaticHiPulse_p0_ACSMWckFreqSwStaticHiWidth;
	rand uvm_reg_field ACSMWckFreqSwStaticHiWidth;
	rand uvm_reg_field ACSMWckFreqSwTogglePulse_p0_ACSMWckFreqSwToggleDelay;
	rand uvm_reg_field ACSMWckFreqSwToggleDelay;
	rand uvm_reg_field ACSMWckFreqSwTogglePulse_p0_ACSMWckFreqSwToggleDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwToggleDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwTogglePulse_p0_ACSMWckFreqSwToggleWidth;
	rand uvm_reg_field ACSMWckFreqSwToggleWidth;
	rand uvm_reg_field ACSMWckFreqSwFastTogglePulse_p0_ACSMWckFreqSwFastToggleDelay;
	rand uvm_reg_field ACSMWckFreqSwFastToggleDelay;
	rand uvm_reg_field ACSMWckFreqSwFastTogglePulse_p0_ACSMWckFreqSwFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwFastToggleDelayReserved;
	rand uvm_reg_field ACSMWckFreqSwFastTogglePulse_p0_ACSMWckFreqSwFastToggleWidth;
	rand uvm_reg_field ACSMWckFreqSwFastToggleWidth;
	rand uvm_reg_field ACSMWckFreeRunMode_p0_ACSMWckFreeRunMode_p0;
	rand uvm_reg_field ACSMLowSpeedClockEnable_ACSMLowSpeedClockEnable;
	rand uvm_reg_field ACSMLowSpeedClockDelay_ACSMLowSpeedClockDelay;
	rand uvm_reg_field ACSMRptCntOverride_p0_ACSMRptCntOverride_p0;
	rand uvm_reg_field ACSMRptCntDbl_p0_ACSMRptCntDbl_p0;
	uvm_reg_field ACSMParityStatus_ACSMParityStatus;
	rand uvm_reg_field HwtLpCsEnBypass_HwtLpCsEnBypass;
	rand uvm_reg_field ACSMNopAddr_ACSMNopAddr;
	rand uvm_reg_field SnoopCntrl_SnoopCntrl;
	rand uvm_reg_field ACSMParityInvert_ACSMParityInvert;
	rand uvm_reg_field AcsmPsIndx_AcsmPsIndx;
	rand uvm_reg_field AcsmDynPtrCtrl_AcsmDynPtrCtrl;
	rand uvm_reg_field FspState_DramFsp0xPhyPs;
	rand uvm_reg_field DramFsp0xPhyPs;
	rand uvm_reg_field FspState_DramFsp1xPhyPs;
	rand uvm_reg_field DramFsp1xPhyPs;
	rand uvm_reg_field FspState_DramFsp2xPhyPs;
	rand uvm_reg_field DramFsp2xPhyPs;
	rand uvm_reg_field AcsmMapTable0_AcsmMapTableVal0;
	rand uvm_reg_field AcsmMapTableVal0;
	rand uvm_reg_field AcsmMapTable0_AcsmMapTableVal1;
	rand uvm_reg_field AcsmMapTableVal1;
	rand uvm_reg_field AcsmMapTable1_AcsmMapTableVal2;
	rand uvm_reg_field AcsmMapTableVal2;
	rand uvm_reg_field AcsmMapTable1_AcsmMapTableVal3;
	rand uvm_reg_field AcsmMapTableVal3;
	rand uvm_reg_field AcsmMapTable2_AcsmMapTableVal4;
	rand uvm_reg_field AcsmMapTableVal4;
	rand uvm_reg_field AcsmMapTable2_AcsmMapTableVal5;
	rand uvm_reg_field AcsmMapTableVal5;
	rand uvm_reg_field AcsmMapTable3_AcsmMapTableVal6;
	rand uvm_reg_field AcsmMapTableVal6;
	rand uvm_reg_field AcsmMapTable3_AcsmMapTableVal7;
	rand uvm_reg_field AcsmMapTableVal7;
	rand uvm_reg_field AcsmMapTable4_AcsmMapTableVal8;
	rand uvm_reg_field AcsmMapTableVal8;
	rand uvm_reg_field AcsmMapTable4_AcsmMapTableVal9;
	rand uvm_reg_field AcsmMapTableVal9;
	rand uvm_reg_field AcsmMapTable5_AcsmMapTableVal10;
	rand uvm_reg_field AcsmMapTableVal10;
	rand uvm_reg_field AcsmMapTable5_AcsmMapTableVal11;
	rand uvm_reg_field AcsmMapTableVal11;
	rand uvm_reg_field AcsmMapTable6_AcsmMapTableVal12;
	rand uvm_reg_field AcsmMapTableVal12;
	rand uvm_reg_field AcsmMapTable6_AcsmMapTableVal13;
	rand uvm_reg_field AcsmMapTableVal13;
	rand uvm_reg_field AcsmMapTable7_AcsmMapTableVal14;
	rand uvm_reg_field AcsmMapTableVal14;
	rand uvm_reg_field AcsmMapTable7_AcsmMapTableVal15;
	rand uvm_reg_field AcsmMapTableVal15;
	rand uvm_reg_field AcsmMapTable8_AcsmMapTableVal16;
	rand uvm_reg_field AcsmMapTableVal16;
	rand uvm_reg_field AcsmMapTable8_AcsmMapTableVal17;
	rand uvm_reg_field AcsmMapTableVal17;
	rand uvm_reg_field AcsmMapTable9_AcsmMapTableVal18;
	rand uvm_reg_field AcsmMapTableVal18;
	rand uvm_reg_field AcsmMapTable9_AcsmMapTableVal19;
	rand uvm_reg_field AcsmMapTableVal19;
	rand uvm_reg_field AcsmMapTable10_AcsmMapTableVal20;
	rand uvm_reg_field AcsmMapTableVal20;
	rand uvm_reg_field AcsmMapTable10_AcsmMapTableVal21;
	rand uvm_reg_field AcsmMapTableVal21;
	rand uvm_reg_field AcsmMapTable11_AcsmMapTableVal22;
	rand uvm_reg_field AcsmMapTableVal22;
	rand uvm_reg_field AcsmMapTable11_AcsmMapTableVal23;
	rand uvm_reg_field AcsmMapTableVal23;
	rand uvm_reg_field AcsmMapTable12_AcsmMapTableVal24;
	rand uvm_reg_field AcsmMapTableVal24;
	rand uvm_reg_field AcsmMapTable12_AcsmMapTableVal25;
	rand uvm_reg_field AcsmMapTableVal25;
	rand uvm_reg_field AcsmMapTable13_AcsmMapTableVal26;
	rand uvm_reg_field AcsmMapTableVal26;
	rand uvm_reg_field AcsmMapTable13_AcsmMapTableVal27;
	rand uvm_reg_field AcsmMapTableVal27;
	rand uvm_reg_field AcsmMapTable14_AcsmMapTableVal28;
	rand uvm_reg_field AcsmMapTableVal28;
	rand uvm_reg_field AcsmMapTable14_AcsmMapTableVal29;
	rand uvm_reg_field AcsmMapTableVal29;
	rand uvm_reg_field AcsmMapTable15_AcsmMapTableVal30;
	rand uvm_reg_field AcsmMapTableVal30;
	rand uvm_reg_field AcsmMapTable15_AcsmMapTableVal31;
	rand uvm_reg_field AcsmMapTableVal31;
	rand uvm_reg_field AcsmMapTable16_AcsmMapTableVal32;
	rand uvm_reg_field AcsmMapTableVal32;
	rand uvm_reg_field AcsmMapTable16_AcsmMapTableVal33;
	rand uvm_reg_field AcsmMapTableVal33;
	rand uvm_reg_field AcsmMapTable17_AcsmMapTableVal34;
	rand uvm_reg_field AcsmMapTableVal34;
	rand uvm_reg_field AcsmMapTable17_AcsmMapTableVal35;
	rand uvm_reg_field AcsmMapTableVal35;
	rand uvm_reg_field AcsmMapTable18_AcsmMapTableVal36;
	rand uvm_reg_field AcsmMapTableVal36;
	rand uvm_reg_field AcsmMapTable18_AcsmMapTableVal37;
	rand uvm_reg_field AcsmMapTableVal37;
	rand uvm_reg_field AcsmMapTable19_AcsmMapTableVal38;
	rand uvm_reg_field AcsmMapTableVal38;
	rand uvm_reg_field AcsmMapTable19_AcsmMapTableVal39;
	rand uvm_reg_field AcsmMapTableVal39;
	rand uvm_reg_field AcsmMapTable20_AcsmMapTableVal40;
	rand uvm_reg_field AcsmMapTableVal40;
	rand uvm_reg_field AcsmMapTable20_AcsmMapTableVal41;
	rand uvm_reg_field AcsmMapTableVal41;
	rand uvm_reg_field AcsmMapTable21_AcsmMapTableVal42;
	rand uvm_reg_field AcsmMapTableVal42;
	rand uvm_reg_field AcsmMapTable21_AcsmMapTableVal43;
	rand uvm_reg_field AcsmMapTableVal43;
	rand uvm_reg_field AcsmMapTable22_AcsmMapTableVal44;
	rand uvm_reg_field AcsmMapTableVal44;
	rand uvm_reg_field AcsmMapTable22_AcsmMapTableVal45;
	rand uvm_reg_field AcsmMapTableVal45;
	rand uvm_reg_field AcsmMapTable23_AcsmMapTableVal46;
	rand uvm_reg_field AcsmMapTableVal46;
	rand uvm_reg_field AcsmMapTable23_AcsmMapTableVal47;
	rand uvm_reg_field AcsmMapTableVal47;
	rand uvm_reg_field AcsmMapTable24_AcsmMapTableVal48;
	rand uvm_reg_field AcsmMapTableVal48;
	rand uvm_reg_field AcsmMapTable24_AcsmMapTableVal49;
	rand uvm_reg_field AcsmMapTableVal49;
	rand uvm_reg_field AcsmMapTable25_AcsmMapTableVal50;
	rand uvm_reg_field AcsmMapTableVal50;
	rand uvm_reg_field AcsmMapTable25_AcsmMapTableVal51;
	rand uvm_reg_field AcsmMapTableVal51;
	rand uvm_reg_field AcsmMapTable26_AcsmMapTableVal52;
	rand uvm_reg_field AcsmMapTableVal52;
	rand uvm_reg_field AcsmMapTable26_AcsmMapTableVal53;
	rand uvm_reg_field AcsmMapTableVal53;
	rand uvm_reg_field AcsmMapTable27_AcsmMapTableVal54;
	rand uvm_reg_field AcsmMapTableVal54;
	rand uvm_reg_field AcsmMapTable27_AcsmMapTableVal55;
	rand uvm_reg_field AcsmMapTableVal55;
	rand uvm_reg_field AcsmMapTable28_AcsmMapTableVal56;
	rand uvm_reg_field AcsmMapTableVal56;
	rand uvm_reg_field AcsmMapTable28_AcsmMapTableVal57;
	rand uvm_reg_field AcsmMapTableVal57;
	rand uvm_reg_field AcsmMapTable29_AcsmMapTableVal58;
	rand uvm_reg_field AcsmMapTableVal58;
	rand uvm_reg_field AcsmMapTable29_AcsmMapTableVal59;
	rand uvm_reg_field AcsmMapTableVal59;
	rand uvm_reg_field AcsmMapTable30_AcsmMapTableVal60;
	rand uvm_reg_field AcsmMapTableVal60;
	rand uvm_reg_field AcsmMapTable30_AcsmMapTableVal61;
	rand uvm_reg_field AcsmMapTableVal61;
	rand uvm_reg_field AcsmMapTable31_AcsmMapTableVal62;
	rand uvm_reg_field AcsmMapTableVal62;
	rand uvm_reg_field AcsmMapTable31_AcsmMapTableVal63;
	rand uvm_reg_field AcsmMapTableVal63;
	rand uvm_reg_field AcsmMapTable32_AcsmMapTableVal64;
	rand uvm_reg_field AcsmMapTableVal64;
	rand uvm_reg_field AcsmMapTable32_AcsmMapTableVal65;
	rand uvm_reg_field AcsmMapTableVal65;
	rand uvm_reg_field AcsmMapTable33_AcsmMapTableVal66;
	rand uvm_reg_field AcsmMapTableVal66;
	rand uvm_reg_field AcsmMapTable33_AcsmMapTableVal67;
	rand uvm_reg_field AcsmMapTableVal67;
	rand uvm_reg_field AcsmMapTable34_AcsmMapTableVal68;
	rand uvm_reg_field AcsmMapTableVal68;
	rand uvm_reg_field AcsmMapTable34_AcsmMapTableVal69;
	rand uvm_reg_field AcsmMapTableVal69;
	rand uvm_reg_field AcsmMapTable35_AcsmMapTableVal70;
	rand uvm_reg_field AcsmMapTableVal70;
	rand uvm_reg_field AcsmMapTable35_AcsmMapTableVal71;
	rand uvm_reg_field AcsmMapTableVal71;
	rand uvm_reg_field AcsmMapTable36_AcsmMapTableVal72;
	rand uvm_reg_field AcsmMapTableVal72;
	rand uvm_reg_field AcsmMapTable36_AcsmMapTableVal73;
	rand uvm_reg_field AcsmMapTableVal73;
	rand uvm_reg_field AcsmMapTable37_AcsmMapTableVal74;
	rand uvm_reg_field AcsmMapTableVal74;
	rand uvm_reg_field AcsmMapTable37_AcsmMapTableVal75;
	rand uvm_reg_field AcsmMapTableVal75;
	rand uvm_reg_field AcsmMapTable38_AcsmMapTableVal76;
	rand uvm_reg_field AcsmMapTableVal76;
	rand uvm_reg_field AcsmMapTable38_AcsmMapTableVal77;
	rand uvm_reg_field AcsmMapTableVal77;
	rand uvm_reg_field AcsmMapTable39_AcsmMapTableVal78;
	rand uvm_reg_field AcsmMapTableVal78;
	rand uvm_reg_field AcsmMapTable39_AcsmMapTableVal79;
	rand uvm_reg_field AcsmMapTableVal79;
	rand uvm_reg_field AcsmMapTable40_AcsmMapTableVal80;
	rand uvm_reg_field AcsmMapTableVal80;
	rand uvm_reg_field AcsmMapTable40_AcsmMapTableVal81;
	rand uvm_reg_field AcsmMapTableVal81;
	rand uvm_reg_field AcsmMapTable41_AcsmMapTableVal82;
	rand uvm_reg_field AcsmMapTableVal82;
	rand uvm_reg_field AcsmMapTable41_AcsmMapTableVal83;
	rand uvm_reg_field AcsmMapTableVal83;
	rand uvm_reg_field AcsmMapTable42_AcsmMapTableVal84;
	rand uvm_reg_field AcsmMapTableVal84;
	rand uvm_reg_field AcsmMapTable42_AcsmMapTableVal85;
	rand uvm_reg_field AcsmMapTableVal85;
	rand uvm_reg_field AcsmMapTable43_AcsmMapTableVal86;
	rand uvm_reg_field AcsmMapTableVal86;
	rand uvm_reg_field AcsmMapTable43_AcsmMapTableVal87;
	rand uvm_reg_field AcsmMapTableVal87;
	rand uvm_reg_field AcsmMapTable44_AcsmMapTableVal88;
	rand uvm_reg_field AcsmMapTableVal88;
	rand uvm_reg_field AcsmMapTable44_AcsmMapTableVal89;
	rand uvm_reg_field AcsmMapTableVal89;
	rand uvm_reg_field AcsmMapTable45_AcsmMapTableVal90;
	rand uvm_reg_field AcsmMapTableVal90;
	rand uvm_reg_field AcsmMapTable45_AcsmMapTableVal91;
	rand uvm_reg_field AcsmMapTableVal91;
	rand uvm_reg_field AcsmMapTable46_AcsmMapTableVal92;
	rand uvm_reg_field AcsmMapTableVal92;
	rand uvm_reg_field AcsmMapTable46_AcsmMapTableVal93;
	rand uvm_reg_field AcsmMapTableVal93;
	rand uvm_reg_field AcsmMapTable47_AcsmMapTableVal94;
	rand uvm_reg_field AcsmMapTableVal94;
	rand uvm_reg_field AcsmMapTable47_AcsmMapTableVal95;
	rand uvm_reg_field AcsmMapTableVal95;
	rand uvm_reg_field AcsmMapTable48_AcsmMapTableVal96;
	rand uvm_reg_field AcsmMapTableVal96;
	rand uvm_reg_field AcsmMapTable48_AcsmMapTableVal97;
	rand uvm_reg_field AcsmMapTableVal97;
	rand uvm_reg_field AcsmMapTable49_AcsmMapTableVal98;
	rand uvm_reg_field AcsmMapTableVal98;
	rand uvm_reg_field AcsmMapTable49_AcsmMapTableVal99;
	rand uvm_reg_field AcsmMapTableVal99;
	rand uvm_reg_field AcsmMapTable50_AcsmMapTableVal100;
	rand uvm_reg_field AcsmMapTableVal100;
	rand uvm_reg_field AcsmMapTable50_AcsmMapTableVal101;
	rand uvm_reg_field AcsmMapTableVal101;
	rand uvm_reg_field AcsmMapTable51_AcsmMapTableVal102;
	rand uvm_reg_field AcsmMapTableVal102;
	rand uvm_reg_field AcsmMapTable51_AcsmMapTableVal103;
	rand uvm_reg_field AcsmMapTableVal103;
	rand uvm_reg_field AcsmMapTable52_AcsmMapTableVal104;
	rand uvm_reg_field AcsmMapTableVal104;
	rand uvm_reg_field AcsmMapTable52_AcsmMapTableVal105;
	rand uvm_reg_field AcsmMapTableVal105;
	rand uvm_reg_field AcsmMapTable53_AcsmMapTableVal106;
	rand uvm_reg_field AcsmMapTableVal106;
	rand uvm_reg_field AcsmMapTable53_AcsmMapTableVal107;
	rand uvm_reg_field AcsmMapTableVal107;
	rand uvm_reg_field AcsmMapTable54_AcsmMapTableVal108;
	rand uvm_reg_field AcsmMapTableVal108;
	rand uvm_reg_field AcsmMapTable54_AcsmMapTableVal109;
	rand uvm_reg_field AcsmMapTableVal109;
	rand uvm_reg_field AcsmMapTable55_AcsmMapTableVal110;
	rand uvm_reg_field AcsmMapTableVal110;
	rand uvm_reg_field AcsmMapTable55_AcsmMapTableVal111;
	rand uvm_reg_field AcsmMapTableVal111;
	rand uvm_reg_field AcsmMapTable56_AcsmMapTableVal112;
	rand uvm_reg_field AcsmMapTableVal112;
	rand uvm_reg_field AcsmMapTable56_AcsmMapTableVal113;
	rand uvm_reg_field AcsmMapTableVal113;
	rand uvm_reg_field AcsmMapTable57_AcsmMapTableVal114;
	rand uvm_reg_field AcsmMapTableVal114;
	rand uvm_reg_field AcsmMapTable57_AcsmMapTableVal115;
	rand uvm_reg_field AcsmMapTableVal115;
	rand uvm_reg_field AcsmMapTable58_AcsmMapTableVal116;
	rand uvm_reg_field AcsmMapTableVal116;
	rand uvm_reg_field AcsmMapTable58_AcsmMapTableVal117;
	rand uvm_reg_field AcsmMapTableVal117;
	rand uvm_reg_field AcsmMapTable59_AcsmMapTableVal118;
	rand uvm_reg_field AcsmMapTableVal118;
	rand uvm_reg_field AcsmMapTable59_AcsmMapTableVal119;
	rand uvm_reg_field AcsmMapTableVal119;
	rand uvm_reg_field AcsmMapTable60_AcsmMapTableVal120;
	rand uvm_reg_field AcsmMapTableVal120;
	rand uvm_reg_field AcsmMapTable60_AcsmMapTableVal121;
	rand uvm_reg_field AcsmMapTableVal121;
	rand uvm_reg_field AcsmMapTable61_AcsmMapTableVal122;
	rand uvm_reg_field AcsmMapTableVal122;
	rand uvm_reg_field AcsmMapTable61_AcsmMapTableVal123;
	rand uvm_reg_field AcsmMapTableVal123;
	rand uvm_reg_field AcsmMapTable62_AcsmMapTableVal124;
	rand uvm_reg_field AcsmMapTableVal124;
	rand uvm_reg_field AcsmMapTable62_AcsmMapTableVal125;
	rand uvm_reg_field AcsmMapTableVal125;
	rand uvm_reg_field AcsmMapTable63_AcsmMapTableVal126;
	rand uvm_reg_field AcsmMapTableVal126;
	rand uvm_reg_field AcsmMapTable63_AcsmMapTableVal127;
	rand uvm_reg_field AcsmMapTableVal127;
	rand uvm_reg_field AcsmStartAddrXlatVal0_AcsmStartAddrXlatVal0;
	rand uvm_reg_field AcsmStartAddrXlatVal1_AcsmStartAddrXlatVal1;
	rand uvm_reg_field AcsmStartAddrXlatVal2_AcsmStartAddrXlatVal2;
	rand uvm_reg_field AcsmStartAddrXlatVal3_AcsmStartAddrXlatVal3;
	rand uvm_reg_field AcsmStartAddrXlatVal4_AcsmStartAddrXlatVal4;
	rand uvm_reg_field AcsmStartAddrXlatVal5_AcsmStartAddrXlatVal5;
	rand uvm_reg_field AcsmStartAddrXlatVal6_AcsmStartAddrXlatVal6;
	rand uvm_reg_field AcsmStartAddrXlatVal7_AcsmStartAddrXlatVal7;
	rand uvm_reg_field AcsmStartAddrXlatVal8_AcsmStartAddrXlatVal8;
	rand uvm_reg_field AcsmStartAddrXlatVal9_AcsmStartAddrXlatVal9;
	rand uvm_reg_field AcsmStartAddrXlatVal10_AcsmStartAddrXlatVal10;
	rand uvm_reg_field AcsmStartAddrXlatVal11_AcsmStartAddrXlatVal11;
	rand uvm_reg_field AcsmStartAddrXlatVal12_AcsmStartAddrXlatVal12;
	rand uvm_reg_field AcsmStartAddrXlatVal13_AcsmStartAddrXlatVal13;
	rand uvm_reg_field AcsmStartAddrXlatVal14_AcsmStartAddrXlatVal14;
	rand uvm_reg_field AcsmStartAddrXlatVal15_AcsmStartAddrXlatVal15;
	rand uvm_reg_field AcsmStartAddrXlatVal16_AcsmStartAddrXlatVal16;
	rand uvm_reg_field AcsmStartAddrXlatVal17_AcsmStartAddrXlatVal17;
	rand uvm_reg_field AcsmStartAddrXlatVal18_AcsmStartAddrXlatVal18;
	rand uvm_reg_field AcsmStartAddrXlatVal19_AcsmStartAddrXlatVal19;
	rand uvm_reg_field AcsmStartAddrXlatVal20_AcsmStartAddrXlatVal20;
	rand uvm_reg_field AcsmStartAddrXlatVal21_AcsmStartAddrXlatVal21;
	rand uvm_reg_field AcsmStartAddrXlatVal22_AcsmStartAddrXlatVal22;
	rand uvm_reg_field AcsmStartAddrXlatVal23_AcsmStartAddrXlatVal23;
	rand uvm_reg_field AcsmStartAddrXlatVal24_AcsmStartAddrXlatVal24;
	rand uvm_reg_field AcsmStartAddrXlatVal25_AcsmStartAddrXlatVal25;
	rand uvm_reg_field AcsmStartAddrXlatVal26_AcsmStartAddrXlatVal26;
	rand uvm_reg_field AcsmStartAddrXlatVal27_AcsmStartAddrXlatVal27;
	rand uvm_reg_field AcsmStartAddrXlatVal28_AcsmStartAddrXlatVal28;
	rand uvm_reg_field AcsmStartAddrXlatVal29_AcsmStartAddrXlatVal29;
	rand uvm_reg_field AcsmStartAddrXlatVal30_AcsmStartAddrXlatVal30;
	rand uvm_reg_field AcsmStartAddrXlatVal31_AcsmStartAddrXlatVal31;
	rand uvm_reg_field AcsmStartAddrXlatVal32_AcsmStartAddrXlatVal32;
	rand uvm_reg_field AcsmStartAddrXlatVal33_AcsmStartAddrXlatVal33;
	rand uvm_reg_field AcsmStartAddrXlatVal34_AcsmStartAddrXlatVal34;
	rand uvm_reg_field AcsmStartAddrXlatVal35_AcsmStartAddrXlatVal35;
	rand uvm_reg_field AcsmStartAddrXlatVal36_AcsmStartAddrXlatVal36;
	rand uvm_reg_field AcsmStartAddrXlatVal37_AcsmStartAddrXlatVal37;
	rand uvm_reg_field AcsmStartAddrXlatVal38_AcsmStartAddrXlatVal38;
	rand uvm_reg_field AcsmStartAddrXlatVal39_AcsmStartAddrXlatVal39;
	rand uvm_reg_field AcsmStartAddrXlatVal40_AcsmStartAddrXlatVal40;
	rand uvm_reg_field AcsmStartAddrXlatVal41_AcsmStartAddrXlatVal41;
	rand uvm_reg_field AcsmStartAddrXlatVal42_AcsmStartAddrXlatVal42;
	rand uvm_reg_field AcsmStartAddrXlatVal43_AcsmStartAddrXlatVal43;
	rand uvm_reg_field AcsmStartAddrXlatVal44_AcsmStartAddrXlatVal44;
	rand uvm_reg_field AcsmStartAddrXlatVal45_AcsmStartAddrXlatVal45;
	rand uvm_reg_field AcsmStartAddrXlatVal46_AcsmStartAddrXlatVal46;
	rand uvm_reg_field AcsmStartAddrXlatVal47_AcsmStartAddrXlatVal47;
	rand uvm_reg_field AcsmStartAddrXlatVal48_AcsmStartAddrXlatVal48;
	rand uvm_reg_field AcsmStartAddrXlatVal49_AcsmStartAddrXlatVal49;
	rand uvm_reg_field AcsmStartAddrXlatVal50_AcsmStartAddrXlatVal50;
	rand uvm_reg_field AcsmStartAddrXlatVal51_AcsmStartAddrXlatVal51;
	rand uvm_reg_field AcsmStartAddrXlatVal52_AcsmStartAddrXlatVal52;
	rand uvm_reg_field AcsmStartAddrXlatVal53_AcsmStartAddrXlatVal53;
	rand uvm_reg_field AcsmStartAddrXlatVal54_AcsmStartAddrXlatVal54;
	rand uvm_reg_field AcsmStartAddrXlatVal55_AcsmStartAddrXlatVal55;
	rand uvm_reg_field AcsmStartAddrXlatVal56_AcsmStartAddrXlatVal56;
	rand uvm_reg_field AcsmStartAddrXlatVal57_AcsmStartAddrXlatVal57;
	rand uvm_reg_field AcsmStartAddrXlatVal58_AcsmStartAddrXlatVal58;
	rand uvm_reg_field AcsmStartAddrXlatVal59_AcsmStartAddrXlatVal59;
	rand uvm_reg_field AcsmStartAddrXlatVal60_AcsmStartAddrXlatVal60;
	rand uvm_reg_field AcsmStartAddrXlatVal61_AcsmStartAddrXlatVal61;
	rand uvm_reg_field AcsmStartAddrXlatVal62_AcsmStartAddrXlatVal62;
	rand uvm_reg_field AcsmStartAddrXlatVal63_AcsmStartAddrXlatVal63;
	rand uvm_reg_field AcsmStopAddrXlatVal0_AcsmStopAddrXlatVal0;
	rand uvm_reg_field AcsmStopAddrXlatVal1_AcsmStopAddrXlatVal1;
	rand uvm_reg_field AcsmStopAddrXlatVal2_AcsmStopAddrXlatVal2;
	rand uvm_reg_field AcsmStopAddrXlatVal3_AcsmStopAddrXlatVal3;
	rand uvm_reg_field AcsmStopAddrXlatVal4_AcsmStopAddrXlatVal4;
	rand uvm_reg_field AcsmStopAddrXlatVal5_AcsmStopAddrXlatVal5;
	rand uvm_reg_field AcsmStopAddrXlatVal6_AcsmStopAddrXlatVal6;
	rand uvm_reg_field AcsmStopAddrXlatVal7_AcsmStopAddrXlatVal7;
	rand uvm_reg_field AcsmStopAddrXlatVal8_AcsmStopAddrXlatVal8;
	rand uvm_reg_field AcsmStopAddrXlatVal9_AcsmStopAddrXlatVal9;
	rand uvm_reg_field AcsmStopAddrXlatVal10_AcsmStopAddrXlatVal10;
	rand uvm_reg_field AcsmStopAddrXlatVal11_AcsmStopAddrXlatVal11;
	rand uvm_reg_field AcsmStopAddrXlatVal12_AcsmStopAddrXlatVal12;
	rand uvm_reg_field AcsmStopAddrXlatVal13_AcsmStopAddrXlatVal13;
	rand uvm_reg_field AcsmStopAddrXlatVal14_AcsmStopAddrXlatVal14;
	rand uvm_reg_field AcsmStopAddrXlatVal15_AcsmStopAddrXlatVal15;
	rand uvm_reg_field AcsmStopAddrXlatVal16_AcsmStopAddrXlatVal16;
	rand uvm_reg_field AcsmStopAddrXlatVal17_AcsmStopAddrXlatVal17;
	rand uvm_reg_field AcsmStopAddrXlatVal18_AcsmStopAddrXlatVal18;
	rand uvm_reg_field AcsmStopAddrXlatVal19_AcsmStopAddrXlatVal19;
	rand uvm_reg_field AcsmStopAddrXlatVal20_AcsmStopAddrXlatVal20;
	rand uvm_reg_field AcsmStopAddrXlatVal21_AcsmStopAddrXlatVal21;
	rand uvm_reg_field AcsmStopAddrXlatVal22_AcsmStopAddrXlatVal22;
	rand uvm_reg_field AcsmStopAddrXlatVal23_AcsmStopAddrXlatVal23;
	rand uvm_reg_field AcsmStopAddrXlatVal24_AcsmStopAddrXlatVal24;
	rand uvm_reg_field AcsmStopAddrXlatVal25_AcsmStopAddrXlatVal25;
	rand uvm_reg_field AcsmStopAddrXlatVal26_AcsmStopAddrXlatVal26;
	rand uvm_reg_field AcsmStopAddrXlatVal27_AcsmStopAddrXlatVal27;
	rand uvm_reg_field AcsmStopAddrXlatVal28_AcsmStopAddrXlatVal28;
	rand uvm_reg_field AcsmStopAddrXlatVal29_AcsmStopAddrXlatVal29;
	rand uvm_reg_field AcsmStopAddrXlatVal30_AcsmStopAddrXlatVal30;
	rand uvm_reg_field AcsmStopAddrXlatVal31_AcsmStopAddrXlatVal31;
	rand uvm_reg_field AcsmStopAddrXlatVal32_AcsmStopAddrXlatVal32;
	rand uvm_reg_field AcsmStopAddrXlatVal33_AcsmStopAddrXlatVal33;
	rand uvm_reg_field AcsmStopAddrXlatVal34_AcsmStopAddrXlatVal34;
	rand uvm_reg_field AcsmStopAddrXlatVal35_AcsmStopAddrXlatVal35;
	rand uvm_reg_field AcsmStopAddrXlatVal36_AcsmStopAddrXlatVal36;
	rand uvm_reg_field AcsmStopAddrXlatVal37_AcsmStopAddrXlatVal37;
	rand uvm_reg_field AcsmStopAddrXlatVal38_AcsmStopAddrXlatVal38;
	rand uvm_reg_field AcsmStopAddrXlatVal39_AcsmStopAddrXlatVal39;
	rand uvm_reg_field AcsmStopAddrXlatVal40_AcsmStopAddrXlatVal40;
	rand uvm_reg_field AcsmStopAddrXlatVal41_AcsmStopAddrXlatVal41;
	rand uvm_reg_field AcsmStopAddrXlatVal42_AcsmStopAddrXlatVal42;
	rand uvm_reg_field AcsmStopAddrXlatVal43_AcsmStopAddrXlatVal43;
	rand uvm_reg_field AcsmStopAddrXlatVal44_AcsmStopAddrXlatVal44;
	rand uvm_reg_field AcsmStopAddrXlatVal45_AcsmStopAddrXlatVal45;
	rand uvm_reg_field AcsmStopAddrXlatVal46_AcsmStopAddrXlatVal46;
	rand uvm_reg_field AcsmStopAddrXlatVal47_AcsmStopAddrXlatVal47;
	rand uvm_reg_field AcsmStopAddrXlatVal48_AcsmStopAddrXlatVal48;
	rand uvm_reg_field AcsmStopAddrXlatVal49_AcsmStopAddrXlatVal49;
	rand uvm_reg_field AcsmStopAddrXlatVal50_AcsmStopAddrXlatVal50;
	rand uvm_reg_field AcsmStopAddrXlatVal51_AcsmStopAddrXlatVal51;
	rand uvm_reg_field AcsmStopAddrXlatVal52_AcsmStopAddrXlatVal52;
	rand uvm_reg_field AcsmStopAddrXlatVal53_AcsmStopAddrXlatVal53;
	rand uvm_reg_field AcsmStopAddrXlatVal54_AcsmStopAddrXlatVal54;
	rand uvm_reg_field AcsmStopAddrXlatVal55_AcsmStopAddrXlatVal55;
	rand uvm_reg_field AcsmStopAddrXlatVal56_AcsmStopAddrXlatVal56;
	rand uvm_reg_field AcsmStopAddrXlatVal57_AcsmStopAddrXlatVal57;
	rand uvm_reg_field AcsmStopAddrXlatVal58_AcsmStopAddrXlatVal58;
	rand uvm_reg_field AcsmStopAddrXlatVal59_AcsmStopAddrXlatVal59;
	rand uvm_reg_field AcsmStopAddrXlatVal60_AcsmStopAddrXlatVal60;
	rand uvm_reg_field AcsmStopAddrXlatVal61_AcsmStopAddrXlatVal61;
	rand uvm_reg_field AcsmStopAddrXlatVal62_AcsmStopAddrXlatVal62;
	rand uvm_reg_field AcsmStopAddrXlatVal63_AcsmStopAddrXlatVal63;


	covergroup cg_addr (input string name);
	option.per_instance = 1;
option.name = get_name();

	PpgcGenCtrl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h0 };
		option.weight = 1;
	}

	PpgcGenDbiCtrl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1 };
		option.weight = 1;
	}

	PpgcGenDbiConfig : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2 };
		option.weight = 1;
	}

	PpgcGenLaneMuxSel0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3 };
		option.weight = 1;
	}

	PpgcGenLaneMuxSel1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h4 };
		option.weight = 1;
	}

	EnPhyUpdZQCalUpdate : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h5 };
		option.weight = 1;
	}

	BlockDfiInterface : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6 };
		option.weight = 1;
	}

	BlockDfiInterfaceStatus : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h7 };
		option.weight = 1;
	}

	DfiCustMode_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hB };
		option.weight = 1;
	}

	HwtMRL_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hD };
		option.weight = 1;
	}

	RegRet : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE };
		option.weight = 1;
	}

	DisableZQupdateOnSnoop : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hF };
		option.weight = 1;
	}

	Prbs0GenModeSel : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h10 };
		option.weight = 1;
	}

	Prbs0GenUiMuxSel : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h11 };
		option.weight = 1;
	}

	Prbs0GenTapDly0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h12 };
		option.weight = 1;
	}

	Prbs0GenTapDly1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h13 };
		option.weight = 1;
	}

	Prbs0GenTapDly2 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h14 };
		option.weight = 1;
	}

	Prbs0GenTapDly3 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h15 };
		option.weight = 1;
	}

	Prbs0GenTapDly4 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h16 };
		option.weight = 1;
	}

	Prbs0GenTapDly5 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h17 };
		option.weight = 1;
	}

	Prbs0GenTapDly6 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h18 };
		option.weight = 1;
	}

	Prbs0GenTapDly7 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h19 };
		option.weight = 1;
	}

	MtestMuxSel : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1A };
		option.weight = 1;
	}

	Prbs0GenStateLo : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1B };
		option.weight = 1;
	}

	Prbs0GenStateHi : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1C };
		option.weight = 1;
	}

	Prbs1GenModeSel : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20 };
		option.weight = 1;
	}

	Prbs1GenUiMuxSel : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h21 };
		option.weight = 1;
	}

	Prbs1GenTapDly0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h22 };
		option.weight = 1;
	}

	Prbs1GenTapDly1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h23 };
		option.weight = 1;
	}

	Prbs1GenTapDly2 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h24 };
		option.weight = 1;
	}

	Prbs1GenTapDly3 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h25 };
		option.weight = 1;
	}

	Prbs1GenTapDly4 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h26 };
		option.weight = 1;
	}

	Prbs1GenTapDly5 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h27 };
		option.weight = 1;
	}

	Prbs1GenTapDly6 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h28 };
		option.weight = 1;
	}

	Prbs1GenTapDly7 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h29 };
		option.weight = 1;
	}

	Prbs1GenStateLo : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2B };
		option.weight = 1;
	}

	Prbs1GenStateHi : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2C };
		option.weight = 1;
	}

	Prbs2GenModeSel : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h30 };
		option.weight = 1;
	}

	Prbs2GenUiMuxSel : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h31 };
		option.weight = 1;
	}

	Prbs2GenTapDly0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h32 };
		option.weight = 1;
	}

	Prbs2GenTapDly1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h33 };
		option.weight = 1;
	}

	Prbs2GenTapDly2 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h34 };
		option.weight = 1;
	}

	Prbs2GenTapDly3 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h35 };
		option.weight = 1;
	}

	Prbs2GenTapDly4 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h36 };
		option.weight = 1;
	}

	Prbs2GenTapDly5 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h37 };
		option.weight = 1;
	}

	Prbs2GenTapDly6 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h38 };
		option.weight = 1;
	}

	Prbs2GenTapDly7 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h39 };
		option.weight = 1;
	}

	Prbs2GenStateLo : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B };
		option.weight = 1;
	}

	Prbs2GenStateHi : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C };
		option.weight = 1;
	}

	PPTTrainSetup_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h40 };
		option.weight = 1;
	}

	PhyMstrFreqOverride_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h41 };
		option.weight = 1;
	}

	DfiInitComplete : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h49 };
		option.weight = 1;
	}

	PPGCParityInvert : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h4D };
		option.weight = 1;
	}

	PMIEnable : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h54 };
		option.weight = 1;
	}

	Dfi0Status : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h5A };
		option.weight = 1;
	}

	Dfi1Status : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h5B };
		option.weight = 1;
	}

	DfiHandshakeDelays0_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h66 };
		option.weight = 1;
	}

	DFIPHYUPD0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h67 };
		option.weight = 1;
	}

	DfiLpCtrlEn0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h68 };
		option.weight = 1;
	}

	DfiLpDataEn0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h69 };
		option.weight = 1;
	}

	DynOdtEnCntrl0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6A };
		option.weight = 1;
	}

	DfiRespHandshakeDelays0_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6B };
		option.weight = 1;
	}

	HwtLpCsEnA : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h72 };
		option.weight = 1;
	}

	HwtLpCsEnB : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h73 };
		option.weight = 1;
	}

	HwtCtrl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h77 };
		option.weight = 1;
	}

	HwtControlOvr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h7A };
		option.weight = 1;
	}

	ScratchPadPPGC : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h7D };
		option.weight = 1;
	}

	HwtControlVal : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h7E };
		option.weight = 1;
	}

	ForceHWTClkGaterEnables : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h80 };
		option.weight = 1;
	}

	MasUpdGoodCtr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hB5 };
		option.weight = 1;
	}

	PhyUpd0GoodCtr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hB6 };
		option.weight = 1;
	}

	PhyUpd1GoodCtr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hB7 };
		option.weight = 1;
	}

	CtlUpd0GoodCtr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hB8 };
		option.weight = 1;
	}

	CtlUpd1GoodCtr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hB9 };
		option.weight = 1;
	}

	MasUpdFailCtr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hBA };
		option.weight = 1;
	}

	PhyUpd0FailCtr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hBB };
		option.weight = 1;
	}

	PhyUpd1FailCtr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hBC };
		option.weight = 1;
	}

	PhyPerfCtrEnable : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hBD };
		option.weight = 1;
	}

	DfiHandshakeDelays1_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE6 };
		option.weight = 1;
	}

	DFIPHYUPD1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE7 };
		option.weight = 1;
	}

	DfiLpCtrlEn1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE8 };
		option.weight = 1;
	}

	DfiLpDataEn1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE9 };
		option.weight = 1;
	}

	DynOdtEnCntrl1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hEA };
		option.weight = 1;
	}

	DfiRespHandshakeDelays1_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hEB };
		option.weight = 1;
	}

	FspSkipList : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hF0 };
		option.weight = 1;
	}

	PPGCReserved0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hFA };
		option.weight = 1;
	}

	PUBReservedP1_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hFF };
		option.weight = 1;
	}

	PhyInterruptOverride : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h11A };
		option.weight = 1;
	}

	PhyInterruptEnable : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h11B };
		option.weight = 1;
	}

	PhyInterruptFWControl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h11C };
		option.weight = 1;
	}

	PhyInterruptMask : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h11D };
		option.weight = 1;
	}

	PhyInterruptClear : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h11E };
		option.weight = 1;
	}

	PhyInterruptStatus : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h11F };
		option.weight = 1;
	}

	ACSMRunCtrl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h120 };
		option.weight = 1;
	}

	ACSMDone : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h121 };
		option.weight = 1;
	}

	ACSMStartAddr_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h122 };
		option.weight = 1;
	}

	ACSMStopAddr_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h123 };
		option.weight = 1;
	}

	ACSMLastAddr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h124 };
		option.weight = 1;
	}

	ACSMAlgaIncVal : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h125 };
		option.weight = 1;
	}

	ACSMAddressMask : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h126 };
		option.weight = 1;
	}

	ACSMOuterLoopRepeatCnt : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h127 };
		option.weight = 1;
	}

	ACSMCkeControl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h128 };
		option.weight = 1;
	}

	ACSMCkeStatus : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h129 };
		option.weight = 1;
	}

	ACSMWckEnControl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h12A };
		option.weight = 1;
	}

	ACSMWckEnStatus : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h12B };
		option.weight = 1;
	}

	ACSMRxEnPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h12C };
		option.weight = 1;
	}

	ACSMRxValPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h12D };
		option.weight = 1;
	}

	ACSMTxEnPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h12E };
		option.weight = 1;
	}

	ACSMWrcsPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h12F };
		option.weight = 1;
	}

	ACSMRdcsPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h130 };
		option.weight = 1;
	}

	ACSMInfiniteOLRC : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h131 };
		option.weight = 1;
	}

	ACSMDefaultAddr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h132 };
		option.weight = 1;
	}

	ACSMDefaultCs : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h133 };
		option.weight = 1;
	}

	ACSMStaticCtrl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h134 };
		option.weight = 1;
	}

	ACSMWckWriteStaticLoPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h135 };
		option.weight = 1;
	}

	ACSMWckWriteStaticHiPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h136 };
		option.weight = 1;
	}

	ACSMWckWriteTogglePulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h137 };
		option.weight = 1;
	}

	ACSMWckWriteFastTogglePulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h138 };
		option.weight = 1;
	}

	ACSMWckReadStaticLoPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h139 };
		option.weight = 1;
	}

	ACSMWckReadStaticHiPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h13A };
		option.weight = 1;
	}

	ACSMWckReadTogglePulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h13B };
		option.weight = 1;
	}

	ACSMWckReadFastTogglePulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h13C };
		option.weight = 1;
	}

	ACSMWckFreqSwStaticLoPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h13D };
		option.weight = 1;
	}

	ACSMWckFreqSwStaticHiPulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h13E };
		option.weight = 1;
	}

	ACSMWckFreqSwTogglePulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h13F };
		option.weight = 1;
	}

	ACSMWckFreqSwFastTogglePulse_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h140 };
		option.weight = 1;
	}

	ACSMWckFreeRunMode_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h141 };
		option.weight = 1;
	}

	ACSMLowSpeedClockEnable : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h142 };
		option.weight = 1;
	}

	ACSMLowSpeedClockDelay : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h144 };
		option.weight = 1;
	}

	ACSMRptCntOverride_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h145 };
		option.weight = 1;
	}

	ACSMRptCntDbl_p0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h146 };
		option.weight = 1;
	}

	ACSMParityStatus : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h147 };
		option.weight = 1;
	}

	HwtLpCsEnBypass : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h174 };
		option.weight = 1;
	}

	ACSMNopAddr : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h18A };
		option.weight = 1;
	}

	SnoopCntrl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1A7 };
		option.weight = 1;
	}

	ACSMParityInvert : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1A8 };
		option.weight = 1;
	}

	AcsmPsIndx : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1A9 };
		option.weight = 1;
	}

	AcsmDynPtrCtrl : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1AA };
		option.weight = 1;
	}

	FspState : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1EF };
		option.weight = 1;
	}

	AcsmMapTable0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h200 };
		option.weight = 1;
	}

	AcsmMapTable1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h201 };
		option.weight = 1;
	}

	AcsmMapTable2 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h202 };
		option.weight = 1;
	}

	AcsmMapTable3 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h203 };
		option.weight = 1;
	}

	AcsmMapTable4 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h204 };
		option.weight = 1;
	}

	AcsmMapTable5 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h205 };
		option.weight = 1;
	}

	AcsmMapTable6 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h206 };
		option.weight = 1;
	}

	AcsmMapTable7 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h207 };
		option.weight = 1;
	}

	AcsmMapTable8 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h208 };
		option.weight = 1;
	}

	AcsmMapTable9 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h209 };
		option.weight = 1;
	}

	AcsmMapTable10 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20A };
		option.weight = 1;
	}

	AcsmMapTable11 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20B };
		option.weight = 1;
	}

	AcsmMapTable12 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20C };
		option.weight = 1;
	}

	AcsmMapTable13 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20D };
		option.weight = 1;
	}

	AcsmMapTable14 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20E };
		option.weight = 1;
	}

	AcsmMapTable15 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20F };
		option.weight = 1;
	}

	AcsmMapTable16 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h210 };
		option.weight = 1;
	}

	AcsmMapTable17 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h211 };
		option.weight = 1;
	}

	AcsmMapTable18 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h212 };
		option.weight = 1;
	}

	AcsmMapTable19 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h213 };
		option.weight = 1;
	}

	AcsmMapTable20 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h214 };
		option.weight = 1;
	}

	AcsmMapTable21 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h215 };
		option.weight = 1;
	}

	AcsmMapTable22 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h216 };
		option.weight = 1;
	}

	AcsmMapTable23 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h217 };
		option.weight = 1;
	}

	AcsmMapTable24 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h218 };
		option.weight = 1;
	}

	AcsmMapTable25 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h219 };
		option.weight = 1;
	}

	AcsmMapTable26 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h21A };
		option.weight = 1;
	}

	AcsmMapTable27 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h21B };
		option.weight = 1;
	}

	AcsmMapTable28 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h21C };
		option.weight = 1;
	}

	AcsmMapTable29 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h21D };
		option.weight = 1;
	}

	AcsmMapTable30 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h21E };
		option.weight = 1;
	}

	AcsmMapTable31 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h21F };
		option.weight = 1;
	}

	AcsmMapTable32 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h220 };
		option.weight = 1;
	}

	AcsmMapTable33 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h221 };
		option.weight = 1;
	}

	AcsmMapTable34 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h222 };
		option.weight = 1;
	}

	AcsmMapTable35 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h223 };
		option.weight = 1;
	}

	AcsmMapTable36 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h224 };
		option.weight = 1;
	}

	AcsmMapTable37 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h225 };
		option.weight = 1;
	}

	AcsmMapTable38 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h226 };
		option.weight = 1;
	}

	AcsmMapTable39 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h227 };
		option.weight = 1;
	}

	AcsmMapTable40 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h228 };
		option.weight = 1;
	}

	AcsmMapTable41 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h229 };
		option.weight = 1;
	}

	AcsmMapTable42 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h22A };
		option.weight = 1;
	}

	AcsmMapTable43 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h22B };
		option.weight = 1;
	}

	AcsmMapTable44 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h22C };
		option.weight = 1;
	}

	AcsmMapTable45 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h22D };
		option.weight = 1;
	}

	AcsmMapTable46 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h22E };
		option.weight = 1;
	}

	AcsmMapTable47 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h22F };
		option.weight = 1;
	}

	AcsmMapTable48 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h230 };
		option.weight = 1;
	}

	AcsmMapTable49 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h231 };
		option.weight = 1;
	}

	AcsmMapTable50 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h232 };
		option.weight = 1;
	}

	AcsmMapTable51 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h233 };
		option.weight = 1;
	}

	AcsmMapTable52 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h234 };
		option.weight = 1;
	}

	AcsmMapTable53 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h235 };
		option.weight = 1;
	}

	AcsmMapTable54 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h236 };
		option.weight = 1;
	}

	AcsmMapTable55 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h237 };
		option.weight = 1;
	}

	AcsmMapTable56 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h238 };
		option.weight = 1;
	}

	AcsmMapTable57 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h239 };
		option.weight = 1;
	}

	AcsmMapTable58 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h23A };
		option.weight = 1;
	}

	AcsmMapTable59 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h23B };
		option.weight = 1;
	}

	AcsmMapTable60 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h23C };
		option.weight = 1;
	}

	AcsmMapTable61 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h23D };
		option.weight = 1;
	}

	AcsmMapTable62 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h23E };
		option.weight = 1;
	}

	AcsmMapTable63 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h23F };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h324 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h325 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal2 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h326 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal3 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h327 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal4 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h328 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal5 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h329 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal6 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h32A };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal7 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h32B };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal8 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h32C };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal9 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h32D };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal10 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h32E };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal11 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h32F };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal12 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h330 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal13 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h331 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal14 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h332 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal15 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h333 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal16 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h334 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal17 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h335 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal18 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h336 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal19 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h337 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal20 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h338 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal21 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h339 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal22 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h33A };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal23 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h33B };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal24 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h33C };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal25 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h33D };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal26 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h33E };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal27 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h33F };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal28 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h340 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal29 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h341 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal30 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h342 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal31 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h343 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal32 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h344 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal33 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h345 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal34 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h346 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal35 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h347 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal36 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h348 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal37 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h349 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal38 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h34A };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal39 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h34B };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal40 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h34C };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal41 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h34D };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal42 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h34E };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal43 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h34F };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal44 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h350 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal45 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h351 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal46 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h352 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal47 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h353 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal48 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h354 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal49 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h355 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal50 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h356 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal51 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h357 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal52 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h358 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal53 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h359 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal54 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h35A };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal55 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h35B };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal56 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h35C };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal57 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h35D };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal58 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h35E };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal59 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h35F };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal60 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h360 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal61 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h361 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal62 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h362 };
		option.weight = 1;
	}

	AcsmStartAddrXlatVal63 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h363 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h38B };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h38C };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal2 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h38D };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal3 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h38E };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal4 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h38F };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal5 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h390 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal6 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h391 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal7 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h392 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal8 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h393 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal9 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h394 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal10 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h395 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal11 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h396 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal12 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h397 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal13 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h398 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal14 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h399 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal15 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h39A };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal16 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h39B };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal17 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h39C };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal18 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h39D };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal19 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h39E };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal20 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h39F };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal21 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A0 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal22 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A1 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal23 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A2 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal24 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A3 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal25 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A4 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal26 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A5 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal27 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A6 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal28 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A7 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal29 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A8 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal30 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3A9 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal31 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3AA };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal32 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3AB };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal33 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3AC };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal34 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3AD };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal35 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3AE };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal36 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3AF };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal37 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B0 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal38 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B1 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal39 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B2 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal40 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B3 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal41 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B4 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal42 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B5 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal43 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B6 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal44 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B7 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal45 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B8 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal46 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3B9 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal47 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3BA };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal48 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3BB };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal49 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3BC };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal50 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3BD };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal51 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3BE };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal52 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3BF };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal53 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C0 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal54 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C1 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal55 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C2 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal56 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C3 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal57 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C4 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal58 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C5 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal59 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C6 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal60 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C7 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal61 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C8 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal62 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C9 };
		option.weight = 1;
	}

	AcsmStopAddrXlatVal63 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3CA };
		option.weight = 1;
	}
endgroup
	function new(string name = "DWC_DDRPHYA_PPGC0_p0");
		super.new(name, build_coverage(UVM_CVR_ADDR_MAP));
		add_coverage(build_coverage(UVM_CVR_ADDR_MAP));
		if (has_coverage(UVM_CVR_ADDR_MAP))
			cg_addr = new("cg_addr");
	endfunction: new

   virtual function void build();
      this.default_map = create_map("", 0, 4, UVM_LITTLE_ENDIAN, 0);
      this.PpgcGenCtrl = ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenCtrl::type_id::create("PpgcGenCtrl",,get_full_name());
      if(this.PpgcGenCtrl.has_coverage(UVM_CVR_ALL))
      	this.PpgcGenCtrl.cg_bits.option.name = {get_name(), ".", "PpgcGenCtrl_bits"};
      this.PpgcGenCtrl.configure(this, null, "");
      this.PpgcGenCtrl.build();
      this.default_map.add_reg(this.PpgcGenCtrl, `UVM_REG_ADDR_WIDTH'h0, "RW", 0);
		this.PpgcGenCtrl_PpgcGenCtrl = this.PpgcGenCtrl.PpgcGenCtrl;
      this.PpgcGenDbiCtrl = ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiCtrl::type_id::create("PpgcGenDbiCtrl",,get_full_name());
      if(this.PpgcGenDbiCtrl.has_coverage(UVM_CVR_ALL))
      	this.PpgcGenDbiCtrl.cg_bits.option.name = {get_name(), ".", "PpgcGenDbiCtrl_bits"};
      this.PpgcGenDbiCtrl.configure(this, null, "");
      this.PpgcGenDbiCtrl.build();
      this.default_map.add_reg(this.PpgcGenDbiCtrl, `UVM_REG_ADDR_WIDTH'h1, "RW", 0);
		this.PpgcGenDbiCtrl_PpgcGenDbiCtrl = this.PpgcGenDbiCtrl.PpgcGenDbiCtrl;
      this.PpgcGenDbiConfig = ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenDbiConfig::type_id::create("PpgcGenDbiConfig",,get_full_name());
      if(this.PpgcGenDbiConfig.has_coverage(UVM_CVR_ALL))
      	this.PpgcGenDbiConfig.cg_bits.option.name = {get_name(), ".", "PpgcGenDbiConfig_bits"};
      this.PpgcGenDbiConfig.configure(this, null, "");
      this.PpgcGenDbiConfig.build();
      this.default_map.add_reg(this.PpgcGenDbiConfig, `UVM_REG_ADDR_WIDTH'h2, "RW", 0);
		this.PpgcGenDbiConfig_PpgcGenDbiConfig = this.PpgcGenDbiConfig.PpgcGenDbiConfig;
      this.PpgcGenLaneMuxSel0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel0::type_id::create("PpgcGenLaneMuxSel0",,get_full_name());
      if(this.PpgcGenLaneMuxSel0.has_coverage(UVM_CVR_ALL))
      	this.PpgcGenLaneMuxSel0.cg_bits.option.name = {get_name(), ".", "PpgcGenLaneMuxSel0_bits"};
      this.PpgcGenLaneMuxSel0.configure(this, null, "");
      this.PpgcGenLaneMuxSel0.build();
      this.default_map.add_reg(this.PpgcGenLaneMuxSel0, `UVM_REG_ADDR_WIDTH'h3, "RW", 0);
		this.PpgcGenLaneMuxSel0_PpgcGenLaneMuxSel0 = this.PpgcGenLaneMuxSel0.PpgcGenLaneMuxSel0;
      this.PpgcGenLaneMuxSel1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_PpgcGenLaneMuxSel1::type_id::create("PpgcGenLaneMuxSel1",,get_full_name());
      if(this.PpgcGenLaneMuxSel1.has_coverage(UVM_CVR_ALL))
      	this.PpgcGenLaneMuxSel1.cg_bits.option.name = {get_name(), ".", "PpgcGenLaneMuxSel1_bits"};
      this.PpgcGenLaneMuxSel1.configure(this, null, "");
      this.PpgcGenLaneMuxSel1.build();
      this.default_map.add_reg(this.PpgcGenLaneMuxSel1, `UVM_REG_ADDR_WIDTH'h4, "RW", 0);
		this.PpgcGenLaneMuxSel1_PpgcGenLaneMuxSel1 = this.PpgcGenLaneMuxSel1.PpgcGenLaneMuxSel1;
      this.EnPhyUpdZQCalUpdate = ral_reg_DWC_DDRPHYA_PPGC0_p0_EnPhyUpdZQCalUpdate::type_id::create("EnPhyUpdZQCalUpdate",,get_full_name());
      if(this.EnPhyUpdZQCalUpdate.has_coverage(UVM_CVR_ALL))
      	this.EnPhyUpdZQCalUpdate.cg_bits.option.name = {get_name(), ".", "EnPhyUpdZQCalUpdate_bits"};
      this.EnPhyUpdZQCalUpdate.configure(this, null, "");
      this.EnPhyUpdZQCalUpdate.build();
      this.default_map.add_reg(this.EnPhyUpdZQCalUpdate, `UVM_REG_ADDR_WIDTH'h5, "RW", 0);
		this.EnPhyUpdZQCalUpdate_EnPhyUpdZQCalUpdate = this.EnPhyUpdZQCalUpdate.EnPhyUpdZQCalUpdate;
      this.BlockDfiInterface = ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterface::type_id::create("BlockDfiInterface",,get_full_name());
      if(this.BlockDfiInterface.has_coverage(UVM_CVR_ALL))
      	this.BlockDfiInterface.cg_bits.option.name = {get_name(), ".", "BlockDfiInterface_bits"};
      this.BlockDfiInterface.configure(this, null, "");
      this.BlockDfiInterface.build();
      this.default_map.add_reg(this.BlockDfiInterface, `UVM_REG_ADDR_WIDTH'h6, "RW", 0);
		this.BlockDfiInterface_BlockDfiInterfaceEn = this.BlockDfiInterface.BlockDfiInterfaceEn;
		this.BlockDfiInterfaceEn = this.BlockDfiInterface.BlockDfiInterfaceEn;
		this.BlockDfiInterface_BlockDfiInterfaceStatusReset = this.BlockDfiInterface.BlockDfiInterfaceStatusReset;
		this.BlockDfiInterfaceStatusReset = this.BlockDfiInterface.BlockDfiInterfaceStatusReset;
		this.BlockDfiInterface_PmuBusy = this.BlockDfiInterface.PmuBusy;
		this.PmuBusy = this.BlockDfiInterface.PmuBusy;
      this.BlockDfiInterfaceStatus = ral_reg_DWC_DDRPHYA_PPGC0_p0_BlockDfiInterfaceStatus::type_id::create("BlockDfiInterfaceStatus",,get_full_name());
      if(this.BlockDfiInterfaceStatus.has_coverage(UVM_CVR_ALL))
      	this.BlockDfiInterfaceStatus.cg_bits.option.name = {get_name(), ".", "BlockDfiInterfaceStatus_bits"};
      this.BlockDfiInterfaceStatus.configure(this, null, "");
      this.BlockDfiInterfaceStatus.build();
      this.default_map.add_reg(this.BlockDfiInterfaceStatus, `UVM_REG_ADDR_WIDTH'h7, "RO", 0);
		this.BlockDfiInterfaceStatus_BlockDfiInterfaceStatus = this.BlockDfiInterfaceStatus.BlockDfiInterfaceStatus;
      this.DfiCustMode_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiCustMode_p0::type_id::create("DfiCustMode_p0",,get_full_name());
      if(this.DfiCustMode_p0.has_coverage(UVM_CVR_ALL))
      	this.DfiCustMode_p0.cg_bits.option.name = {get_name(), ".", "DfiCustMode_p0_bits"};
      this.DfiCustMode_p0.configure(this, null, "");
      this.DfiCustMode_p0.build();
      this.default_map.add_reg(this.DfiCustMode_p0, `UVM_REG_ADDR_WIDTH'hB, "RW", 0);
		this.DfiCustMode_p0_DfiCustMode_p0 = this.DfiCustMode_p0.DfiCustMode_p0;
      this.HwtMRL_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtMRL_p0::type_id::create("HwtMRL_p0",,get_full_name());
      if(this.HwtMRL_p0.has_coverage(UVM_CVR_ALL))
      	this.HwtMRL_p0.cg_bits.option.name = {get_name(), ".", "HwtMRL_p0_bits"};
      this.HwtMRL_p0.configure(this, null, "");
      this.HwtMRL_p0.build();
      this.default_map.add_reg(this.HwtMRL_p0, `UVM_REG_ADDR_WIDTH'hD, "RW", 0);
		this.HwtMRL_p0_HwtMRL_p0 = this.HwtMRL_p0.HwtMRL_p0;
      this.RegRet = ral_reg_DWC_DDRPHYA_PPGC0_p0_RegRet::type_id::create("RegRet",,get_full_name());
      if(this.RegRet.has_coverage(UVM_CVR_ALL))
      	this.RegRet.cg_bits.option.name = {get_name(), ".", "RegRet_bits"};
      this.RegRet.configure(this, null, "");
      this.RegRet.build();
      this.default_map.add_reg(this.RegRet, `UVM_REG_ADDR_WIDTH'hE, "RW", 0);
		this.RegRet_RegRet = this.RegRet.RegRet;
      this.DisableZQupdateOnSnoop = ral_reg_DWC_DDRPHYA_PPGC0_p0_DisableZQupdateOnSnoop::type_id::create("DisableZQupdateOnSnoop",,get_full_name());
      if(this.DisableZQupdateOnSnoop.has_coverage(UVM_CVR_ALL))
      	this.DisableZQupdateOnSnoop.cg_bits.option.name = {get_name(), ".", "DisableZQupdateOnSnoop_bits"};
      this.DisableZQupdateOnSnoop.configure(this, null, "");
      this.DisableZQupdateOnSnoop.build();
      this.default_map.add_reg(this.DisableZQupdateOnSnoop, `UVM_REG_ADDR_WIDTH'hF, "RW", 0);
		this.DisableZQupdateOnSnoop_DisableZQupdateOnSnoop = this.DisableZQupdateOnSnoop.DisableZQupdateOnSnoop;
      this.Prbs0GenModeSel = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenModeSel::type_id::create("Prbs0GenModeSel",,get_full_name());
      if(this.Prbs0GenModeSel.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenModeSel.cg_bits.option.name = {get_name(), ".", "Prbs0GenModeSel_bits"};
      this.Prbs0GenModeSel.configure(this, null, "");
      this.Prbs0GenModeSel.build();
      this.default_map.add_reg(this.Prbs0GenModeSel, `UVM_REG_ADDR_WIDTH'h10, "RW", 0);
		this.Prbs0GenModeSel_Prbs0GenModeSel = this.Prbs0GenModeSel.Prbs0GenModeSel;
      this.Prbs0GenUiMuxSel = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenUiMuxSel::type_id::create("Prbs0GenUiMuxSel",,get_full_name());
      if(this.Prbs0GenUiMuxSel.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenUiMuxSel.cg_bits.option.name = {get_name(), ".", "Prbs0GenUiMuxSel_bits"};
      this.Prbs0GenUiMuxSel.configure(this, null, "");
      this.Prbs0GenUiMuxSel.build();
      this.default_map.add_reg(this.Prbs0GenUiMuxSel, `UVM_REG_ADDR_WIDTH'h11, "RW", 0);
		this.Prbs0GenUiMuxSel_Prbs0GenUiMuxSel = this.Prbs0GenUiMuxSel.Prbs0GenUiMuxSel;
      this.Prbs0GenTapDly0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly0::type_id::create("Prbs0GenTapDly0",,get_full_name());
      if(this.Prbs0GenTapDly0.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenTapDly0.cg_bits.option.name = {get_name(), ".", "Prbs0GenTapDly0_bits"};
      this.Prbs0GenTapDly0.configure(this, null, "");
      this.Prbs0GenTapDly0.build();
      this.default_map.add_reg(this.Prbs0GenTapDly0, `UVM_REG_ADDR_WIDTH'h12, "RW", 0);
		this.Prbs0GenTapDly0_Prbs0GenTapDly0 = this.Prbs0GenTapDly0.Prbs0GenTapDly0;
      this.Prbs0GenTapDly1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly1::type_id::create("Prbs0GenTapDly1",,get_full_name());
      if(this.Prbs0GenTapDly1.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenTapDly1.cg_bits.option.name = {get_name(), ".", "Prbs0GenTapDly1_bits"};
      this.Prbs0GenTapDly1.configure(this, null, "");
      this.Prbs0GenTapDly1.build();
      this.default_map.add_reg(this.Prbs0GenTapDly1, `UVM_REG_ADDR_WIDTH'h13, "RW", 0);
		this.Prbs0GenTapDly1_Prbs0GenTapDly1 = this.Prbs0GenTapDly1.Prbs0GenTapDly1;
      this.Prbs0GenTapDly2 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly2::type_id::create("Prbs0GenTapDly2",,get_full_name());
      if(this.Prbs0GenTapDly2.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenTapDly2.cg_bits.option.name = {get_name(), ".", "Prbs0GenTapDly2_bits"};
      this.Prbs0GenTapDly2.configure(this, null, "");
      this.Prbs0GenTapDly2.build();
      this.default_map.add_reg(this.Prbs0GenTapDly2, `UVM_REG_ADDR_WIDTH'h14, "RW", 0);
		this.Prbs0GenTapDly2_Prbs0GenTapDly2 = this.Prbs0GenTapDly2.Prbs0GenTapDly2;
      this.Prbs0GenTapDly3 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly3::type_id::create("Prbs0GenTapDly3",,get_full_name());
      if(this.Prbs0GenTapDly3.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenTapDly3.cg_bits.option.name = {get_name(), ".", "Prbs0GenTapDly3_bits"};
      this.Prbs0GenTapDly3.configure(this, null, "");
      this.Prbs0GenTapDly3.build();
      this.default_map.add_reg(this.Prbs0GenTapDly3, `UVM_REG_ADDR_WIDTH'h15, "RW", 0);
		this.Prbs0GenTapDly3_Prbs0GenTapDly3 = this.Prbs0GenTapDly3.Prbs0GenTapDly3;
      this.Prbs0GenTapDly4 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly4::type_id::create("Prbs0GenTapDly4",,get_full_name());
      if(this.Prbs0GenTapDly4.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenTapDly4.cg_bits.option.name = {get_name(), ".", "Prbs0GenTapDly4_bits"};
      this.Prbs0GenTapDly4.configure(this, null, "");
      this.Prbs0GenTapDly4.build();
      this.default_map.add_reg(this.Prbs0GenTapDly4, `UVM_REG_ADDR_WIDTH'h16, "RW", 0);
		this.Prbs0GenTapDly4_Prbs0GenTapDly4 = this.Prbs0GenTapDly4.Prbs0GenTapDly4;
      this.Prbs0GenTapDly5 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly5::type_id::create("Prbs0GenTapDly5",,get_full_name());
      if(this.Prbs0GenTapDly5.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenTapDly5.cg_bits.option.name = {get_name(), ".", "Prbs0GenTapDly5_bits"};
      this.Prbs0GenTapDly5.configure(this, null, "");
      this.Prbs0GenTapDly5.build();
      this.default_map.add_reg(this.Prbs0GenTapDly5, `UVM_REG_ADDR_WIDTH'h17, "RW", 0);
		this.Prbs0GenTapDly5_Prbs0GenTapDly5 = this.Prbs0GenTapDly5.Prbs0GenTapDly5;
      this.Prbs0GenTapDly6 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly6::type_id::create("Prbs0GenTapDly6",,get_full_name());
      if(this.Prbs0GenTapDly6.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenTapDly6.cg_bits.option.name = {get_name(), ".", "Prbs0GenTapDly6_bits"};
      this.Prbs0GenTapDly6.configure(this, null, "");
      this.Prbs0GenTapDly6.build();
      this.default_map.add_reg(this.Prbs0GenTapDly6, `UVM_REG_ADDR_WIDTH'h18, "RW", 0);
		this.Prbs0GenTapDly6_Prbs0GenTapDly6 = this.Prbs0GenTapDly6.Prbs0GenTapDly6;
      this.Prbs0GenTapDly7 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenTapDly7::type_id::create("Prbs0GenTapDly7",,get_full_name());
      if(this.Prbs0GenTapDly7.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenTapDly7.cg_bits.option.name = {get_name(), ".", "Prbs0GenTapDly7_bits"};
      this.Prbs0GenTapDly7.configure(this, null, "");
      this.Prbs0GenTapDly7.build();
      this.default_map.add_reg(this.Prbs0GenTapDly7, `UVM_REG_ADDR_WIDTH'h19, "RW", 0);
		this.Prbs0GenTapDly7_Prbs0GenTapDly7 = this.Prbs0GenTapDly7.Prbs0GenTapDly7;
      this.MtestMuxSel = ral_reg_DWC_DDRPHYA_PPGC0_p0_MtestMuxSel::type_id::create("MtestMuxSel",,get_full_name());
      if(this.MtestMuxSel.has_coverage(UVM_CVR_ALL))
      	this.MtestMuxSel.cg_bits.option.name = {get_name(), ".", "MtestMuxSel_bits"};
      this.MtestMuxSel.configure(this, null, "");
      this.MtestMuxSel.build();
      this.default_map.add_reg(this.MtestMuxSel, `UVM_REG_ADDR_WIDTH'h1A, "RW", 0);
		this.MtestMuxSel_MtestMuxSel = this.MtestMuxSel.MtestMuxSel;
      this.Prbs0GenStateLo = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateLo::type_id::create("Prbs0GenStateLo",,get_full_name());
      if(this.Prbs0GenStateLo.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenStateLo.cg_bits.option.name = {get_name(), ".", "Prbs0GenStateLo_bits"};
      this.Prbs0GenStateLo.configure(this, null, "");
      this.Prbs0GenStateLo.build();
      this.default_map.add_reg(this.Prbs0GenStateLo, `UVM_REG_ADDR_WIDTH'h1B, "RW", 0);
		this.Prbs0GenStateLo_Prbs0GenStateLo = this.Prbs0GenStateLo.Prbs0GenStateLo;
      this.Prbs0GenStateHi = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs0GenStateHi::type_id::create("Prbs0GenStateHi",,get_full_name());
      if(this.Prbs0GenStateHi.has_coverage(UVM_CVR_ALL))
      	this.Prbs0GenStateHi.cg_bits.option.name = {get_name(), ".", "Prbs0GenStateHi_bits"};
      this.Prbs0GenStateHi.configure(this, null, "");
      this.Prbs0GenStateHi.build();
      this.default_map.add_reg(this.Prbs0GenStateHi, `UVM_REG_ADDR_WIDTH'h1C, "RW", 0);
		this.Prbs0GenStateHi_Prbs0GenStateHi = this.Prbs0GenStateHi.Prbs0GenStateHi;
      this.Prbs1GenModeSel = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenModeSel::type_id::create("Prbs1GenModeSel",,get_full_name());
      if(this.Prbs1GenModeSel.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenModeSel.cg_bits.option.name = {get_name(), ".", "Prbs1GenModeSel_bits"};
      this.Prbs1GenModeSel.configure(this, null, "");
      this.Prbs1GenModeSel.build();
      this.default_map.add_reg(this.Prbs1GenModeSel, `UVM_REG_ADDR_WIDTH'h20, "RW", 0);
		this.Prbs1GenModeSel_Prbs1GenModeSel = this.Prbs1GenModeSel.Prbs1GenModeSel;
      this.Prbs1GenUiMuxSel = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenUiMuxSel::type_id::create("Prbs1GenUiMuxSel",,get_full_name());
      if(this.Prbs1GenUiMuxSel.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenUiMuxSel.cg_bits.option.name = {get_name(), ".", "Prbs1GenUiMuxSel_bits"};
      this.Prbs1GenUiMuxSel.configure(this, null, "");
      this.Prbs1GenUiMuxSel.build();
      this.default_map.add_reg(this.Prbs1GenUiMuxSel, `UVM_REG_ADDR_WIDTH'h21, "RW", 0);
		this.Prbs1GenUiMuxSel_Prbs1GenUiMuxSel = this.Prbs1GenUiMuxSel.Prbs1GenUiMuxSel;
      this.Prbs1GenTapDly0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly0::type_id::create("Prbs1GenTapDly0",,get_full_name());
      if(this.Prbs1GenTapDly0.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenTapDly0.cg_bits.option.name = {get_name(), ".", "Prbs1GenTapDly0_bits"};
      this.Prbs1GenTapDly0.configure(this, null, "");
      this.Prbs1GenTapDly0.build();
      this.default_map.add_reg(this.Prbs1GenTapDly0, `UVM_REG_ADDR_WIDTH'h22, "RW", 0);
		this.Prbs1GenTapDly0_Prbs1GenTapDly0 = this.Prbs1GenTapDly0.Prbs1GenTapDly0;
      this.Prbs1GenTapDly1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly1::type_id::create("Prbs1GenTapDly1",,get_full_name());
      if(this.Prbs1GenTapDly1.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenTapDly1.cg_bits.option.name = {get_name(), ".", "Prbs1GenTapDly1_bits"};
      this.Prbs1GenTapDly1.configure(this, null, "");
      this.Prbs1GenTapDly1.build();
      this.default_map.add_reg(this.Prbs1GenTapDly1, `UVM_REG_ADDR_WIDTH'h23, "RW", 0);
		this.Prbs1GenTapDly1_Prbs1GenTapDly1 = this.Prbs1GenTapDly1.Prbs1GenTapDly1;
      this.Prbs1GenTapDly2 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly2::type_id::create("Prbs1GenTapDly2",,get_full_name());
      if(this.Prbs1GenTapDly2.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenTapDly2.cg_bits.option.name = {get_name(), ".", "Prbs1GenTapDly2_bits"};
      this.Prbs1GenTapDly2.configure(this, null, "");
      this.Prbs1GenTapDly2.build();
      this.default_map.add_reg(this.Prbs1GenTapDly2, `UVM_REG_ADDR_WIDTH'h24, "RW", 0);
		this.Prbs1GenTapDly2_Prbs1GenTapDly2 = this.Prbs1GenTapDly2.Prbs1GenTapDly2;
      this.Prbs1GenTapDly3 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly3::type_id::create("Prbs1GenTapDly3",,get_full_name());
      if(this.Prbs1GenTapDly3.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenTapDly3.cg_bits.option.name = {get_name(), ".", "Prbs1GenTapDly3_bits"};
      this.Prbs1GenTapDly3.configure(this, null, "");
      this.Prbs1GenTapDly3.build();
      this.default_map.add_reg(this.Prbs1GenTapDly3, `UVM_REG_ADDR_WIDTH'h25, "RW", 0);
		this.Prbs1GenTapDly3_Prbs1GenTapDly3 = this.Prbs1GenTapDly3.Prbs1GenTapDly3;
      this.Prbs1GenTapDly4 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly4::type_id::create("Prbs1GenTapDly4",,get_full_name());
      if(this.Prbs1GenTapDly4.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenTapDly4.cg_bits.option.name = {get_name(), ".", "Prbs1GenTapDly4_bits"};
      this.Prbs1GenTapDly4.configure(this, null, "");
      this.Prbs1GenTapDly4.build();
      this.default_map.add_reg(this.Prbs1GenTapDly4, `UVM_REG_ADDR_WIDTH'h26, "RW", 0);
		this.Prbs1GenTapDly4_Prbs1GenTapDly4 = this.Prbs1GenTapDly4.Prbs1GenTapDly4;
      this.Prbs1GenTapDly5 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly5::type_id::create("Prbs1GenTapDly5",,get_full_name());
      if(this.Prbs1GenTapDly5.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenTapDly5.cg_bits.option.name = {get_name(), ".", "Prbs1GenTapDly5_bits"};
      this.Prbs1GenTapDly5.configure(this, null, "");
      this.Prbs1GenTapDly5.build();
      this.default_map.add_reg(this.Prbs1GenTapDly5, `UVM_REG_ADDR_WIDTH'h27, "RW", 0);
		this.Prbs1GenTapDly5_Prbs1GenTapDly5 = this.Prbs1GenTapDly5.Prbs1GenTapDly5;
      this.Prbs1GenTapDly6 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly6::type_id::create("Prbs1GenTapDly6",,get_full_name());
      if(this.Prbs1GenTapDly6.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenTapDly6.cg_bits.option.name = {get_name(), ".", "Prbs1GenTapDly6_bits"};
      this.Prbs1GenTapDly6.configure(this, null, "");
      this.Prbs1GenTapDly6.build();
      this.default_map.add_reg(this.Prbs1GenTapDly6, `UVM_REG_ADDR_WIDTH'h28, "RW", 0);
		this.Prbs1GenTapDly6_Prbs1GenTapDly6 = this.Prbs1GenTapDly6.Prbs1GenTapDly6;
      this.Prbs1GenTapDly7 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenTapDly7::type_id::create("Prbs1GenTapDly7",,get_full_name());
      if(this.Prbs1GenTapDly7.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenTapDly7.cg_bits.option.name = {get_name(), ".", "Prbs1GenTapDly7_bits"};
      this.Prbs1GenTapDly7.configure(this, null, "");
      this.Prbs1GenTapDly7.build();
      this.default_map.add_reg(this.Prbs1GenTapDly7, `UVM_REG_ADDR_WIDTH'h29, "RW", 0);
		this.Prbs1GenTapDly7_Prbs1GenTapDly7 = this.Prbs1GenTapDly7.Prbs1GenTapDly7;
      this.Prbs1GenStateLo = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateLo::type_id::create("Prbs1GenStateLo",,get_full_name());
      if(this.Prbs1GenStateLo.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenStateLo.cg_bits.option.name = {get_name(), ".", "Prbs1GenStateLo_bits"};
      this.Prbs1GenStateLo.configure(this, null, "");
      this.Prbs1GenStateLo.build();
      this.default_map.add_reg(this.Prbs1GenStateLo, `UVM_REG_ADDR_WIDTH'h2B, "RW", 0);
		this.Prbs1GenStateLo_Prbs1GenStateLo = this.Prbs1GenStateLo.Prbs1GenStateLo;
      this.Prbs1GenStateHi = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs1GenStateHi::type_id::create("Prbs1GenStateHi",,get_full_name());
      if(this.Prbs1GenStateHi.has_coverage(UVM_CVR_ALL))
      	this.Prbs1GenStateHi.cg_bits.option.name = {get_name(), ".", "Prbs1GenStateHi_bits"};
      this.Prbs1GenStateHi.configure(this, null, "");
      this.Prbs1GenStateHi.build();
      this.default_map.add_reg(this.Prbs1GenStateHi, `UVM_REG_ADDR_WIDTH'h2C, "RW", 0);
		this.Prbs1GenStateHi_Prbs1GenStateHi = this.Prbs1GenStateHi.Prbs1GenStateHi;
      this.Prbs2GenModeSel = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenModeSel::type_id::create("Prbs2GenModeSel",,get_full_name());
      if(this.Prbs2GenModeSel.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenModeSel.cg_bits.option.name = {get_name(), ".", "Prbs2GenModeSel_bits"};
      this.Prbs2GenModeSel.configure(this, null, "");
      this.Prbs2GenModeSel.build();
      this.default_map.add_reg(this.Prbs2GenModeSel, `UVM_REG_ADDR_WIDTH'h30, "RW", 0);
		this.Prbs2GenModeSel_Prbs2GenModeSel = this.Prbs2GenModeSel.Prbs2GenModeSel;
      this.Prbs2GenUiMuxSel = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenUiMuxSel::type_id::create("Prbs2GenUiMuxSel",,get_full_name());
      if(this.Prbs2GenUiMuxSel.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenUiMuxSel.cg_bits.option.name = {get_name(), ".", "Prbs2GenUiMuxSel_bits"};
      this.Prbs2GenUiMuxSel.configure(this, null, "");
      this.Prbs2GenUiMuxSel.build();
      this.default_map.add_reg(this.Prbs2GenUiMuxSel, `UVM_REG_ADDR_WIDTH'h31, "RW", 0);
		this.Prbs2GenUiMuxSel_Prbs2GenUiMuxSel = this.Prbs2GenUiMuxSel.Prbs2GenUiMuxSel;
      this.Prbs2GenTapDly0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly0::type_id::create("Prbs2GenTapDly0",,get_full_name());
      if(this.Prbs2GenTapDly0.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenTapDly0.cg_bits.option.name = {get_name(), ".", "Prbs2GenTapDly0_bits"};
      this.Prbs2GenTapDly0.configure(this, null, "");
      this.Prbs2GenTapDly0.build();
      this.default_map.add_reg(this.Prbs2GenTapDly0, `UVM_REG_ADDR_WIDTH'h32, "RW", 0);
		this.Prbs2GenTapDly0_Prbs2GenTapDly0 = this.Prbs2GenTapDly0.Prbs2GenTapDly0;
      this.Prbs2GenTapDly1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly1::type_id::create("Prbs2GenTapDly1",,get_full_name());
      if(this.Prbs2GenTapDly1.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenTapDly1.cg_bits.option.name = {get_name(), ".", "Prbs2GenTapDly1_bits"};
      this.Prbs2GenTapDly1.configure(this, null, "");
      this.Prbs2GenTapDly1.build();
      this.default_map.add_reg(this.Prbs2GenTapDly1, `UVM_REG_ADDR_WIDTH'h33, "RW", 0);
		this.Prbs2GenTapDly1_Prbs2GenTapDly1 = this.Prbs2GenTapDly1.Prbs2GenTapDly1;
      this.Prbs2GenTapDly2 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly2::type_id::create("Prbs2GenTapDly2",,get_full_name());
      if(this.Prbs2GenTapDly2.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenTapDly2.cg_bits.option.name = {get_name(), ".", "Prbs2GenTapDly2_bits"};
      this.Prbs2GenTapDly2.configure(this, null, "");
      this.Prbs2GenTapDly2.build();
      this.default_map.add_reg(this.Prbs2GenTapDly2, `UVM_REG_ADDR_WIDTH'h34, "RW", 0);
		this.Prbs2GenTapDly2_Prbs2GenTapDly2 = this.Prbs2GenTapDly2.Prbs2GenTapDly2;
      this.Prbs2GenTapDly3 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly3::type_id::create("Prbs2GenTapDly3",,get_full_name());
      if(this.Prbs2GenTapDly3.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenTapDly3.cg_bits.option.name = {get_name(), ".", "Prbs2GenTapDly3_bits"};
      this.Prbs2GenTapDly3.configure(this, null, "");
      this.Prbs2GenTapDly3.build();
      this.default_map.add_reg(this.Prbs2GenTapDly3, `UVM_REG_ADDR_WIDTH'h35, "RW", 0);
		this.Prbs2GenTapDly3_Prbs2GenTapDly3 = this.Prbs2GenTapDly3.Prbs2GenTapDly3;
      this.Prbs2GenTapDly4 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly4::type_id::create("Prbs2GenTapDly4",,get_full_name());
      if(this.Prbs2GenTapDly4.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenTapDly4.cg_bits.option.name = {get_name(), ".", "Prbs2GenTapDly4_bits"};
      this.Prbs2GenTapDly4.configure(this, null, "");
      this.Prbs2GenTapDly4.build();
      this.default_map.add_reg(this.Prbs2GenTapDly4, `UVM_REG_ADDR_WIDTH'h36, "RW", 0);
		this.Prbs2GenTapDly4_Prbs2GenTapDly4 = this.Prbs2GenTapDly4.Prbs2GenTapDly4;
      this.Prbs2GenTapDly5 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly5::type_id::create("Prbs2GenTapDly5",,get_full_name());
      if(this.Prbs2GenTapDly5.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenTapDly5.cg_bits.option.name = {get_name(), ".", "Prbs2GenTapDly5_bits"};
      this.Prbs2GenTapDly5.configure(this, null, "");
      this.Prbs2GenTapDly5.build();
      this.default_map.add_reg(this.Prbs2GenTapDly5, `UVM_REG_ADDR_WIDTH'h37, "RW", 0);
		this.Prbs2GenTapDly5_Prbs2GenTapDly5 = this.Prbs2GenTapDly5.Prbs2GenTapDly5;
      this.Prbs2GenTapDly6 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly6::type_id::create("Prbs2GenTapDly6",,get_full_name());
      if(this.Prbs2GenTapDly6.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenTapDly6.cg_bits.option.name = {get_name(), ".", "Prbs2GenTapDly6_bits"};
      this.Prbs2GenTapDly6.configure(this, null, "");
      this.Prbs2GenTapDly6.build();
      this.default_map.add_reg(this.Prbs2GenTapDly6, `UVM_REG_ADDR_WIDTH'h38, "RW", 0);
		this.Prbs2GenTapDly6_Prbs2GenTapDly6 = this.Prbs2GenTapDly6.Prbs2GenTapDly6;
      this.Prbs2GenTapDly7 = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenTapDly7::type_id::create("Prbs2GenTapDly7",,get_full_name());
      if(this.Prbs2GenTapDly7.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenTapDly7.cg_bits.option.name = {get_name(), ".", "Prbs2GenTapDly7_bits"};
      this.Prbs2GenTapDly7.configure(this, null, "");
      this.Prbs2GenTapDly7.build();
      this.default_map.add_reg(this.Prbs2GenTapDly7, `UVM_REG_ADDR_WIDTH'h39, "RW", 0);
		this.Prbs2GenTapDly7_Prbs2GenTapDly7 = this.Prbs2GenTapDly7.Prbs2GenTapDly7;
      this.Prbs2GenStateLo = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateLo::type_id::create("Prbs2GenStateLo",,get_full_name());
      if(this.Prbs2GenStateLo.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenStateLo.cg_bits.option.name = {get_name(), ".", "Prbs2GenStateLo_bits"};
      this.Prbs2GenStateLo.configure(this, null, "");
      this.Prbs2GenStateLo.build();
      this.default_map.add_reg(this.Prbs2GenStateLo, `UVM_REG_ADDR_WIDTH'h3B, "RW", 0);
		this.Prbs2GenStateLo_Prbs2GenStateLo = this.Prbs2GenStateLo.Prbs2GenStateLo;
      this.Prbs2GenStateHi = ral_reg_DWC_DDRPHYA_PPGC0_p0_Prbs2GenStateHi::type_id::create("Prbs2GenStateHi",,get_full_name());
      if(this.Prbs2GenStateHi.has_coverage(UVM_CVR_ALL))
      	this.Prbs2GenStateHi.cg_bits.option.name = {get_name(), ".", "Prbs2GenStateHi_bits"};
      this.Prbs2GenStateHi.configure(this, null, "");
      this.Prbs2GenStateHi.build();
      this.default_map.add_reg(this.Prbs2GenStateHi, `UVM_REG_ADDR_WIDTH'h3C, "RW", 0);
		this.Prbs2GenStateHi_Prbs2GenStateHi = this.Prbs2GenStateHi.Prbs2GenStateHi;
      this.PPTTrainSetup_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_PPTTrainSetup_p0::type_id::create("PPTTrainSetup_p0",,get_full_name());
      if(this.PPTTrainSetup_p0.has_coverage(UVM_CVR_ALL))
      	this.PPTTrainSetup_p0.cg_bits.option.name = {get_name(), ".", "PPTTrainSetup_p0_bits"};
      this.PPTTrainSetup_p0.configure(this, null, "");
      this.PPTTrainSetup_p0.build();
      this.default_map.add_reg(this.PPTTrainSetup_p0, `UVM_REG_ADDR_WIDTH'h40, "RW", 0);
		this.PPTTrainSetup_p0_PhyMstrTrainInterval = this.PPTTrainSetup_p0.PhyMstrTrainInterval;
		this.PhyMstrTrainInterval = this.PPTTrainSetup_p0.PhyMstrTrainInterval;
		this.PPTTrainSetup_p0_PhyMstrMaxReqToAck = this.PPTTrainSetup_p0.PhyMstrMaxReqToAck;
		this.PhyMstrMaxReqToAck = this.PPTTrainSetup_p0.PhyMstrMaxReqToAck;
      this.PhyMstrFreqOverride_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyMstrFreqOverride_p0::type_id::create("PhyMstrFreqOverride_p0",,get_full_name());
      if(this.PhyMstrFreqOverride_p0.has_coverage(UVM_CVR_ALL))
      	this.PhyMstrFreqOverride_p0.cg_bits.option.name = {get_name(), ".", "PhyMstrFreqOverride_p0_bits"};
      this.PhyMstrFreqOverride_p0.configure(this, null, "");
      this.PhyMstrFreqOverride_p0.build();
      this.default_map.add_reg(this.PhyMstrFreqOverride_p0, `UVM_REG_ADDR_WIDTH'h41, "RW", 0);
		this.PhyMstrFreqOverride_p0_PhyMstrFreqOverride_p0 = this.PhyMstrFreqOverride_p0.PhyMstrFreqOverride_p0;
      this.DfiInitComplete = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiInitComplete::type_id::create("DfiInitComplete",,get_full_name());
      if(this.DfiInitComplete.has_coverage(UVM_CVR_ALL))
      	this.DfiInitComplete.cg_bits.option.name = {get_name(), ".", "DfiInitComplete_bits"};
      this.DfiInitComplete.configure(this, null, "");
      this.DfiInitComplete.build();
      this.default_map.add_reg(this.DfiInitComplete, `UVM_REG_ADDR_WIDTH'h49, "RW", 0);
		this.DfiInitComplete_DfiInitComplete = this.DfiInitComplete.DfiInitComplete;
      this.PPGCParityInvert = ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCParityInvert::type_id::create("PPGCParityInvert",,get_full_name());
      if(this.PPGCParityInvert.has_coverage(UVM_CVR_ALL))
      	this.PPGCParityInvert.cg_bits.option.name = {get_name(), ".", "PPGCParityInvert_bits"};
      this.PPGCParityInvert.configure(this, null, "");
      this.PPGCParityInvert.build();
      this.default_map.add_reg(this.PPGCParityInvert, `UVM_REG_ADDR_WIDTH'h4D, "RW", 0);
		this.PPGCParityInvert_PPGCParityInvert = this.PPGCParityInvert.PPGCParityInvert;
      this.PMIEnable = ral_reg_DWC_DDRPHYA_PPGC0_p0_PMIEnable::type_id::create("PMIEnable",,get_full_name());
      if(this.PMIEnable.has_coverage(UVM_CVR_ALL))
      	this.PMIEnable.cg_bits.option.name = {get_name(), ".", "PMIEnable_bits"};
      this.PMIEnable.configure(this, null, "");
      this.PMIEnable.build();
      this.default_map.add_reg(this.PMIEnable, `UVM_REG_ADDR_WIDTH'h54, "RW", 0);
		this.PMIEnable_PMIEnable = this.PMIEnable.PMIEnable;
      this.Dfi0Status = ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi0Status::type_id::create("Dfi0Status",,get_full_name());
      if(this.Dfi0Status.has_coverage(UVM_CVR_ALL))
      	this.Dfi0Status.cg_bits.option.name = {get_name(), ".", "Dfi0Status_bits"};
      this.Dfi0Status.configure(this, null, "");
      this.Dfi0Status.build();
      this.default_map.add_reg(this.Dfi0Status, `UVM_REG_ADDR_WIDTH'h5A, "RO", 0);
		this.Dfi0Status_Dfi0Status = this.Dfi0Status.Dfi0Status;
      this.Dfi1Status = ral_reg_DWC_DDRPHYA_PPGC0_p0_Dfi1Status::type_id::create("Dfi1Status",,get_full_name());
      if(this.Dfi1Status.has_coverage(UVM_CVR_ALL))
      	this.Dfi1Status.cg_bits.option.name = {get_name(), ".", "Dfi1Status_bits"};
      this.Dfi1Status.configure(this, null, "");
      this.Dfi1Status.build();
      this.default_map.add_reg(this.Dfi1Status, `UVM_REG_ADDR_WIDTH'h5B, "RO", 0);
		this.Dfi1Status_Dfi1Status = this.Dfi1Status.Dfi1Status;
      this.DfiHandshakeDelays0_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays0_p0::type_id::create("DfiHandshakeDelays0_p0",,get_full_name());
      if(this.DfiHandshakeDelays0_p0.has_coverage(UVM_CVR_ALL))
      	this.DfiHandshakeDelays0_p0.cg_bits.option.name = {get_name(), ".", "DfiHandshakeDelays0_p0_bits"};
      this.DfiHandshakeDelays0_p0.configure(this, null, "");
      this.DfiHandshakeDelays0_p0.build();
      this.default_map.add_reg(this.DfiHandshakeDelays0_p0, `UVM_REG_ADDR_WIDTH'h66, "RW", 0);
		this.DfiHandshakeDelays0_p0_PhyUpdAckDelay0 = this.DfiHandshakeDelays0_p0.PhyUpdAckDelay0;
		this.PhyUpdAckDelay0 = this.DfiHandshakeDelays0_p0.PhyUpdAckDelay0;
		this.DfiHandshakeDelays0_p0_PhyUpdReqDelay0 = this.DfiHandshakeDelays0_p0.PhyUpdReqDelay0;
		this.PhyUpdReqDelay0 = this.DfiHandshakeDelays0_p0.PhyUpdReqDelay0;
		this.DfiHandshakeDelays0_p0_CtrlUpdReqDelay0 = this.DfiHandshakeDelays0_p0.CtrlUpdReqDelay0;
		this.CtrlUpdReqDelay0 = this.DfiHandshakeDelays0_p0.CtrlUpdReqDelay0;
      this.DFIPHYUPD0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD0::type_id::create("DFIPHYUPD0",,get_full_name());
      if(this.DFIPHYUPD0.has_coverage(UVM_CVR_ALL))
      	this.DFIPHYUPD0.cg_bits.option.name = {get_name(), ".", "DFIPHYUPD0_bits"};
      this.DFIPHYUPD0.configure(this, null, "");
      this.DFIPHYUPD0.build();
      this.default_map.add_reg(this.DFIPHYUPD0, `UVM_REG_ADDR_WIDTH'h67, "RW", 0);
		this.DFIPHYUPD0_DFIPHYUPDCNT0 = this.DFIPHYUPD0.DFIPHYUPDCNT0;
		this.DFIPHYUPDCNT0 = this.DFIPHYUPD0.DFIPHYUPDCNT0;
		this.DFIPHYUPD0_DFIPHYUPDRESP0 = this.DFIPHYUPD0.DFIPHYUPDRESP0;
		this.DFIPHYUPDRESP0 = this.DFIPHYUPD0.DFIPHYUPDRESP0;
      this.DfiLpCtrlEn0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn0::type_id::create("DfiLpCtrlEn0",,get_full_name());
      if(this.DfiLpCtrlEn0.has_coverage(UVM_CVR_ALL))
      	this.DfiLpCtrlEn0.cg_bits.option.name = {get_name(), ".", "DfiLpCtrlEn0_bits"};
      this.DfiLpCtrlEn0.configure(this, null, "");
      this.DfiLpCtrlEn0.build();
      this.default_map.add_reg(this.DfiLpCtrlEn0, `UVM_REG_ADDR_WIDTH'h68, "RW", 0);
		this.DfiLpCtrlEn0_DfiLpCtrlEn0 = this.DfiLpCtrlEn0.DfiLpCtrlEn0;
      this.DfiLpDataEn0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn0::type_id::create("DfiLpDataEn0",,get_full_name());
      if(this.DfiLpDataEn0.has_coverage(UVM_CVR_ALL))
      	this.DfiLpDataEn0.cg_bits.option.name = {get_name(), ".", "DfiLpDataEn0_bits"};
      this.DfiLpDataEn0.configure(this, null, "");
      this.DfiLpDataEn0.build();
      this.default_map.add_reg(this.DfiLpDataEn0, `UVM_REG_ADDR_WIDTH'h69, "RW", 0);
		this.DfiLpDataEn0_DfiLpDataEn0 = this.DfiLpDataEn0.DfiLpDataEn0;
      this.DynOdtEnCntrl0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl0::type_id::create("DynOdtEnCntrl0",,get_full_name());
      if(this.DynOdtEnCntrl0.has_coverage(UVM_CVR_ALL))
      	this.DynOdtEnCntrl0.cg_bits.option.name = {get_name(), ".", "DynOdtEnCntrl0_bits"};
      this.DynOdtEnCntrl0.configure(this, null, "");
      this.DynOdtEnCntrl0.build();
      this.default_map.add_reg(this.DynOdtEnCntrl0, `UVM_REG_ADDR_WIDTH'h6A, "RW", 0);
		this.DynOdtEnCntrl0_DbyteDynOdtEn0 = this.DynOdtEnCntrl0.DbyteDynOdtEn0;
		this.DbyteDynOdtEn0 = this.DynOdtEnCntrl0.DbyteDynOdtEn0;
      this.DfiRespHandshakeDelays0_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays0_p0::type_id::create("DfiRespHandshakeDelays0_p0",,get_full_name());
      if(this.DfiRespHandshakeDelays0_p0.has_coverage(UVM_CVR_ALL))
      	this.DfiRespHandshakeDelays0_p0.cg_bits.option.name = {get_name(), ".", "DfiRespHandshakeDelays0_p0_bits"};
      this.DfiRespHandshakeDelays0_p0.configure(this, null, "");
      this.DfiRespHandshakeDelays0_p0.build();
      this.default_map.add_reg(this.DfiRespHandshakeDelays0_p0, `UVM_REG_ADDR_WIDTH'h6B, "RW", 0);
		this.DfiRespHandshakeDelays0_p0_LpCtrlAckDelay0 = this.DfiRespHandshakeDelays0_p0.LpCtrlAckDelay0;
		this.LpCtrlAckDelay0 = this.DfiRespHandshakeDelays0_p0.LpCtrlAckDelay0;
		this.DfiRespHandshakeDelays0_p0_LpDataAckDelay0 = this.DfiRespHandshakeDelays0_p0.LpDataAckDelay0;
		this.LpDataAckDelay0 = this.DfiRespHandshakeDelays0_p0.LpDataAckDelay0;
		this.DfiRespHandshakeDelays0_p0_CtrlUpdAckDelay0 = this.DfiRespHandshakeDelays0_p0.CtrlUpdAckDelay0;
		this.CtrlUpdAckDelay0 = this.DfiRespHandshakeDelays0_p0.CtrlUpdAckDelay0;
		this.DfiRespHandshakeDelays0_p0_LpAssertAckDelay0 = this.DfiRespHandshakeDelays0_p0.LpAssertAckDelay0;
		this.LpAssertAckDelay0 = this.DfiRespHandshakeDelays0_p0.LpAssertAckDelay0;
      this.HwtLpCsEnA = ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnA::type_id::create("HwtLpCsEnA",,get_full_name());
      if(this.HwtLpCsEnA.has_coverage(UVM_CVR_ALL))
      	this.HwtLpCsEnA.cg_bits.option.name = {get_name(), ".", "HwtLpCsEnA_bits"};
      this.HwtLpCsEnA.configure(this, null, "");
      this.HwtLpCsEnA.build();
      this.default_map.add_reg(this.HwtLpCsEnA, `UVM_REG_ADDR_WIDTH'h72, "RW", 0);
		this.HwtLpCsEnA_HwtLpCsEnA = this.HwtLpCsEnA.HwtLpCsEnA;
      this.HwtLpCsEnB = ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnB::type_id::create("HwtLpCsEnB",,get_full_name());
      if(this.HwtLpCsEnB.has_coverage(UVM_CVR_ALL))
      	this.HwtLpCsEnB.cg_bits.option.name = {get_name(), ".", "HwtLpCsEnB_bits"};
      this.HwtLpCsEnB.configure(this, null, "");
      this.HwtLpCsEnB.build();
      this.default_map.add_reg(this.HwtLpCsEnB, `UVM_REG_ADDR_WIDTH'h73, "RW", 0);
		this.HwtLpCsEnB_HwtLpCsEnB = this.HwtLpCsEnB.HwtLpCsEnB;
      this.HwtCtrl = ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtCtrl::type_id::create("HwtCtrl",,get_full_name());
      if(this.HwtCtrl.has_coverage(UVM_CVR_ALL))
      	this.HwtCtrl.cg_bits.option.name = {get_name(), ".", "HwtCtrl_bits"};
      this.HwtCtrl.configure(this, null, "");
      this.HwtCtrl.build();
      this.default_map.add_reg(this.HwtCtrl, `UVM_REG_ADDR_WIDTH'h77, "RW", 0);
		this.HwtCtrl_HwtCtrl = this.HwtCtrl.HwtCtrl;
      this.HwtControlOvr = ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlOvr::type_id::create("HwtControlOvr",,get_full_name());
      if(this.HwtControlOvr.has_coverage(UVM_CVR_ALL))
      	this.HwtControlOvr.cg_bits.option.name = {get_name(), ".", "HwtControlOvr_bits"};
      this.HwtControlOvr.configure(this, null, "");
      this.HwtControlOvr.build();
      this.default_map.add_reg(this.HwtControlOvr, `UVM_REG_ADDR_WIDTH'h7A, "RW", 0);
		this.HwtControlOvr_HwtControlOvr = this.HwtControlOvr.HwtControlOvr;
      this.ScratchPadPPGC = ral_reg_DWC_DDRPHYA_PPGC0_p0_ScratchPadPPGC::type_id::create("ScratchPadPPGC",,get_full_name());
      if(this.ScratchPadPPGC.has_coverage(UVM_CVR_ALL))
      	this.ScratchPadPPGC.cg_bits.option.name = {get_name(), ".", "ScratchPadPPGC_bits"};
      this.ScratchPadPPGC.configure(this, null, "");
      this.ScratchPadPPGC.build();
      this.default_map.add_reg(this.ScratchPadPPGC, `UVM_REG_ADDR_WIDTH'h7D, "RW", 0);
		this.ScratchPadPPGC_ScratchPadPPGC = this.ScratchPadPPGC.ScratchPadPPGC;
      this.HwtControlVal = ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtControlVal::type_id::create("HwtControlVal",,get_full_name());
      if(this.HwtControlVal.has_coverage(UVM_CVR_ALL))
      	this.HwtControlVal.cg_bits.option.name = {get_name(), ".", "HwtControlVal_bits"};
      this.HwtControlVal.configure(this, null, "");
      this.HwtControlVal.build();
      this.default_map.add_reg(this.HwtControlVal, `UVM_REG_ADDR_WIDTH'h7E, "RW", 0);
		this.HwtControlVal_HwtControlVal = this.HwtControlVal.HwtControlVal;
      this.ForceHWTClkGaterEnables = ral_reg_DWC_DDRPHYA_PPGC0_p0_ForceHWTClkGaterEnables::type_id::create("ForceHWTClkGaterEnables",,get_full_name());
      if(this.ForceHWTClkGaterEnables.has_coverage(UVM_CVR_ALL))
      	this.ForceHWTClkGaterEnables.cg_bits.option.name = {get_name(), ".", "ForceHWTClkGaterEnables_bits"};
      this.ForceHWTClkGaterEnables.configure(this, null, "");
      this.ForceHWTClkGaterEnables.build();
      this.default_map.add_reg(this.ForceHWTClkGaterEnables, `UVM_REG_ADDR_WIDTH'h80, "RW", 0);
		this.ForceHWTClkGaterEnables_ForceACSMClkEnHigh = this.ForceHWTClkGaterEnables.ForceACSMClkEnHigh;
		this.ForceACSMClkEnHigh = this.ForceHWTClkGaterEnables.ForceACSMClkEnHigh;
		this.ForceHWTClkGaterEnables_ForceACSMClkEnLow = this.ForceHWTClkGaterEnables.ForceACSMClkEnLow;
		this.ForceACSMClkEnLow = this.ForceHWTClkGaterEnables.ForceACSMClkEnLow;
		this.ForceHWTClkGaterEnables_ForcePIEClkEnHigh = this.ForceHWTClkGaterEnables.ForcePIEClkEnHigh;
		this.ForcePIEClkEnHigh = this.ForceHWTClkGaterEnables.ForcePIEClkEnHigh;
		this.ForceHWTClkGaterEnables_ForcePIEClkEnLow = this.ForceHWTClkGaterEnables.ForcePIEClkEnLow;
		this.ForcePIEClkEnLow = this.ForceHWTClkGaterEnables.ForcePIEClkEnLow;
      this.MasUpdGoodCtr = ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdGoodCtr::type_id::create("MasUpdGoodCtr",,get_full_name());
      if(this.MasUpdGoodCtr.has_coverage(UVM_CVR_ALL))
      	this.MasUpdGoodCtr.cg_bits.option.name = {get_name(), ".", "MasUpdGoodCtr_bits"};
      this.MasUpdGoodCtr.configure(this, null, "");
      this.MasUpdGoodCtr.build();
      this.default_map.add_reg(this.MasUpdGoodCtr, `UVM_REG_ADDR_WIDTH'hB5, "RO", 0);
		this.MasUpdGoodCtr_MasUpdGoodCtr = this.MasUpdGoodCtr.MasUpdGoodCtr;
      this.PhyUpd0GoodCtr = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0GoodCtr::type_id::create("PhyUpd0GoodCtr",,get_full_name());
      if(this.PhyUpd0GoodCtr.has_coverage(UVM_CVR_ALL))
      	this.PhyUpd0GoodCtr.cg_bits.option.name = {get_name(), ".", "PhyUpd0GoodCtr_bits"};
      this.PhyUpd0GoodCtr.configure(this, null, "");
      this.PhyUpd0GoodCtr.build();
      this.default_map.add_reg(this.PhyUpd0GoodCtr, `UVM_REG_ADDR_WIDTH'hB6, "RO", 0);
		this.PhyUpd0GoodCtr_PhyUpd0GoodCtr = this.PhyUpd0GoodCtr.PhyUpd0GoodCtr;
      this.PhyUpd1GoodCtr = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1GoodCtr::type_id::create("PhyUpd1GoodCtr",,get_full_name());
      if(this.PhyUpd1GoodCtr.has_coverage(UVM_CVR_ALL))
      	this.PhyUpd1GoodCtr.cg_bits.option.name = {get_name(), ".", "PhyUpd1GoodCtr_bits"};
      this.PhyUpd1GoodCtr.configure(this, null, "");
      this.PhyUpd1GoodCtr.build();
      this.default_map.add_reg(this.PhyUpd1GoodCtr, `UVM_REG_ADDR_WIDTH'hB7, "RO", 0);
		this.PhyUpd1GoodCtr_PhyUpd1GoodCtr = this.PhyUpd1GoodCtr.PhyUpd1GoodCtr;
      this.CtlUpd0GoodCtr = ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd0GoodCtr::type_id::create("CtlUpd0GoodCtr",,get_full_name());
      if(this.CtlUpd0GoodCtr.has_coverage(UVM_CVR_ALL))
      	this.CtlUpd0GoodCtr.cg_bits.option.name = {get_name(), ".", "CtlUpd0GoodCtr_bits"};
      this.CtlUpd0GoodCtr.configure(this, null, "");
      this.CtlUpd0GoodCtr.build();
      this.default_map.add_reg(this.CtlUpd0GoodCtr, `UVM_REG_ADDR_WIDTH'hB8, "RO", 0);
		this.CtlUpd0GoodCtr_CtlUpd0GoodCtr = this.CtlUpd0GoodCtr.CtlUpd0GoodCtr;
      this.CtlUpd1GoodCtr = ral_reg_DWC_DDRPHYA_PPGC0_p0_CtlUpd1GoodCtr::type_id::create("CtlUpd1GoodCtr",,get_full_name());
      if(this.CtlUpd1GoodCtr.has_coverage(UVM_CVR_ALL))
      	this.CtlUpd1GoodCtr.cg_bits.option.name = {get_name(), ".", "CtlUpd1GoodCtr_bits"};
      this.CtlUpd1GoodCtr.configure(this, null, "");
      this.CtlUpd1GoodCtr.build();
      this.default_map.add_reg(this.CtlUpd1GoodCtr, `UVM_REG_ADDR_WIDTH'hB9, "RO", 0);
		this.CtlUpd1GoodCtr_CtlUpd1GoodCtr = this.CtlUpd1GoodCtr.CtlUpd1GoodCtr;
      this.MasUpdFailCtr = ral_reg_DWC_DDRPHYA_PPGC0_p0_MasUpdFailCtr::type_id::create("MasUpdFailCtr",,get_full_name());
      if(this.MasUpdFailCtr.has_coverage(UVM_CVR_ALL))
      	this.MasUpdFailCtr.cg_bits.option.name = {get_name(), ".", "MasUpdFailCtr_bits"};
      this.MasUpdFailCtr.configure(this, null, "");
      this.MasUpdFailCtr.build();
      this.default_map.add_reg(this.MasUpdFailCtr, `UVM_REG_ADDR_WIDTH'hBA, "RO", 0);
		this.MasUpdFailCtr_MasUpdFailCtr = this.MasUpdFailCtr.MasUpdFailCtr;
      this.PhyUpd0FailCtr = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd0FailCtr::type_id::create("PhyUpd0FailCtr",,get_full_name());
      if(this.PhyUpd0FailCtr.has_coverage(UVM_CVR_ALL))
      	this.PhyUpd0FailCtr.cg_bits.option.name = {get_name(), ".", "PhyUpd0FailCtr_bits"};
      this.PhyUpd0FailCtr.configure(this, null, "");
      this.PhyUpd0FailCtr.build();
      this.default_map.add_reg(this.PhyUpd0FailCtr, `UVM_REG_ADDR_WIDTH'hBB, "RO", 0);
		this.PhyUpd0FailCtr_PhyUpd0FailCtr = this.PhyUpd0FailCtr.PhyUpd0FailCtr;
      this.PhyUpd1FailCtr = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyUpd1FailCtr::type_id::create("PhyUpd1FailCtr",,get_full_name());
      if(this.PhyUpd1FailCtr.has_coverage(UVM_CVR_ALL))
      	this.PhyUpd1FailCtr.cg_bits.option.name = {get_name(), ".", "PhyUpd1FailCtr_bits"};
      this.PhyUpd1FailCtr.configure(this, null, "");
      this.PhyUpd1FailCtr.build();
      this.default_map.add_reg(this.PhyUpd1FailCtr, `UVM_REG_ADDR_WIDTH'hBC, "RO", 0);
		this.PhyUpd1FailCtr_PhyUpd1FailCtr = this.PhyUpd1FailCtr.PhyUpd1FailCtr;
      this.PhyPerfCtrEnable = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyPerfCtrEnable::type_id::create("PhyPerfCtrEnable",,get_full_name());
      if(this.PhyPerfCtrEnable.has_coverage(UVM_CVR_ALL))
      	this.PhyPerfCtrEnable.cg_bits.option.name = {get_name(), ".", "PhyPerfCtrEnable_bits"};
      this.PhyPerfCtrEnable.configure(this, null, "");
      this.PhyPerfCtrEnable.build();
      this.default_map.add_reg(this.PhyPerfCtrEnable, `UVM_REG_ADDR_WIDTH'hBD, "RW", 0);
		this.PhyPerfCtrEnable_MasUpdGoodCtl = this.PhyPerfCtrEnable.MasUpdGoodCtl;
		this.MasUpdGoodCtl = this.PhyPerfCtrEnable.MasUpdGoodCtl;
		this.PhyPerfCtrEnable_PhyUpd0GoodCtl = this.PhyPerfCtrEnable.PhyUpd0GoodCtl;
		this.PhyUpd0GoodCtl = this.PhyPerfCtrEnable.PhyUpd0GoodCtl;
		this.PhyPerfCtrEnable_PhyUpd1GoodCtl = this.PhyPerfCtrEnable.PhyUpd1GoodCtl;
		this.PhyUpd1GoodCtl = this.PhyPerfCtrEnable.PhyUpd1GoodCtl;
		this.PhyPerfCtrEnable_CtlUpd0GoodCtl = this.PhyPerfCtrEnable.CtlUpd0GoodCtl;
		this.CtlUpd0GoodCtl = this.PhyPerfCtrEnable.CtlUpd0GoodCtl;
		this.PhyPerfCtrEnable_CtlUpd1GoodCtl = this.PhyPerfCtrEnable.CtlUpd1GoodCtl;
		this.CtlUpd1GoodCtl = this.PhyPerfCtrEnable.CtlUpd1GoodCtl;
		this.PhyPerfCtrEnable_MasUpdFailCtl = this.PhyPerfCtrEnable.MasUpdFailCtl;
		this.MasUpdFailCtl = this.PhyPerfCtrEnable.MasUpdFailCtl;
		this.PhyPerfCtrEnable_PhyUpd0FailCtl = this.PhyPerfCtrEnable.PhyUpd0FailCtl;
		this.PhyUpd0FailCtl = this.PhyPerfCtrEnable.PhyUpd0FailCtl;
		this.PhyPerfCtrEnable_PhyUpd1FailCtl = this.PhyPerfCtrEnable.PhyUpd1FailCtl;
		this.PhyUpd1FailCtl = this.PhyPerfCtrEnable.PhyUpd1FailCtl;
      this.DfiHandshakeDelays1_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiHandshakeDelays1_p0::type_id::create("DfiHandshakeDelays1_p0",,get_full_name());
      if(this.DfiHandshakeDelays1_p0.has_coverage(UVM_CVR_ALL))
      	this.DfiHandshakeDelays1_p0.cg_bits.option.name = {get_name(), ".", "DfiHandshakeDelays1_p0_bits"};
      this.DfiHandshakeDelays1_p0.configure(this, null, "");
      this.DfiHandshakeDelays1_p0.build();
      this.default_map.add_reg(this.DfiHandshakeDelays1_p0, `UVM_REG_ADDR_WIDTH'hE6, "RW", 0);
		this.DfiHandshakeDelays1_p0_PhyUpdAckDelay1 = this.DfiHandshakeDelays1_p0.PhyUpdAckDelay1;
		this.PhyUpdAckDelay1 = this.DfiHandshakeDelays1_p0.PhyUpdAckDelay1;
		this.DfiHandshakeDelays1_p0_PhyUpdReqDelay1 = this.DfiHandshakeDelays1_p0.PhyUpdReqDelay1;
		this.PhyUpdReqDelay1 = this.DfiHandshakeDelays1_p0.PhyUpdReqDelay1;
		this.DfiHandshakeDelays1_p0_CtrlUpdReqDelay1 = this.DfiHandshakeDelays1_p0.CtrlUpdReqDelay1;
		this.CtrlUpdReqDelay1 = this.DfiHandshakeDelays1_p0.CtrlUpdReqDelay1;
      this.DFIPHYUPD1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DFIPHYUPD1::type_id::create("DFIPHYUPD1",,get_full_name());
      if(this.DFIPHYUPD1.has_coverage(UVM_CVR_ALL))
      	this.DFIPHYUPD1.cg_bits.option.name = {get_name(), ".", "DFIPHYUPD1_bits"};
      this.DFIPHYUPD1.configure(this, null, "");
      this.DFIPHYUPD1.build();
      this.default_map.add_reg(this.DFIPHYUPD1, `UVM_REG_ADDR_WIDTH'hE7, "RW", 0);
		this.DFIPHYUPD1_DFIPHYUPDCNT1 = this.DFIPHYUPD1.DFIPHYUPDCNT1;
		this.DFIPHYUPDCNT1 = this.DFIPHYUPD1.DFIPHYUPDCNT1;
		this.DFIPHYUPD1_DFIPHYUPDRESP1 = this.DFIPHYUPD1.DFIPHYUPDRESP1;
		this.DFIPHYUPDRESP1 = this.DFIPHYUPD1.DFIPHYUPDRESP1;
      this.DfiLpCtrlEn1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpCtrlEn1::type_id::create("DfiLpCtrlEn1",,get_full_name());
      if(this.DfiLpCtrlEn1.has_coverage(UVM_CVR_ALL))
      	this.DfiLpCtrlEn1.cg_bits.option.name = {get_name(), ".", "DfiLpCtrlEn1_bits"};
      this.DfiLpCtrlEn1.configure(this, null, "");
      this.DfiLpCtrlEn1.build();
      this.default_map.add_reg(this.DfiLpCtrlEn1, `UVM_REG_ADDR_WIDTH'hE8, "RW", 0);
		this.DfiLpCtrlEn1_DfiLpCtrlEn1 = this.DfiLpCtrlEn1.DfiLpCtrlEn1;
      this.DfiLpDataEn1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiLpDataEn1::type_id::create("DfiLpDataEn1",,get_full_name());
      if(this.DfiLpDataEn1.has_coverage(UVM_CVR_ALL))
      	this.DfiLpDataEn1.cg_bits.option.name = {get_name(), ".", "DfiLpDataEn1_bits"};
      this.DfiLpDataEn1.configure(this, null, "");
      this.DfiLpDataEn1.build();
      this.default_map.add_reg(this.DfiLpDataEn1, `UVM_REG_ADDR_WIDTH'hE9, "RW", 0);
		this.DfiLpDataEn1_DfiLpDataEn1 = this.DfiLpDataEn1.DfiLpDataEn1;
      this.DynOdtEnCntrl1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DynOdtEnCntrl1::type_id::create("DynOdtEnCntrl1",,get_full_name());
      if(this.DynOdtEnCntrl1.has_coverage(UVM_CVR_ALL))
      	this.DynOdtEnCntrl1.cg_bits.option.name = {get_name(), ".", "DynOdtEnCntrl1_bits"};
      this.DynOdtEnCntrl1.configure(this, null, "");
      this.DynOdtEnCntrl1.build();
      this.default_map.add_reg(this.DynOdtEnCntrl1, `UVM_REG_ADDR_WIDTH'hEA, "RW", 0);
		this.DynOdtEnCntrl1_DbyteDynOdtEn1 = this.DynOdtEnCntrl1.DbyteDynOdtEn1;
		this.DbyteDynOdtEn1 = this.DynOdtEnCntrl1.DbyteDynOdtEn1;
      this.DfiRespHandshakeDelays1_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_DfiRespHandshakeDelays1_p0::type_id::create("DfiRespHandshakeDelays1_p0",,get_full_name());
      if(this.DfiRespHandshakeDelays1_p0.has_coverage(UVM_CVR_ALL))
      	this.DfiRespHandshakeDelays1_p0.cg_bits.option.name = {get_name(), ".", "DfiRespHandshakeDelays1_p0_bits"};
      this.DfiRespHandshakeDelays1_p0.configure(this, null, "");
      this.DfiRespHandshakeDelays1_p0.build();
      this.default_map.add_reg(this.DfiRespHandshakeDelays1_p0, `UVM_REG_ADDR_WIDTH'hEB, "RW", 0);
		this.DfiRespHandshakeDelays1_p0_LpCtrlAckDelay1 = this.DfiRespHandshakeDelays1_p0.LpCtrlAckDelay1;
		this.LpCtrlAckDelay1 = this.DfiRespHandshakeDelays1_p0.LpCtrlAckDelay1;
		this.DfiRespHandshakeDelays1_p0_LpDataAckDelay1 = this.DfiRespHandshakeDelays1_p0.LpDataAckDelay1;
		this.LpDataAckDelay1 = this.DfiRespHandshakeDelays1_p0.LpDataAckDelay1;
		this.DfiRespHandshakeDelays1_p0_CtrlUpdAckDelay1 = this.DfiRespHandshakeDelays1_p0.CtrlUpdAckDelay1;
		this.CtrlUpdAckDelay1 = this.DfiRespHandshakeDelays1_p0.CtrlUpdAckDelay1;
		this.DfiRespHandshakeDelays1_p0_LpAssertAckDelay1 = this.DfiRespHandshakeDelays1_p0.LpAssertAckDelay1;
		this.LpAssertAckDelay1 = this.DfiRespHandshakeDelays1_p0.LpAssertAckDelay1;
      this.FspSkipList = ral_reg_DWC_DDRPHYA_PPGC0_p0_FspSkipList::type_id::create("FspSkipList",,get_full_name());
      if(this.FspSkipList.has_coverage(UVM_CVR_ALL))
      	this.FspSkipList.cg_bits.option.name = {get_name(), ".", "FspSkipList_bits"};
      this.FspSkipList.configure(this, null, "");
      this.FspSkipList.build();
      this.default_map.add_reg(this.FspSkipList, `UVM_REG_ADDR_WIDTH'hF0, "RW", 0);
		this.FspSkipList_FspPStateSkip0 = this.FspSkipList.FspPStateSkip0;
		this.FspPStateSkip0 = this.FspSkipList.FspPStateSkip0;
		this.FspSkipList_FspPStateSkip1 = this.FspSkipList.FspPStateSkip1;
		this.FspPStateSkip1 = this.FspSkipList.FspPStateSkip1;
		this.FspSkipList_FspPStateSkip2 = this.FspSkipList.FspPStateSkip2;
		this.FspPStateSkip2 = this.FspSkipList.FspPStateSkip2;
		this.FspSkipList_FspPStateSkip3 = this.FspSkipList.FspPStateSkip3;
		this.FspPStateSkip3 = this.FspSkipList.FspPStateSkip3;
      this.PPGCReserved0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_PPGCReserved0::type_id::create("PPGCReserved0",,get_full_name());
      if(this.PPGCReserved0.has_coverage(UVM_CVR_ALL))
      	this.PPGCReserved0.cg_bits.option.name = {get_name(), ".", "PPGCReserved0_bits"};
      this.PPGCReserved0.configure(this, null, "");
      this.PPGCReserved0.build();
      this.default_map.add_reg(this.PPGCReserved0, `UVM_REG_ADDR_WIDTH'hFA, "RW", 0);
		this.PPGCReserved0_PPGCReserved0 = this.PPGCReserved0.PPGCReserved0;
      this.PUBReservedP1_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_PUBReservedP1_p0::type_id::create("PUBReservedP1_p0",,get_full_name());
      if(this.PUBReservedP1_p0.has_coverage(UVM_CVR_ALL))
      	this.PUBReservedP1_p0.cg_bits.option.name = {get_name(), ".", "PUBReservedP1_p0_bits"};
      this.PUBReservedP1_p0.configure(this, null, "");
      this.PUBReservedP1_p0.build();
      this.default_map.add_reg(this.PUBReservedP1_p0, `UVM_REG_ADDR_WIDTH'hFF, "RW", 0);
		this.PUBReservedP1_p0_PUBReservedP1_p0 = this.PUBReservedP1_p0.PUBReservedP1_p0;
      this.PhyInterruptOverride = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptOverride::type_id::create("PhyInterruptOverride",,get_full_name());
      if(this.PhyInterruptOverride.has_coverage(UVM_CVR_ALL))
      	this.PhyInterruptOverride.cg_bits.option.name = {get_name(), ".", "PhyInterruptOverride_bits"};
      this.PhyInterruptOverride.configure(this, null, "");
      this.PhyInterruptOverride.build();
      this.default_map.add_reg(this.PhyInterruptOverride, `UVM_REG_ADDR_WIDTH'h11A, "RW", 0);
		this.PhyInterruptOverride_PhyInterruptOverride = this.PhyInterruptOverride.PhyInterruptOverride;
      this.PhyInterruptEnable = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptEnable::type_id::create("PhyInterruptEnable",,get_full_name());
      if(this.PhyInterruptEnable.has_coverage(UVM_CVR_ALL))
      	this.PhyInterruptEnable.cg_bits.option.name = {get_name(), ".", "PhyInterruptEnable_bits"};
      this.PhyInterruptEnable.configure(this, null, "");
      this.PhyInterruptEnable.build();
      this.default_map.add_reg(this.PhyInterruptEnable, `UVM_REG_ADDR_WIDTH'h11B, "RW", 0);
		this.PhyInterruptEnable_PhyTrngCmpltEn = this.PhyInterruptEnable.PhyTrngCmpltEn;
		this.PhyTrngCmpltEn = this.PhyInterruptEnable.PhyTrngCmpltEn;
		this.PhyInterruptEnable_PhyInitCmpltEn = this.PhyInterruptEnable.PhyInitCmpltEn;
		this.PhyInitCmpltEn = this.PhyInterruptEnable.PhyInitCmpltEn;
		this.PhyInterruptEnable_PhyTrngFailEn = this.PhyInterruptEnable.PhyTrngFailEn;
		this.PhyTrngFailEn = this.PhyInterruptEnable.PhyTrngFailEn;
		this.PhyInterruptEnable_PhyFWReservedEn = this.PhyInterruptEnable.PhyFWReservedEn;
		this.PhyFWReservedEn = this.PhyInterruptEnable.PhyFWReservedEn;
		this.PhyInterruptEnable_PhyAcsmParityErrEn = this.PhyInterruptEnable.PhyAcsmParityErrEn;
		this.PhyAcsmParityErrEn = this.PhyInterruptEnable.PhyAcsmParityErrEn;
		this.PhyInterruptEnable_PhyPIEParityErrEn = this.PhyInterruptEnable.PhyPIEParityErrEn;
		this.PhyPIEParityErrEn = this.PhyInterruptEnable.PhyPIEParityErrEn;
		this.PhyInterruptEnable_PhyRdfPtrChkErrEn = this.PhyInterruptEnable.PhyRdfPtrChkErrEn;
		this.PhyRdfPtrChkErrEn = this.PhyInterruptEnable.PhyRdfPtrChkErrEn;
		this.PhyInterruptEnable_PhyEccEn = this.PhyInterruptEnable.PhyEccEn;
		this.PhyEccEn = this.PhyInterruptEnable.PhyEccEn;
		this.PhyInterruptEnable_PhyPIEProgErrEn = this.PhyInterruptEnable.PhyPIEProgErrEn;
		this.PhyPIEProgErrEn = this.PhyInterruptEnable.PhyPIEProgErrEn;
		this.PhyInterruptEnable_PhyHWReservedEn = this.PhyInterruptEnable.PhyHWReservedEn;
		this.PhyHWReservedEn = this.PhyInterruptEnable.PhyHWReservedEn;
      this.PhyInterruptFWControl = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptFWControl::type_id::create("PhyInterruptFWControl",,get_full_name());
      if(this.PhyInterruptFWControl.has_coverage(UVM_CVR_ALL))
      	this.PhyInterruptFWControl.cg_bits.option.name = {get_name(), ".", "PhyInterruptFWControl_bits"};
      this.PhyInterruptFWControl.configure(this, null, "");
      this.PhyInterruptFWControl.build();
      this.default_map.add_reg(this.PhyInterruptFWControl, `UVM_REG_ADDR_WIDTH'h11C, "RW", 0);
		this.PhyInterruptFWControl_PhyTrngCmpltFW = this.PhyInterruptFWControl.PhyTrngCmpltFW;
		this.PhyTrngCmpltFW = this.PhyInterruptFWControl.PhyTrngCmpltFW;
		this.PhyInterruptFWControl_PhyInitCmpltFW = this.PhyInterruptFWControl.PhyInitCmpltFW;
		this.PhyInitCmpltFW = this.PhyInterruptFWControl.PhyInitCmpltFW;
		this.PhyInterruptFWControl_PhyTrngFailFW = this.PhyInterruptFWControl.PhyTrngFailFW;
		this.PhyTrngFailFW = this.PhyInterruptFWControl.PhyTrngFailFW;
		this.PhyInterruptFWControl_PhyFWReservedFW = this.PhyInterruptFWControl.PhyFWReservedFW;
		this.PhyFWReservedFW = this.PhyInterruptFWControl.PhyFWReservedFW;
      this.PhyInterruptMask = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptMask::type_id::create("PhyInterruptMask",,get_full_name());
      if(this.PhyInterruptMask.has_coverage(UVM_CVR_ALL))
      	this.PhyInterruptMask.cg_bits.option.name = {get_name(), ".", "PhyInterruptMask_bits"};
      this.PhyInterruptMask.configure(this, null, "");
      this.PhyInterruptMask.build();
      this.default_map.add_reg(this.PhyInterruptMask, `UVM_REG_ADDR_WIDTH'h11D, "RW", 0);
		this.PhyInterruptMask_PhyTrngCmpltMsk = this.PhyInterruptMask.PhyTrngCmpltMsk;
		this.PhyTrngCmpltMsk = this.PhyInterruptMask.PhyTrngCmpltMsk;
		this.PhyInterruptMask_PhyInitCmpltMsk = this.PhyInterruptMask.PhyInitCmpltMsk;
		this.PhyInitCmpltMsk = this.PhyInterruptMask.PhyInitCmpltMsk;
		this.PhyInterruptMask_PhyTrngFailMsk = this.PhyInterruptMask.PhyTrngFailMsk;
		this.PhyTrngFailMsk = this.PhyInterruptMask.PhyTrngFailMsk;
		this.PhyInterruptMask_PhyFWReservedMsk = this.PhyInterruptMask.PhyFWReservedMsk;
		this.PhyFWReservedMsk = this.PhyInterruptMask.PhyFWReservedMsk;
		this.PhyInterruptMask_PhyAcsmParityErrMsk = this.PhyInterruptMask.PhyAcsmParityErrMsk;
		this.PhyAcsmParityErrMsk = this.PhyInterruptMask.PhyAcsmParityErrMsk;
		this.PhyInterruptMask_PhyPIEParityErrMsk = this.PhyInterruptMask.PhyPIEParityErrMsk;
		this.PhyPIEParityErrMsk = this.PhyInterruptMask.PhyPIEParityErrMsk;
		this.PhyInterruptMask_PhyRdfPtrChkErrMsk = this.PhyInterruptMask.PhyRdfPtrChkErrMsk;
		this.PhyRdfPtrChkErrMsk = this.PhyInterruptMask.PhyRdfPtrChkErrMsk;
		this.PhyInterruptMask_PhyEccMsk = this.PhyInterruptMask.PhyEccMsk;
		this.PhyEccMsk = this.PhyInterruptMask.PhyEccMsk;
		this.PhyInterruptMask_PhyPIEProgErrMsk = this.PhyInterruptMask.PhyPIEProgErrMsk;
		this.PhyPIEProgErrMsk = this.PhyInterruptMask.PhyPIEProgErrMsk;
		this.PhyInterruptMask_PhyHWReservedMsk = this.PhyInterruptMask.PhyHWReservedMsk;
		this.PhyHWReservedMsk = this.PhyInterruptMask.PhyHWReservedMsk;
      this.PhyInterruptClear = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptClear::type_id::create("PhyInterruptClear",,get_full_name());
      if(this.PhyInterruptClear.has_coverage(UVM_CVR_ALL))
      	this.PhyInterruptClear.cg_bits.option.name = {get_name(), ".", "PhyInterruptClear_bits"};
      this.PhyInterruptClear.configure(this, null, "");
      this.PhyInterruptClear.build();
      this.default_map.add_reg(this.PhyInterruptClear, `UVM_REG_ADDR_WIDTH'h11E, "RW", 0);
		this.PhyInterruptClear_PhyTrngCmpltClr = this.PhyInterruptClear.PhyTrngCmpltClr;
		this.PhyTrngCmpltClr = this.PhyInterruptClear.PhyTrngCmpltClr;
		this.PhyInterruptClear_PhyInitCmpltClr = this.PhyInterruptClear.PhyInitCmpltClr;
		this.PhyInitCmpltClr = this.PhyInterruptClear.PhyInitCmpltClr;
		this.PhyInterruptClear_PhyTrngFailClr = this.PhyInterruptClear.PhyTrngFailClr;
		this.PhyTrngFailClr = this.PhyInterruptClear.PhyTrngFailClr;
		this.PhyInterruptClear_PhyFWReservedClr = this.PhyInterruptClear.PhyFWReservedClr;
		this.PhyFWReservedClr = this.PhyInterruptClear.PhyFWReservedClr;
		this.PhyInterruptClear_PhyAcsmParityErrClr = this.PhyInterruptClear.PhyAcsmParityErrClr;
		this.PhyAcsmParityErrClr = this.PhyInterruptClear.PhyAcsmParityErrClr;
		this.PhyInterruptClear_PhyPIEParityErrClr = this.PhyInterruptClear.PhyPIEParityErrClr;
		this.PhyPIEParityErrClr = this.PhyInterruptClear.PhyPIEParityErrClr;
		this.PhyInterruptClear_PhyRdfPtrChkErrClr = this.PhyInterruptClear.PhyRdfPtrChkErrClr;
		this.PhyRdfPtrChkErrClr = this.PhyInterruptClear.PhyRdfPtrChkErrClr;
		this.PhyInterruptClear_PhyEccClr = this.PhyInterruptClear.PhyEccClr;
		this.PhyEccClr = this.PhyInterruptClear.PhyEccClr;
		this.PhyInterruptClear_PhyPIEProgErrClr = this.PhyInterruptClear.PhyPIEProgErrClr;
		this.PhyPIEProgErrClr = this.PhyInterruptClear.PhyPIEProgErrClr;
		this.PhyInterruptClear_PhyHWReservedClr = this.PhyInterruptClear.PhyHWReservedClr;
		this.PhyHWReservedClr = this.PhyInterruptClear.PhyHWReservedClr;
      this.PhyInterruptStatus = ral_reg_DWC_DDRPHYA_PPGC0_p0_PhyInterruptStatus::type_id::create("PhyInterruptStatus",,get_full_name());
      if(this.PhyInterruptStatus.has_coverage(UVM_CVR_ALL))
      	this.PhyInterruptStatus.cg_bits.option.name = {get_name(), ".", "PhyInterruptStatus_bits"};
      this.PhyInterruptStatus.configure(this, null, "");
      this.PhyInterruptStatus.build();
      this.default_map.add_reg(this.PhyInterruptStatus, `UVM_REG_ADDR_WIDTH'h11F, "RO", 0);
		this.PhyInterruptStatus_PhyTrngCmplt = this.PhyInterruptStatus.PhyTrngCmplt;
		this.PhyTrngCmplt = this.PhyInterruptStatus.PhyTrngCmplt;
		this.PhyInterruptStatus_PhyInitCmplt = this.PhyInterruptStatus.PhyInitCmplt;
		this.PhyInitCmplt = this.PhyInterruptStatus.PhyInitCmplt;
		this.PhyInterruptStatus_PhyTrngFail = this.PhyInterruptStatus.PhyTrngFail;
		this.PhyTrngFail = this.PhyInterruptStatus.PhyTrngFail;
		this.PhyInterruptStatus_PhyFWReserved = this.PhyInterruptStatus.PhyFWReserved;
		this.PhyFWReserved = this.PhyInterruptStatus.PhyFWReserved;
		this.PhyInterruptStatus_PhyAcsmParityErr = this.PhyInterruptStatus.PhyAcsmParityErr;
		this.PhyAcsmParityErr = this.PhyInterruptStatus.PhyAcsmParityErr;
		this.PhyInterruptStatus_PhyPIEParityErr = this.PhyInterruptStatus.PhyPIEParityErr;
		this.PhyPIEParityErr = this.PhyInterruptStatus.PhyPIEParityErr;
		this.PhyInterruptStatus_PhyRdfPtrChkErr = this.PhyInterruptStatus.PhyRdfPtrChkErr;
		this.PhyRdfPtrChkErr = this.PhyInterruptStatus.PhyRdfPtrChkErr;
		this.PhyInterruptStatus_PhyEccErr = this.PhyInterruptStatus.PhyEccErr;
		this.PhyEccErr = this.PhyInterruptStatus.PhyEccErr;
		this.PhyInterruptStatus_PhyPIEProgErr = this.PhyInterruptStatus.PhyPIEProgErr;
		this.PhyPIEProgErr = this.PhyInterruptStatus.PhyPIEProgErr;
		this.PhyInterruptStatus_PhyHWReserved = this.PhyInterruptStatus.PhyHWReserved;
		this.PhyHWReserved = this.PhyInterruptStatus.PhyHWReserved;
      this.ACSMRunCtrl = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRunCtrl::type_id::create("ACSMRunCtrl",,get_full_name());
      if(this.ACSMRunCtrl.has_coverage(UVM_CVR_ALL))
      	this.ACSMRunCtrl.cg_bits.option.name = {get_name(), ".", "ACSMRunCtrl_bits"};
      this.ACSMRunCtrl.configure(this, null, "");
      this.ACSMRunCtrl.build();
      this.default_map.add_reg(this.ACSMRunCtrl, `UVM_REG_ADDR_WIDTH'h120, "RW", 0);
		this.ACSMRunCtrl_ACSMRun = this.ACSMRunCtrl.ACSMRun;
		this.ACSMRun = this.ACSMRunCtrl.ACSMRun;
		this.ACSMRunCtrl_AcsmProgPtr = this.ACSMRunCtrl.AcsmProgPtr;
		this.AcsmProgPtr = this.ACSMRunCtrl.AcsmProgPtr;
		this.ACSMRunCtrl_ACSMXlatEn = this.ACSMRunCtrl.ACSMXlatEn;
		this.ACSMXlatEn = this.ACSMRunCtrl.ACSMXlatEn;
		this.ACSMRunCtrl_ACSMNopFlag = this.ACSMRunCtrl.ACSMNopFlag;
		this.ACSMNopFlag = this.ACSMRunCtrl.ACSMNopFlag;
		this.ACSMRunCtrl_ACSMRptCntOverrideEn = this.ACSMRunCtrl.ACSMRptCntOverrideEn;
		this.ACSMRptCntOverrideEn = this.ACSMRunCtrl.ACSMRptCntOverrideEn;
      this.ACSMDone = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDone::type_id::create("ACSMDone",,get_full_name());
      if(this.ACSMDone.has_coverage(UVM_CVR_ALL))
      	this.ACSMDone.cg_bits.option.name = {get_name(), ".", "ACSMDone_bits"};
      this.ACSMDone.configure(this, null, "");
      this.ACSMDone.build();
      this.default_map.add_reg(this.ACSMDone, `UVM_REG_ADDR_WIDTH'h121, "RO", 0);
		this.ACSMDone_ACSMDone = this.ACSMDone.ACSMDone;
      this.ACSMStartAddr_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStartAddr_p0::type_id::create("ACSMStartAddr_p0",,get_full_name());
      if(this.ACSMStartAddr_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMStartAddr_p0.cg_bits.option.name = {get_name(), ".", "ACSMStartAddr_p0_bits"};
      this.ACSMStartAddr_p0.configure(this, null, "");
      this.ACSMStartAddr_p0.build();
      this.default_map.add_reg(this.ACSMStartAddr_p0, `UVM_REG_ADDR_WIDTH'h122, "RW", 0);
		this.ACSMStartAddr_p0_ACSMStartAddr_p0 = this.ACSMStartAddr_p0.ACSMStartAddr_p0;
      this.ACSMStopAddr_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStopAddr_p0::type_id::create("ACSMStopAddr_p0",,get_full_name());
      if(this.ACSMStopAddr_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMStopAddr_p0.cg_bits.option.name = {get_name(), ".", "ACSMStopAddr_p0_bits"};
      this.ACSMStopAddr_p0.configure(this, null, "");
      this.ACSMStopAddr_p0.build();
      this.default_map.add_reg(this.ACSMStopAddr_p0, `UVM_REG_ADDR_WIDTH'h123, "RW", 0);
		this.ACSMStopAddr_p0_ACSMStopAddr_p0 = this.ACSMStopAddr_p0.ACSMStopAddr_p0;
      this.ACSMLastAddr = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLastAddr::type_id::create("ACSMLastAddr",,get_full_name());
      if(this.ACSMLastAddr.has_coverage(UVM_CVR_ALL))
      	this.ACSMLastAddr.cg_bits.option.name = {get_name(), ".", "ACSMLastAddr_bits"};
      this.ACSMLastAddr.configure(this, null, "");
      this.ACSMLastAddr.build();
      this.default_map.add_reg(this.ACSMLastAddr, `UVM_REG_ADDR_WIDTH'h124, "RO", 0);
		this.ACSMLastAddr_ACSMLastAddr = this.ACSMLastAddr.ACSMLastAddr;
      this.ACSMAlgaIncVal = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAlgaIncVal::type_id::create("ACSMAlgaIncVal",,get_full_name());
      if(this.ACSMAlgaIncVal.has_coverage(UVM_CVR_ALL))
      	this.ACSMAlgaIncVal.cg_bits.option.name = {get_name(), ".", "ACSMAlgaIncVal_bits"};
      this.ACSMAlgaIncVal.configure(this, null, "");
      this.ACSMAlgaIncVal.build();
      this.default_map.add_reg(this.ACSMAlgaIncVal, `UVM_REG_ADDR_WIDTH'h125, "RW", 0);
		this.ACSMAlgaIncVal_ACSMAlgaIncVal = this.ACSMAlgaIncVal.ACSMAlgaIncVal;
      this.ACSMAddressMask = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMAddressMask::type_id::create("ACSMAddressMask",,get_full_name());
      if(this.ACSMAddressMask.has_coverage(UVM_CVR_ALL))
      	this.ACSMAddressMask.cg_bits.option.name = {get_name(), ".", "ACSMAddressMask_bits"};
      this.ACSMAddressMask.configure(this, null, "");
      this.ACSMAddressMask.build();
      this.default_map.add_reg(this.ACSMAddressMask, `UVM_REG_ADDR_WIDTH'h126, "RW", 0);
		this.ACSMAddressMask_ACSMAddressMask = this.ACSMAddressMask.ACSMAddressMask;
      this.ACSMOuterLoopRepeatCnt = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMOuterLoopRepeatCnt::type_id::create("ACSMOuterLoopRepeatCnt",,get_full_name());
      if(this.ACSMOuterLoopRepeatCnt.has_coverage(UVM_CVR_ALL))
      	this.ACSMOuterLoopRepeatCnt.cg_bits.option.name = {get_name(), ".", "ACSMOuterLoopRepeatCnt_bits"};
      this.ACSMOuterLoopRepeatCnt.configure(this, null, "");
      this.ACSMOuterLoopRepeatCnt.build();
      this.default_map.add_reg(this.ACSMOuterLoopRepeatCnt, `UVM_REG_ADDR_WIDTH'h127, "RW", 0);
		this.ACSMOuterLoopRepeatCnt_ACSMOuterLoopRepeatCnt = this.ACSMOuterLoopRepeatCnt.ACSMOuterLoopRepeatCnt;
      this.ACSMCkeControl = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeControl::type_id::create("ACSMCkeControl",,get_full_name());
      if(this.ACSMCkeControl.has_coverage(UVM_CVR_ALL))
      	this.ACSMCkeControl.cg_bits.option.name = {get_name(), ".", "ACSMCkeControl_bits"};
      this.ACSMCkeControl.configure(this, null, "");
      this.ACSMCkeControl.build();
      this.default_map.add_reg(this.ACSMCkeControl, `UVM_REG_ADDR_WIDTH'h128, "RW", 0);
		this.ACSMCkeControl_ACSMCkeControl = this.ACSMCkeControl.ACSMCkeControl;
      this.ACSMCkeStatus = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMCkeStatus::type_id::create("ACSMCkeStatus",,get_full_name());
      if(this.ACSMCkeStatus.has_coverage(UVM_CVR_ALL))
      	this.ACSMCkeStatus.cg_bits.option.name = {get_name(), ".", "ACSMCkeStatus_bits"};
      this.ACSMCkeStatus.configure(this, null, "");
      this.ACSMCkeStatus.build();
      this.default_map.add_reg(this.ACSMCkeStatus, `UVM_REG_ADDR_WIDTH'h129, "RO", 0);
		this.ACSMCkeStatus_ACSMCkeStatus = this.ACSMCkeStatus.ACSMCkeStatus;
      this.ACSMWckEnControl = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnControl::type_id::create("ACSMWckEnControl",,get_full_name());
      if(this.ACSMWckEnControl.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckEnControl.cg_bits.option.name = {get_name(), ".", "ACSMWckEnControl_bits"};
      this.ACSMWckEnControl.configure(this, null, "");
      this.ACSMWckEnControl.build();
      this.default_map.add_reg(this.ACSMWckEnControl, `UVM_REG_ADDR_WIDTH'h12A, "RW", 0);
		this.ACSMWckEnControl_ACSMWckEnControl = this.ACSMWckEnControl.ACSMWckEnControl;
      this.ACSMWckEnStatus = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckEnStatus::type_id::create("ACSMWckEnStatus",,get_full_name());
      if(this.ACSMWckEnStatus.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckEnStatus.cg_bits.option.name = {get_name(), ".", "ACSMWckEnStatus_bits"};
      this.ACSMWckEnStatus.configure(this, null, "");
      this.ACSMWckEnStatus.build();
      this.default_map.add_reg(this.ACSMWckEnStatus, `UVM_REG_ADDR_WIDTH'h12B, "RO", 0);
		this.ACSMWckEnStatus_ACSMWckEnStatus = this.ACSMWckEnStatus.ACSMWckEnStatus;
      this.ACSMRxEnPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxEnPulse_p0::type_id::create("ACSMRxEnPulse_p0",,get_full_name());
      if(this.ACSMRxEnPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMRxEnPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMRxEnPulse_p0_bits"};
      this.ACSMRxEnPulse_p0.configure(this, null, "");
      this.ACSMRxEnPulse_p0.build();
      this.default_map.add_reg(this.ACSMRxEnPulse_p0, `UVM_REG_ADDR_WIDTH'h12C, "RW", 0);
		this.ACSMRxEnPulse_p0_ACSMRxEnDelay = this.ACSMRxEnPulse_p0.ACSMRxEnDelay;
		this.ACSMRxEnDelay = this.ACSMRxEnPulse_p0.ACSMRxEnDelay;
		this.ACSMRxEnPulse_p0_ACSMRxEnDelayReserved = this.ACSMRxEnPulse_p0.ACSMRxEnDelayReserved;
		this.ACSMRxEnDelayReserved = this.ACSMRxEnPulse_p0.ACSMRxEnDelayReserved;
		this.ACSMRxEnPulse_p0_ACSMRxEnWidth = this.ACSMRxEnPulse_p0.ACSMRxEnWidth;
		this.ACSMRxEnWidth = this.ACSMRxEnPulse_p0.ACSMRxEnWidth;
      this.ACSMRxValPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRxValPulse_p0::type_id::create("ACSMRxValPulse_p0",,get_full_name());
      if(this.ACSMRxValPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMRxValPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMRxValPulse_p0_bits"};
      this.ACSMRxValPulse_p0.configure(this, null, "");
      this.ACSMRxValPulse_p0.build();
      this.default_map.add_reg(this.ACSMRxValPulse_p0, `UVM_REG_ADDR_WIDTH'h12D, "RW", 0);
		this.ACSMRxValPulse_p0_ACSMRxValDelay = this.ACSMRxValPulse_p0.ACSMRxValDelay;
		this.ACSMRxValDelay = this.ACSMRxValPulse_p0.ACSMRxValDelay;
		this.ACSMRxValPulse_p0_ACSMRxValDelayReserved = this.ACSMRxValPulse_p0.ACSMRxValDelayReserved;
		this.ACSMRxValDelayReserved = this.ACSMRxValPulse_p0.ACSMRxValDelayReserved;
		this.ACSMRxValPulse_p0_ACSMRxValWidth = this.ACSMRxValPulse_p0.ACSMRxValWidth;
		this.ACSMRxValWidth = this.ACSMRxValPulse_p0.ACSMRxValWidth;
      this.ACSMTxEnPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMTxEnPulse_p0::type_id::create("ACSMTxEnPulse_p0",,get_full_name());
      if(this.ACSMTxEnPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMTxEnPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMTxEnPulse_p0_bits"};
      this.ACSMTxEnPulse_p0.configure(this, null, "");
      this.ACSMTxEnPulse_p0.build();
      this.default_map.add_reg(this.ACSMTxEnPulse_p0, `UVM_REG_ADDR_WIDTH'h12E, "RW", 0);
		this.ACSMTxEnPulse_p0_ACSMTxEnDelay = this.ACSMTxEnPulse_p0.ACSMTxEnDelay;
		this.ACSMTxEnDelay = this.ACSMTxEnPulse_p0.ACSMTxEnDelay;
		this.ACSMTxEnPulse_p0_ACSMTxEnDelayReserved = this.ACSMTxEnPulse_p0.ACSMTxEnDelayReserved;
		this.ACSMTxEnDelayReserved = this.ACSMTxEnPulse_p0.ACSMTxEnDelayReserved;
		this.ACSMTxEnPulse_p0_ACSMTxEnWidth = this.ACSMTxEnPulse_p0.ACSMTxEnWidth;
		this.ACSMTxEnWidth = this.ACSMTxEnPulse_p0.ACSMTxEnWidth;
      this.ACSMWrcsPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWrcsPulse_p0::type_id::create("ACSMWrcsPulse_p0",,get_full_name());
      if(this.ACSMWrcsPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWrcsPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWrcsPulse_p0_bits"};
      this.ACSMWrcsPulse_p0.configure(this, null, "");
      this.ACSMWrcsPulse_p0.build();
      this.default_map.add_reg(this.ACSMWrcsPulse_p0, `UVM_REG_ADDR_WIDTH'h12F, "RW", 0);
		this.ACSMWrcsPulse_p0_ACSMWrcsDelay = this.ACSMWrcsPulse_p0.ACSMWrcsDelay;
		this.ACSMWrcsDelay = this.ACSMWrcsPulse_p0.ACSMWrcsDelay;
		this.ACSMWrcsPulse_p0_ACSMWrcsDelayReserved = this.ACSMWrcsPulse_p0.ACSMWrcsDelayReserved;
		this.ACSMWrcsDelayReserved = this.ACSMWrcsPulse_p0.ACSMWrcsDelayReserved;
		this.ACSMWrcsPulse_p0_ACSMWrcsWidth = this.ACSMWrcsPulse_p0.ACSMWrcsWidth;
		this.ACSMWrcsWidth = this.ACSMWrcsPulse_p0.ACSMWrcsWidth;
      this.ACSMRdcsPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRdcsPulse_p0::type_id::create("ACSMRdcsPulse_p0",,get_full_name());
      if(this.ACSMRdcsPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMRdcsPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMRdcsPulse_p0_bits"};
      this.ACSMRdcsPulse_p0.configure(this, null, "");
      this.ACSMRdcsPulse_p0.build();
      this.default_map.add_reg(this.ACSMRdcsPulse_p0, `UVM_REG_ADDR_WIDTH'h130, "RW", 0);
		this.ACSMRdcsPulse_p0_ACSMRdcsDelay = this.ACSMRdcsPulse_p0.ACSMRdcsDelay;
		this.ACSMRdcsDelay = this.ACSMRdcsPulse_p0.ACSMRdcsDelay;
		this.ACSMRdcsPulse_p0_ACSMRdcsDelayReserved = this.ACSMRdcsPulse_p0.ACSMRdcsDelayReserved;
		this.ACSMRdcsDelayReserved = this.ACSMRdcsPulse_p0.ACSMRdcsDelayReserved;
		this.ACSMRdcsPulse_p0_ACSMRdcsWidth = this.ACSMRdcsPulse_p0.ACSMRdcsWidth;
		this.ACSMRdcsWidth = this.ACSMRdcsPulse_p0.ACSMRdcsWidth;
      this.ACSMInfiniteOLRC = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMInfiniteOLRC::type_id::create("ACSMInfiniteOLRC",,get_full_name());
      if(this.ACSMInfiniteOLRC.has_coverage(UVM_CVR_ALL))
      	this.ACSMInfiniteOLRC.cg_bits.option.name = {get_name(), ".", "ACSMInfiniteOLRC_bits"};
      this.ACSMInfiniteOLRC.configure(this, null, "");
      this.ACSMInfiniteOLRC.build();
      this.default_map.add_reg(this.ACSMInfiniteOLRC, `UVM_REG_ADDR_WIDTH'h131, "RW", 0);
		this.ACSMInfiniteOLRC_ACSMInfiniteOLRC = this.ACSMInfiniteOLRC.ACSMInfiniteOLRC;
      this.ACSMDefaultAddr = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultAddr::type_id::create("ACSMDefaultAddr",,get_full_name());
      if(this.ACSMDefaultAddr.has_coverage(UVM_CVR_ALL))
      	this.ACSMDefaultAddr.cg_bits.option.name = {get_name(), ".", "ACSMDefaultAddr_bits"};
      this.ACSMDefaultAddr.configure(this, null, "");
      this.ACSMDefaultAddr.build();
      this.default_map.add_reg(this.ACSMDefaultAddr, `UVM_REG_ADDR_WIDTH'h132, "RW", 0);
		this.ACSMDefaultAddr_ACSMDefaultAddr = this.ACSMDefaultAddr.ACSMDefaultAddr;
      this.ACSMDefaultCs = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMDefaultCs::type_id::create("ACSMDefaultCs",,get_full_name());
      if(this.ACSMDefaultCs.has_coverage(UVM_CVR_ALL))
      	this.ACSMDefaultCs.cg_bits.option.name = {get_name(), ".", "ACSMDefaultCs_bits"};
      this.ACSMDefaultCs.configure(this, null, "");
      this.ACSMDefaultCs.build();
      this.default_map.add_reg(this.ACSMDefaultCs, `UVM_REG_ADDR_WIDTH'h133, "RW", 0);
		this.ACSMDefaultCs_ACSMDefaultCs = this.ACSMDefaultCs.ACSMDefaultCs;
      this.ACSMStaticCtrl = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMStaticCtrl::type_id::create("ACSMStaticCtrl",,get_full_name());
      if(this.ACSMStaticCtrl.has_coverage(UVM_CVR_ALL))
      	this.ACSMStaticCtrl.cg_bits.option.name = {get_name(), ".", "ACSMStaticCtrl_bits"};
      this.ACSMStaticCtrl.configure(this, null, "");
      this.ACSMStaticCtrl.build();
      this.default_map.add_reg(this.ACSMStaticCtrl, `UVM_REG_ADDR_WIDTH'h134, "RW", 0);
		this.ACSMStaticCtrl_ACSMPhaseControl = this.ACSMStaticCtrl.ACSMPhaseControl;
		this.ACSMPhaseControl = this.ACSMStaticCtrl.ACSMPhaseControl;
      this.ACSMWckWriteStaticLoPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticLoPulse_p0::type_id::create("ACSMWckWriteStaticLoPulse_p0",,get_full_name());
      if(this.ACSMWckWriteStaticLoPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckWriteStaticLoPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckWriteStaticLoPulse_p0_bits"};
      this.ACSMWckWriteStaticLoPulse_p0.configure(this, null, "");
      this.ACSMWckWriteStaticLoPulse_p0.build();
      this.default_map.add_reg(this.ACSMWckWriteStaticLoPulse_p0, `UVM_REG_ADDR_WIDTH'h135, "RW", 0);
		this.ACSMWckWriteStaticLoPulse_p0_ACSMWckWriteStaticLoDelay = this.ACSMWckWriteStaticLoPulse_p0.ACSMWckWriteStaticLoDelay;
		this.ACSMWckWriteStaticLoDelay = this.ACSMWckWriteStaticLoPulse_p0.ACSMWckWriteStaticLoDelay;
		this.ACSMWckWriteStaticLoPulse_p0_ACSMWckWriteStaticLoDelayReserved = this.ACSMWckWriteStaticLoPulse_p0.ACSMWckWriteStaticLoDelayReserved;
		this.ACSMWckWriteStaticLoDelayReserved = this.ACSMWckWriteStaticLoPulse_p0.ACSMWckWriteStaticLoDelayReserved;
		this.ACSMWckWriteStaticLoPulse_p0_ACSMWckWriteStaticLoWidth = this.ACSMWckWriteStaticLoPulse_p0.ACSMWckWriteStaticLoWidth;
		this.ACSMWckWriteStaticLoWidth = this.ACSMWckWriteStaticLoPulse_p0.ACSMWckWriteStaticLoWidth;
      this.ACSMWckWriteStaticHiPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteStaticHiPulse_p0::type_id::create("ACSMWckWriteStaticHiPulse_p0",,get_full_name());
      if(this.ACSMWckWriteStaticHiPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckWriteStaticHiPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckWriteStaticHiPulse_p0_bits"};
      this.ACSMWckWriteStaticHiPulse_p0.configure(this, null, "");
      this.ACSMWckWriteStaticHiPulse_p0.build();
      this.default_map.add_reg(this.ACSMWckWriteStaticHiPulse_p0, `UVM_REG_ADDR_WIDTH'h136, "RW", 0);
		this.ACSMWckWriteStaticHiPulse_p0_ACSMWckWriteStaticHiDelay = this.ACSMWckWriteStaticHiPulse_p0.ACSMWckWriteStaticHiDelay;
		this.ACSMWckWriteStaticHiDelay = this.ACSMWckWriteStaticHiPulse_p0.ACSMWckWriteStaticHiDelay;
		this.ACSMWckWriteStaticHiPulse_p0_ACSMWckWriteStaticHiDelayReserved = this.ACSMWckWriteStaticHiPulse_p0.ACSMWckWriteStaticHiDelayReserved;
		this.ACSMWckWriteStaticHiDelayReserved = this.ACSMWckWriteStaticHiPulse_p0.ACSMWckWriteStaticHiDelayReserved;
		this.ACSMWckWriteStaticHiPulse_p0_ACSMWckWriteStaticHiWidth = this.ACSMWckWriteStaticHiPulse_p0.ACSMWckWriteStaticHiWidth;
		this.ACSMWckWriteStaticHiWidth = this.ACSMWckWriteStaticHiPulse_p0.ACSMWckWriteStaticHiWidth;
      this.ACSMWckWriteTogglePulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteTogglePulse_p0::type_id::create("ACSMWckWriteTogglePulse_p0",,get_full_name());
      if(this.ACSMWckWriteTogglePulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckWriteTogglePulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckWriteTogglePulse_p0_bits"};
      this.ACSMWckWriteTogglePulse_p0.configure(this, null, "");
      this.ACSMWckWriteTogglePulse_p0.build();
      this.default_map.add_reg(this.ACSMWckWriteTogglePulse_p0, `UVM_REG_ADDR_WIDTH'h137, "RW", 0);
		this.ACSMWckWriteTogglePulse_p0_ACSMWckWriteToggleDelay = this.ACSMWckWriteTogglePulse_p0.ACSMWckWriteToggleDelay;
		this.ACSMWckWriteToggleDelay = this.ACSMWckWriteTogglePulse_p0.ACSMWckWriteToggleDelay;
		this.ACSMWckWriteTogglePulse_p0_ACSMWckWriteToggleDelayReserved = this.ACSMWckWriteTogglePulse_p0.ACSMWckWriteToggleDelayReserved;
		this.ACSMWckWriteToggleDelayReserved = this.ACSMWckWriteTogglePulse_p0.ACSMWckWriteToggleDelayReserved;
		this.ACSMWckWriteTogglePulse_p0_ACSMWckWriteToggleWidth = this.ACSMWckWriteTogglePulse_p0.ACSMWckWriteToggleWidth;
		this.ACSMWckWriteToggleWidth = this.ACSMWckWriteTogglePulse_p0.ACSMWckWriteToggleWidth;
      this.ACSMWckWriteFastTogglePulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckWriteFastTogglePulse_p0::type_id::create("ACSMWckWriteFastTogglePulse_p0",,get_full_name());
      if(this.ACSMWckWriteFastTogglePulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckWriteFastTogglePulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckWriteFastTogglePulse_p0_bits"};
      this.ACSMWckWriteFastTogglePulse_p0.configure(this, null, "");
      this.ACSMWckWriteFastTogglePulse_p0.build();
      this.default_map.add_reg(this.ACSMWckWriteFastTogglePulse_p0, `UVM_REG_ADDR_WIDTH'h138, "RW", 0);
		this.ACSMWckWriteFastTogglePulse_p0_ACSMWckWriteFastToggleDelay = this.ACSMWckWriteFastTogglePulse_p0.ACSMWckWriteFastToggleDelay;
		this.ACSMWckWriteFastToggleDelay = this.ACSMWckWriteFastTogglePulse_p0.ACSMWckWriteFastToggleDelay;
		this.ACSMWckWriteFastTogglePulse_p0_ACSMWckWriteFastToggleDelayReserved = this.ACSMWckWriteFastTogglePulse_p0.ACSMWckWriteFastToggleDelayReserved;
		this.ACSMWckWriteFastToggleDelayReserved = this.ACSMWckWriteFastTogglePulse_p0.ACSMWckWriteFastToggleDelayReserved;
		this.ACSMWckWriteFastTogglePulse_p0_ACSMWckWriteFastToggleWidth = this.ACSMWckWriteFastTogglePulse_p0.ACSMWckWriteFastToggleWidth;
		this.ACSMWckWriteFastToggleWidth = this.ACSMWckWriteFastTogglePulse_p0.ACSMWckWriteFastToggleWidth;
      this.ACSMWckReadStaticLoPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticLoPulse_p0::type_id::create("ACSMWckReadStaticLoPulse_p0",,get_full_name());
      if(this.ACSMWckReadStaticLoPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckReadStaticLoPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckReadStaticLoPulse_p0_bits"};
      this.ACSMWckReadStaticLoPulse_p0.configure(this, null, "");
      this.ACSMWckReadStaticLoPulse_p0.build();
      this.default_map.add_reg(this.ACSMWckReadStaticLoPulse_p0, `UVM_REG_ADDR_WIDTH'h139, "RW", 0);
		this.ACSMWckReadStaticLoPulse_p0_ACSMWckReadStaticLoDelay = this.ACSMWckReadStaticLoPulse_p0.ACSMWckReadStaticLoDelay;
		this.ACSMWckReadStaticLoDelay = this.ACSMWckReadStaticLoPulse_p0.ACSMWckReadStaticLoDelay;
		this.ACSMWckReadStaticLoPulse_p0_ACSMWckReadStaticLoDelayReserved = this.ACSMWckReadStaticLoPulse_p0.ACSMWckReadStaticLoDelayReserved;
		this.ACSMWckReadStaticLoDelayReserved = this.ACSMWckReadStaticLoPulse_p0.ACSMWckReadStaticLoDelayReserved;
		this.ACSMWckReadStaticLoPulse_p0_ACSMWckReadStaticLoWidth = this.ACSMWckReadStaticLoPulse_p0.ACSMWckReadStaticLoWidth;
		this.ACSMWckReadStaticLoWidth = this.ACSMWckReadStaticLoPulse_p0.ACSMWckReadStaticLoWidth;
      this.ACSMWckReadStaticHiPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadStaticHiPulse_p0::type_id::create("ACSMWckReadStaticHiPulse_p0",,get_full_name());
      if(this.ACSMWckReadStaticHiPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckReadStaticHiPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckReadStaticHiPulse_p0_bits"};
      this.ACSMWckReadStaticHiPulse_p0.configure(this, null, "");
      this.ACSMWckReadStaticHiPulse_p0.build();
      this.default_map.add_reg(this.ACSMWckReadStaticHiPulse_p0, `UVM_REG_ADDR_WIDTH'h13A, "RW", 0);
		this.ACSMWckReadStaticHiPulse_p0_ACSMWckReadStaticHiDelay = this.ACSMWckReadStaticHiPulse_p0.ACSMWckReadStaticHiDelay;
		this.ACSMWckReadStaticHiDelay = this.ACSMWckReadStaticHiPulse_p0.ACSMWckReadStaticHiDelay;
		this.ACSMWckReadStaticHiPulse_p0_ACSMWckReadStaticHiDelayReserved = this.ACSMWckReadStaticHiPulse_p0.ACSMWckReadStaticHiDelayReserved;
		this.ACSMWckReadStaticHiDelayReserved = this.ACSMWckReadStaticHiPulse_p0.ACSMWckReadStaticHiDelayReserved;
		this.ACSMWckReadStaticHiPulse_p0_ACSMWckReadStaticHiWidth = this.ACSMWckReadStaticHiPulse_p0.ACSMWckReadStaticHiWidth;
		this.ACSMWckReadStaticHiWidth = this.ACSMWckReadStaticHiPulse_p0.ACSMWckReadStaticHiWidth;
      this.ACSMWckReadTogglePulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadTogglePulse_p0::type_id::create("ACSMWckReadTogglePulse_p0",,get_full_name());
      if(this.ACSMWckReadTogglePulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckReadTogglePulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckReadTogglePulse_p0_bits"};
      this.ACSMWckReadTogglePulse_p0.configure(this, null, "");
      this.ACSMWckReadTogglePulse_p0.build();
      this.default_map.add_reg(this.ACSMWckReadTogglePulse_p0, `UVM_REG_ADDR_WIDTH'h13B, "RW", 0);
		this.ACSMWckReadTogglePulse_p0_ACSMWckReadToggleDelay = this.ACSMWckReadTogglePulse_p0.ACSMWckReadToggleDelay;
		this.ACSMWckReadToggleDelay = this.ACSMWckReadTogglePulse_p0.ACSMWckReadToggleDelay;
		this.ACSMWckReadTogglePulse_p0_ACSMWckReadToggleDelayReserved = this.ACSMWckReadTogglePulse_p0.ACSMWckReadToggleDelayReserved;
		this.ACSMWckReadToggleDelayReserved = this.ACSMWckReadTogglePulse_p0.ACSMWckReadToggleDelayReserved;
		this.ACSMWckReadTogglePulse_p0_ACSMWckReadToggleWidth = this.ACSMWckReadTogglePulse_p0.ACSMWckReadToggleWidth;
		this.ACSMWckReadToggleWidth = this.ACSMWckReadTogglePulse_p0.ACSMWckReadToggleWidth;
      this.ACSMWckReadFastTogglePulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckReadFastTogglePulse_p0::type_id::create("ACSMWckReadFastTogglePulse_p0",,get_full_name());
      if(this.ACSMWckReadFastTogglePulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckReadFastTogglePulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckReadFastTogglePulse_p0_bits"};
      this.ACSMWckReadFastTogglePulse_p0.configure(this, null, "");
      this.ACSMWckReadFastTogglePulse_p0.build();
      this.default_map.add_reg(this.ACSMWckReadFastTogglePulse_p0, `UVM_REG_ADDR_WIDTH'h13C, "RW", 0);
		this.ACSMWckReadFastTogglePulse_p0_ACSMWckReadFastToggleDelay = this.ACSMWckReadFastTogglePulse_p0.ACSMWckReadFastToggleDelay;
		this.ACSMWckReadFastToggleDelay = this.ACSMWckReadFastTogglePulse_p0.ACSMWckReadFastToggleDelay;
		this.ACSMWckReadFastTogglePulse_p0_ACSMWckReadFastToggleDelayReserved = this.ACSMWckReadFastTogglePulse_p0.ACSMWckReadFastToggleDelayReserved;
		this.ACSMWckReadFastToggleDelayReserved = this.ACSMWckReadFastTogglePulse_p0.ACSMWckReadFastToggleDelayReserved;
		this.ACSMWckReadFastTogglePulse_p0_ACSMWckReadFastToggleWidth = this.ACSMWckReadFastTogglePulse_p0.ACSMWckReadFastToggleWidth;
		this.ACSMWckReadFastToggleWidth = this.ACSMWckReadFastTogglePulse_p0.ACSMWckReadFastToggleWidth;
      this.ACSMWckFreqSwStaticLoPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticLoPulse_p0::type_id::create("ACSMWckFreqSwStaticLoPulse_p0",,get_full_name());
      if(this.ACSMWckFreqSwStaticLoPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckFreqSwStaticLoPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckFreqSwStaticLoPulse_p0_bits"};
      this.ACSMWckFreqSwStaticLoPulse_p0.configure(this, null, "");
      this.ACSMWckFreqSwStaticLoPulse_p0.build();
      this.default_map.add_reg(this.ACSMWckFreqSwStaticLoPulse_p0, `UVM_REG_ADDR_WIDTH'h13D, "RW", 0);
		this.ACSMWckFreqSwStaticLoPulse_p0_ACSMWckFreqSwStaticLoDelay = this.ACSMWckFreqSwStaticLoPulse_p0.ACSMWckFreqSwStaticLoDelay;
		this.ACSMWckFreqSwStaticLoDelay = this.ACSMWckFreqSwStaticLoPulse_p0.ACSMWckFreqSwStaticLoDelay;
		this.ACSMWckFreqSwStaticLoPulse_p0_ACSMWckFreqSwStaticLoDelayReserved = this.ACSMWckFreqSwStaticLoPulse_p0.ACSMWckFreqSwStaticLoDelayReserved;
		this.ACSMWckFreqSwStaticLoDelayReserved = this.ACSMWckFreqSwStaticLoPulse_p0.ACSMWckFreqSwStaticLoDelayReserved;
		this.ACSMWckFreqSwStaticLoPulse_p0_ACSMWckFreqSwStaticLoWidth = this.ACSMWckFreqSwStaticLoPulse_p0.ACSMWckFreqSwStaticLoWidth;
		this.ACSMWckFreqSwStaticLoWidth = this.ACSMWckFreqSwStaticLoPulse_p0.ACSMWckFreqSwStaticLoWidth;
      this.ACSMWckFreqSwStaticHiPulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwStaticHiPulse_p0::type_id::create("ACSMWckFreqSwStaticHiPulse_p0",,get_full_name());
      if(this.ACSMWckFreqSwStaticHiPulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckFreqSwStaticHiPulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckFreqSwStaticHiPulse_p0_bits"};
      this.ACSMWckFreqSwStaticHiPulse_p0.configure(this, null, "");
      this.ACSMWckFreqSwStaticHiPulse_p0.build();
      this.default_map.add_reg(this.ACSMWckFreqSwStaticHiPulse_p0, `UVM_REG_ADDR_WIDTH'h13E, "RW", 0);
		this.ACSMWckFreqSwStaticHiPulse_p0_ACSMWckFreqSwStaticHiDelay = this.ACSMWckFreqSwStaticHiPulse_p0.ACSMWckFreqSwStaticHiDelay;
		this.ACSMWckFreqSwStaticHiDelay = this.ACSMWckFreqSwStaticHiPulse_p0.ACSMWckFreqSwStaticHiDelay;
		this.ACSMWckFreqSwStaticHiPulse_p0_ACSMWckFreqSwStaticHiDelayReserved = this.ACSMWckFreqSwStaticHiPulse_p0.ACSMWckFreqSwStaticHiDelayReserved;
		this.ACSMWckFreqSwStaticHiDelayReserved = this.ACSMWckFreqSwStaticHiPulse_p0.ACSMWckFreqSwStaticHiDelayReserved;
		this.ACSMWckFreqSwStaticHiPulse_p0_ACSMWckFreqSwStaticHiWidth = this.ACSMWckFreqSwStaticHiPulse_p0.ACSMWckFreqSwStaticHiWidth;
		this.ACSMWckFreqSwStaticHiWidth = this.ACSMWckFreqSwStaticHiPulse_p0.ACSMWckFreqSwStaticHiWidth;
      this.ACSMWckFreqSwTogglePulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwTogglePulse_p0::type_id::create("ACSMWckFreqSwTogglePulse_p0",,get_full_name());
      if(this.ACSMWckFreqSwTogglePulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckFreqSwTogglePulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckFreqSwTogglePulse_p0_bits"};
      this.ACSMWckFreqSwTogglePulse_p0.configure(this, null, "");
      this.ACSMWckFreqSwTogglePulse_p0.build();
      this.default_map.add_reg(this.ACSMWckFreqSwTogglePulse_p0, `UVM_REG_ADDR_WIDTH'h13F, "RW", 0);
		this.ACSMWckFreqSwTogglePulse_p0_ACSMWckFreqSwToggleDelay = this.ACSMWckFreqSwTogglePulse_p0.ACSMWckFreqSwToggleDelay;
		this.ACSMWckFreqSwToggleDelay = this.ACSMWckFreqSwTogglePulse_p0.ACSMWckFreqSwToggleDelay;
		this.ACSMWckFreqSwTogglePulse_p0_ACSMWckFreqSwToggleDelayReserved = this.ACSMWckFreqSwTogglePulse_p0.ACSMWckFreqSwToggleDelayReserved;
		this.ACSMWckFreqSwToggleDelayReserved = this.ACSMWckFreqSwTogglePulse_p0.ACSMWckFreqSwToggleDelayReserved;
		this.ACSMWckFreqSwTogglePulse_p0_ACSMWckFreqSwToggleWidth = this.ACSMWckFreqSwTogglePulse_p0.ACSMWckFreqSwToggleWidth;
		this.ACSMWckFreqSwToggleWidth = this.ACSMWckFreqSwTogglePulse_p0.ACSMWckFreqSwToggleWidth;
      this.ACSMWckFreqSwFastTogglePulse_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreqSwFastTogglePulse_p0::type_id::create("ACSMWckFreqSwFastTogglePulse_p0",,get_full_name());
      if(this.ACSMWckFreqSwFastTogglePulse_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckFreqSwFastTogglePulse_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckFreqSwFastTogglePulse_p0_bits"};
      this.ACSMWckFreqSwFastTogglePulse_p0.configure(this, null, "");
      this.ACSMWckFreqSwFastTogglePulse_p0.build();
      this.default_map.add_reg(this.ACSMWckFreqSwFastTogglePulse_p0, `UVM_REG_ADDR_WIDTH'h140, "RW", 0);
		this.ACSMWckFreqSwFastTogglePulse_p0_ACSMWckFreqSwFastToggleDelay = this.ACSMWckFreqSwFastTogglePulse_p0.ACSMWckFreqSwFastToggleDelay;
		this.ACSMWckFreqSwFastToggleDelay = this.ACSMWckFreqSwFastTogglePulse_p0.ACSMWckFreqSwFastToggleDelay;
		this.ACSMWckFreqSwFastTogglePulse_p0_ACSMWckFreqSwFastToggleDelayReserved = this.ACSMWckFreqSwFastTogglePulse_p0.ACSMWckFreqSwFastToggleDelayReserved;
		this.ACSMWckFreqSwFastToggleDelayReserved = this.ACSMWckFreqSwFastTogglePulse_p0.ACSMWckFreqSwFastToggleDelayReserved;
		this.ACSMWckFreqSwFastTogglePulse_p0_ACSMWckFreqSwFastToggleWidth = this.ACSMWckFreqSwFastTogglePulse_p0.ACSMWckFreqSwFastToggleWidth;
		this.ACSMWckFreqSwFastToggleWidth = this.ACSMWckFreqSwFastTogglePulse_p0.ACSMWckFreqSwFastToggleWidth;
      this.ACSMWckFreeRunMode_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMWckFreeRunMode_p0::type_id::create("ACSMWckFreeRunMode_p0",,get_full_name());
      if(this.ACSMWckFreeRunMode_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMWckFreeRunMode_p0.cg_bits.option.name = {get_name(), ".", "ACSMWckFreeRunMode_p0_bits"};
      this.ACSMWckFreeRunMode_p0.configure(this, null, "");
      this.ACSMWckFreeRunMode_p0.build();
      this.default_map.add_reg(this.ACSMWckFreeRunMode_p0, `UVM_REG_ADDR_WIDTH'h141, "RW", 0);
		this.ACSMWckFreeRunMode_p0_ACSMWckFreeRunMode_p0 = this.ACSMWckFreeRunMode_p0.ACSMWckFreeRunMode_p0;
      this.ACSMLowSpeedClockEnable = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockEnable::type_id::create("ACSMLowSpeedClockEnable",,get_full_name());
      if(this.ACSMLowSpeedClockEnable.has_coverage(UVM_CVR_ALL))
      	this.ACSMLowSpeedClockEnable.cg_bits.option.name = {get_name(), ".", "ACSMLowSpeedClockEnable_bits"};
      this.ACSMLowSpeedClockEnable.configure(this, null, "");
      this.ACSMLowSpeedClockEnable.build();
      this.default_map.add_reg(this.ACSMLowSpeedClockEnable, `UVM_REG_ADDR_WIDTH'h142, "RW", 0);
		this.ACSMLowSpeedClockEnable_ACSMLowSpeedClockEnable = this.ACSMLowSpeedClockEnable.ACSMLowSpeedClockEnable;
      this.ACSMLowSpeedClockDelay = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMLowSpeedClockDelay::type_id::create("ACSMLowSpeedClockDelay",,get_full_name());
      if(this.ACSMLowSpeedClockDelay.has_coverage(UVM_CVR_ALL))
      	this.ACSMLowSpeedClockDelay.cg_bits.option.name = {get_name(), ".", "ACSMLowSpeedClockDelay_bits"};
      this.ACSMLowSpeedClockDelay.configure(this, null, "");
      this.ACSMLowSpeedClockDelay.build();
      this.default_map.add_reg(this.ACSMLowSpeedClockDelay, `UVM_REG_ADDR_WIDTH'h144, "RW", 0);
		this.ACSMLowSpeedClockDelay_ACSMLowSpeedClockDelay = this.ACSMLowSpeedClockDelay.ACSMLowSpeedClockDelay;
      this.ACSMRptCntOverride_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntOverride_p0::type_id::create("ACSMRptCntOverride_p0",,get_full_name());
      if(this.ACSMRptCntOverride_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMRptCntOverride_p0.cg_bits.option.name = {get_name(), ".", "ACSMRptCntOverride_p0_bits"};
      this.ACSMRptCntOverride_p0.configure(this, null, "");
      this.ACSMRptCntOverride_p0.build();
      this.default_map.add_reg(this.ACSMRptCntOverride_p0, `UVM_REG_ADDR_WIDTH'h145, "RW", 0);
		this.ACSMRptCntOverride_p0_ACSMRptCntOverride_p0 = this.ACSMRptCntOverride_p0.ACSMRptCntOverride_p0;
      this.ACSMRptCntDbl_p0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMRptCntDbl_p0::type_id::create("ACSMRptCntDbl_p0",,get_full_name());
      if(this.ACSMRptCntDbl_p0.has_coverage(UVM_CVR_ALL))
      	this.ACSMRptCntDbl_p0.cg_bits.option.name = {get_name(), ".", "ACSMRptCntDbl_p0_bits"};
      this.ACSMRptCntDbl_p0.configure(this, null, "");
      this.ACSMRptCntDbl_p0.build();
      this.default_map.add_reg(this.ACSMRptCntDbl_p0, `UVM_REG_ADDR_WIDTH'h146, "RW", 0);
		this.ACSMRptCntDbl_p0_ACSMRptCntDbl_p0 = this.ACSMRptCntDbl_p0.ACSMRptCntDbl_p0;
      this.ACSMParityStatus = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityStatus::type_id::create("ACSMParityStatus",,get_full_name());
      if(this.ACSMParityStatus.has_coverage(UVM_CVR_ALL))
      	this.ACSMParityStatus.cg_bits.option.name = {get_name(), ".", "ACSMParityStatus_bits"};
      this.ACSMParityStatus.configure(this, null, "");
      this.ACSMParityStatus.build();
      this.default_map.add_reg(this.ACSMParityStatus, `UVM_REG_ADDR_WIDTH'h147, "RO", 0);
		this.ACSMParityStatus_ACSMParityStatus = this.ACSMParityStatus.ACSMParityStatus;
      this.HwtLpCsEnBypass = ral_reg_DWC_DDRPHYA_PPGC0_p0_HwtLpCsEnBypass::type_id::create("HwtLpCsEnBypass",,get_full_name());
      if(this.HwtLpCsEnBypass.has_coverage(UVM_CVR_ALL))
      	this.HwtLpCsEnBypass.cg_bits.option.name = {get_name(), ".", "HwtLpCsEnBypass_bits"};
      this.HwtLpCsEnBypass.configure(this, null, "");
      this.HwtLpCsEnBypass.build();
      this.default_map.add_reg(this.HwtLpCsEnBypass, `UVM_REG_ADDR_WIDTH'h174, "RW", 0);
		this.HwtLpCsEnBypass_HwtLpCsEnBypass = this.HwtLpCsEnBypass.HwtLpCsEnBypass;
      this.ACSMNopAddr = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMNopAddr::type_id::create("ACSMNopAddr",,get_full_name());
      if(this.ACSMNopAddr.has_coverage(UVM_CVR_ALL))
      	this.ACSMNopAddr.cg_bits.option.name = {get_name(), ".", "ACSMNopAddr_bits"};
      this.ACSMNopAddr.configure(this, null, "");
      this.ACSMNopAddr.build();
      this.default_map.add_reg(this.ACSMNopAddr, `UVM_REG_ADDR_WIDTH'h18A, "RW", 0);
		this.ACSMNopAddr_ACSMNopAddr = this.ACSMNopAddr.ACSMNopAddr;
      this.SnoopCntrl = ral_reg_DWC_DDRPHYA_PPGC0_p0_SnoopCntrl::type_id::create("SnoopCntrl",,get_full_name());
      if(this.SnoopCntrl.has_coverage(UVM_CVR_ALL))
      	this.SnoopCntrl.cg_bits.option.name = {get_name(), ".", "SnoopCntrl_bits"};
      this.SnoopCntrl.configure(this, null, "");
      this.SnoopCntrl.build();
      this.default_map.add_reg(this.SnoopCntrl, `UVM_REG_ADDR_WIDTH'h1A7, "RW", 0);
		this.SnoopCntrl_SnoopCntrl = this.SnoopCntrl.SnoopCntrl;
      this.ACSMParityInvert = ral_reg_DWC_DDRPHYA_PPGC0_p0_ACSMParityInvert::type_id::create("ACSMParityInvert",,get_full_name());
      if(this.ACSMParityInvert.has_coverage(UVM_CVR_ALL))
      	this.ACSMParityInvert.cg_bits.option.name = {get_name(), ".", "ACSMParityInvert_bits"};
      this.ACSMParityInvert.configure(this, null, "");
      this.ACSMParityInvert.build();
      this.default_map.add_reg(this.ACSMParityInvert, `UVM_REG_ADDR_WIDTH'h1A8, "RW", 0);
		this.ACSMParityInvert_ACSMParityInvert = this.ACSMParityInvert.ACSMParityInvert;
      this.AcsmPsIndx = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmPsIndx::type_id::create("AcsmPsIndx",,get_full_name());
      if(this.AcsmPsIndx.has_coverage(UVM_CVR_ALL))
      	this.AcsmPsIndx.cg_bits.option.name = {get_name(), ".", "AcsmPsIndx_bits"};
      this.AcsmPsIndx.configure(this, null, "");
      this.AcsmPsIndx.build();
      this.default_map.add_reg(this.AcsmPsIndx, `UVM_REG_ADDR_WIDTH'h1A9, "RW", 0);
		this.AcsmPsIndx_AcsmPsIndx = this.AcsmPsIndx.AcsmPsIndx;
      this.AcsmDynPtrCtrl = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmDynPtrCtrl::type_id::create("AcsmDynPtrCtrl",,get_full_name());
      if(this.AcsmDynPtrCtrl.has_coverage(UVM_CVR_ALL))
      	this.AcsmDynPtrCtrl.cg_bits.option.name = {get_name(), ".", "AcsmDynPtrCtrl_bits"};
      this.AcsmDynPtrCtrl.configure(this, null, "");
      this.AcsmDynPtrCtrl.build();
      this.default_map.add_reg(this.AcsmDynPtrCtrl, `UVM_REG_ADDR_WIDTH'h1AA, "RW", 0);
		this.AcsmDynPtrCtrl_AcsmDynPtrCtrl = this.AcsmDynPtrCtrl.AcsmDynPtrCtrl;
      this.FspState = ral_reg_DWC_DDRPHYA_PPGC0_p0_FspState::type_id::create("FspState",,get_full_name());
      if(this.FspState.has_coverage(UVM_CVR_ALL))
      	this.FspState.cg_bits.option.name = {get_name(), ".", "FspState_bits"};
      this.FspState.configure(this, null, "");
      this.FspState.build();
      this.default_map.add_reg(this.FspState, `UVM_REG_ADDR_WIDTH'h1EF, "RW", 0);
		this.FspState_DramFsp0xPhyPs = this.FspState.DramFsp0xPhyPs;
		this.DramFsp0xPhyPs = this.FspState.DramFsp0xPhyPs;
		this.FspState_DramFsp1xPhyPs = this.FspState.DramFsp1xPhyPs;
		this.DramFsp1xPhyPs = this.FspState.DramFsp1xPhyPs;
		this.FspState_DramFsp2xPhyPs = this.FspState.DramFsp2xPhyPs;
		this.DramFsp2xPhyPs = this.FspState.DramFsp2xPhyPs;
      this.AcsmMapTable0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable0::type_id::create("AcsmMapTable0",,get_full_name());
      if(this.AcsmMapTable0.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable0.cg_bits.option.name = {get_name(), ".", "AcsmMapTable0_bits"};
      this.AcsmMapTable0.configure(this, null, "");
      this.AcsmMapTable0.build();
      this.default_map.add_reg(this.AcsmMapTable0, `UVM_REG_ADDR_WIDTH'h200, "RW", 0);
		this.AcsmMapTable0_AcsmMapTableVal0 = this.AcsmMapTable0.AcsmMapTableVal0;
		this.AcsmMapTableVal0 = this.AcsmMapTable0.AcsmMapTableVal0;
		this.AcsmMapTable0_AcsmMapTableVal1 = this.AcsmMapTable0.AcsmMapTableVal1;
		this.AcsmMapTableVal1 = this.AcsmMapTable0.AcsmMapTableVal1;
      this.AcsmMapTable1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable1::type_id::create("AcsmMapTable1",,get_full_name());
      if(this.AcsmMapTable1.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable1.cg_bits.option.name = {get_name(), ".", "AcsmMapTable1_bits"};
      this.AcsmMapTable1.configure(this, null, "");
      this.AcsmMapTable1.build();
      this.default_map.add_reg(this.AcsmMapTable1, `UVM_REG_ADDR_WIDTH'h201, "RW", 0);
		this.AcsmMapTable1_AcsmMapTableVal2 = this.AcsmMapTable1.AcsmMapTableVal2;
		this.AcsmMapTableVal2 = this.AcsmMapTable1.AcsmMapTableVal2;
		this.AcsmMapTable1_AcsmMapTableVal3 = this.AcsmMapTable1.AcsmMapTableVal3;
		this.AcsmMapTableVal3 = this.AcsmMapTable1.AcsmMapTableVal3;
      this.AcsmMapTable2 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable2::type_id::create("AcsmMapTable2",,get_full_name());
      if(this.AcsmMapTable2.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable2.cg_bits.option.name = {get_name(), ".", "AcsmMapTable2_bits"};
      this.AcsmMapTable2.configure(this, null, "");
      this.AcsmMapTable2.build();
      this.default_map.add_reg(this.AcsmMapTable2, `UVM_REG_ADDR_WIDTH'h202, "RW", 0);
		this.AcsmMapTable2_AcsmMapTableVal4 = this.AcsmMapTable2.AcsmMapTableVal4;
		this.AcsmMapTableVal4 = this.AcsmMapTable2.AcsmMapTableVal4;
		this.AcsmMapTable2_AcsmMapTableVal5 = this.AcsmMapTable2.AcsmMapTableVal5;
		this.AcsmMapTableVal5 = this.AcsmMapTable2.AcsmMapTableVal5;
      this.AcsmMapTable3 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable3::type_id::create("AcsmMapTable3",,get_full_name());
      if(this.AcsmMapTable3.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable3.cg_bits.option.name = {get_name(), ".", "AcsmMapTable3_bits"};
      this.AcsmMapTable3.configure(this, null, "");
      this.AcsmMapTable3.build();
      this.default_map.add_reg(this.AcsmMapTable3, `UVM_REG_ADDR_WIDTH'h203, "RW", 0);
		this.AcsmMapTable3_AcsmMapTableVal6 = this.AcsmMapTable3.AcsmMapTableVal6;
		this.AcsmMapTableVal6 = this.AcsmMapTable3.AcsmMapTableVal6;
		this.AcsmMapTable3_AcsmMapTableVal7 = this.AcsmMapTable3.AcsmMapTableVal7;
		this.AcsmMapTableVal7 = this.AcsmMapTable3.AcsmMapTableVal7;
      this.AcsmMapTable4 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable4::type_id::create("AcsmMapTable4",,get_full_name());
      if(this.AcsmMapTable4.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable4.cg_bits.option.name = {get_name(), ".", "AcsmMapTable4_bits"};
      this.AcsmMapTable4.configure(this, null, "");
      this.AcsmMapTable4.build();
      this.default_map.add_reg(this.AcsmMapTable4, `UVM_REG_ADDR_WIDTH'h204, "RW", 0);
		this.AcsmMapTable4_AcsmMapTableVal8 = this.AcsmMapTable4.AcsmMapTableVal8;
		this.AcsmMapTableVal8 = this.AcsmMapTable4.AcsmMapTableVal8;
		this.AcsmMapTable4_AcsmMapTableVal9 = this.AcsmMapTable4.AcsmMapTableVal9;
		this.AcsmMapTableVal9 = this.AcsmMapTable4.AcsmMapTableVal9;
      this.AcsmMapTable5 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable5::type_id::create("AcsmMapTable5",,get_full_name());
      if(this.AcsmMapTable5.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable5.cg_bits.option.name = {get_name(), ".", "AcsmMapTable5_bits"};
      this.AcsmMapTable5.configure(this, null, "");
      this.AcsmMapTable5.build();
      this.default_map.add_reg(this.AcsmMapTable5, `UVM_REG_ADDR_WIDTH'h205, "RW", 0);
		this.AcsmMapTable5_AcsmMapTableVal10 = this.AcsmMapTable5.AcsmMapTableVal10;
		this.AcsmMapTableVal10 = this.AcsmMapTable5.AcsmMapTableVal10;
		this.AcsmMapTable5_AcsmMapTableVal11 = this.AcsmMapTable5.AcsmMapTableVal11;
		this.AcsmMapTableVal11 = this.AcsmMapTable5.AcsmMapTableVal11;
      this.AcsmMapTable6 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable6::type_id::create("AcsmMapTable6",,get_full_name());
      if(this.AcsmMapTable6.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable6.cg_bits.option.name = {get_name(), ".", "AcsmMapTable6_bits"};
      this.AcsmMapTable6.configure(this, null, "");
      this.AcsmMapTable6.build();
      this.default_map.add_reg(this.AcsmMapTable6, `UVM_REG_ADDR_WIDTH'h206, "RW", 0);
		this.AcsmMapTable6_AcsmMapTableVal12 = this.AcsmMapTable6.AcsmMapTableVal12;
		this.AcsmMapTableVal12 = this.AcsmMapTable6.AcsmMapTableVal12;
		this.AcsmMapTable6_AcsmMapTableVal13 = this.AcsmMapTable6.AcsmMapTableVal13;
		this.AcsmMapTableVal13 = this.AcsmMapTable6.AcsmMapTableVal13;
      this.AcsmMapTable7 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable7::type_id::create("AcsmMapTable7",,get_full_name());
      if(this.AcsmMapTable7.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable7.cg_bits.option.name = {get_name(), ".", "AcsmMapTable7_bits"};
      this.AcsmMapTable7.configure(this, null, "");
      this.AcsmMapTable7.build();
      this.default_map.add_reg(this.AcsmMapTable7, `UVM_REG_ADDR_WIDTH'h207, "RW", 0);
		this.AcsmMapTable7_AcsmMapTableVal14 = this.AcsmMapTable7.AcsmMapTableVal14;
		this.AcsmMapTableVal14 = this.AcsmMapTable7.AcsmMapTableVal14;
		this.AcsmMapTable7_AcsmMapTableVal15 = this.AcsmMapTable7.AcsmMapTableVal15;
		this.AcsmMapTableVal15 = this.AcsmMapTable7.AcsmMapTableVal15;
      this.AcsmMapTable8 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable8::type_id::create("AcsmMapTable8",,get_full_name());
      if(this.AcsmMapTable8.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable8.cg_bits.option.name = {get_name(), ".", "AcsmMapTable8_bits"};
      this.AcsmMapTable8.configure(this, null, "");
      this.AcsmMapTable8.build();
      this.default_map.add_reg(this.AcsmMapTable8, `UVM_REG_ADDR_WIDTH'h208, "RW", 0);
		this.AcsmMapTable8_AcsmMapTableVal16 = this.AcsmMapTable8.AcsmMapTableVal16;
		this.AcsmMapTableVal16 = this.AcsmMapTable8.AcsmMapTableVal16;
		this.AcsmMapTable8_AcsmMapTableVal17 = this.AcsmMapTable8.AcsmMapTableVal17;
		this.AcsmMapTableVal17 = this.AcsmMapTable8.AcsmMapTableVal17;
      this.AcsmMapTable9 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable9::type_id::create("AcsmMapTable9",,get_full_name());
      if(this.AcsmMapTable9.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable9.cg_bits.option.name = {get_name(), ".", "AcsmMapTable9_bits"};
      this.AcsmMapTable9.configure(this, null, "");
      this.AcsmMapTable9.build();
      this.default_map.add_reg(this.AcsmMapTable9, `UVM_REG_ADDR_WIDTH'h209, "RW", 0);
		this.AcsmMapTable9_AcsmMapTableVal18 = this.AcsmMapTable9.AcsmMapTableVal18;
		this.AcsmMapTableVal18 = this.AcsmMapTable9.AcsmMapTableVal18;
		this.AcsmMapTable9_AcsmMapTableVal19 = this.AcsmMapTable9.AcsmMapTableVal19;
		this.AcsmMapTableVal19 = this.AcsmMapTable9.AcsmMapTableVal19;
      this.AcsmMapTable10 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable10::type_id::create("AcsmMapTable10",,get_full_name());
      if(this.AcsmMapTable10.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable10.cg_bits.option.name = {get_name(), ".", "AcsmMapTable10_bits"};
      this.AcsmMapTable10.configure(this, null, "");
      this.AcsmMapTable10.build();
      this.default_map.add_reg(this.AcsmMapTable10, `UVM_REG_ADDR_WIDTH'h20A, "RW", 0);
		this.AcsmMapTable10_AcsmMapTableVal20 = this.AcsmMapTable10.AcsmMapTableVal20;
		this.AcsmMapTableVal20 = this.AcsmMapTable10.AcsmMapTableVal20;
		this.AcsmMapTable10_AcsmMapTableVal21 = this.AcsmMapTable10.AcsmMapTableVal21;
		this.AcsmMapTableVal21 = this.AcsmMapTable10.AcsmMapTableVal21;
      this.AcsmMapTable11 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable11::type_id::create("AcsmMapTable11",,get_full_name());
      if(this.AcsmMapTable11.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable11.cg_bits.option.name = {get_name(), ".", "AcsmMapTable11_bits"};
      this.AcsmMapTable11.configure(this, null, "");
      this.AcsmMapTable11.build();
      this.default_map.add_reg(this.AcsmMapTable11, `UVM_REG_ADDR_WIDTH'h20B, "RW", 0);
		this.AcsmMapTable11_AcsmMapTableVal22 = this.AcsmMapTable11.AcsmMapTableVal22;
		this.AcsmMapTableVal22 = this.AcsmMapTable11.AcsmMapTableVal22;
		this.AcsmMapTable11_AcsmMapTableVal23 = this.AcsmMapTable11.AcsmMapTableVal23;
		this.AcsmMapTableVal23 = this.AcsmMapTable11.AcsmMapTableVal23;
      this.AcsmMapTable12 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable12::type_id::create("AcsmMapTable12",,get_full_name());
      if(this.AcsmMapTable12.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable12.cg_bits.option.name = {get_name(), ".", "AcsmMapTable12_bits"};
      this.AcsmMapTable12.configure(this, null, "");
      this.AcsmMapTable12.build();
      this.default_map.add_reg(this.AcsmMapTable12, `UVM_REG_ADDR_WIDTH'h20C, "RW", 0);
		this.AcsmMapTable12_AcsmMapTableVal24 = this.AcsmMapTable12.AcsmMapTableVal24;
		this.AcsmMapTableVal24 = this.AcsmMapTable12.AcsmMapTableVal24;
		this.AcsmMapTable12_AcsmMapTableVal25 = this.AcsmMapTable12.AcsmMapTableVal25;
		this.AcsmMapTableVal25 = this.AcsmMapTable12.AcsmMapTableVal25;
      this.AcsmMapTable13 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable13::type_id::create("AcsmMapTable13",,get_full_name());
      if(this.AcsmMapTable13.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable13.cg_bits.option.name = {get_name(), ".", "AcsmMapTable13_bits"};
      this.AcsmMapTable13.configure(this, null, "");
      this.AcsmMapTable13.build();
      this.default_map.add_reg(this.AcsmMapTable13, `UVM_REG_ADDR_WIDTH'h20D, "RW", 0);
		this.AcsmMapTable13_AcsmMapTableVal26 = this.AcsmMapTable13.AcsmMapTableVal26;
		this.AcsmMapTableVal26 = this.AcsmMapTable13.AcsmMapTableVal26;
		this.AcsmMapTable13_AcsmMapTableVal27 = this.AcsmMapTable13.AcsmMapTableVal27;
		this.AcsmMapTableVal27 = this.AcsmMapTable13.AcsmMapTableVal27;
      this.AcsmMapTable14 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable14::type_id::create("AcsmMapTable14",,get_full_name());
      if(this.AcsmMapTable14.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable14.cg_bits.option.name = {get_name(), ".", "AcsmMapTable14_bits"};
      this.AcsmMapTable14.configure(this, null, "");
      this.AcsmMapTable14.build();
      this.default_map.add_reg(this.AcsmMapTable14, `UVM_REG_ADDR_WIDTH'h20E, "RW", 0);
		this.AcsmMapTable14_AcsmMapTableVal28 = this.AcsmMapTable14.AcsmMapTableVal28;
		this.AcsmMapTableVal28 = this.AcsmMapTable14.AcsmMapTableVal28;
		this.AcsmMapTable14_AcsmMapTableVal29 = this.AcsmMapTable14.AcsmMapTableVal29;
		this.AcsmMapTableVal29 = this.AcsmMapTable14.AcsmMapTableVal29;
      this.AcsmMapTable15 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable15::type_id::create("AcsmMapTable15",,get_full_name());
      if(this.AcsmMapTable15.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable15.cg_bits.option.name = {get_name(), ".", "AcsmMapTable15_bits"};
      this.AcsmMapTable15.configure(this, null, "");
      this.AcsmMapTable15.build();
      this.default_map.add_reg(this.AcsmMapTable15, `UVM_REG_ADDR_WIDTH'h20F, "RW", 0);
		this.AcsmMapTable15_AcsmMapTableVal30 = this.AcsmMapTable15.AcsmMapTableVal30;
		this.AcsmMapTableVal30 = this.AcsmMapTable15.AcsmMapTableVal30;
		this.AcsmMapTable15_AcsmMapTableVal31 = this.AcsmMapTable15.AcsmMapTableVal31;
		this.AcsmMapTableVal31 = this.AcsmMapTable15.AcsmMapTableVal31;
      this.AcsmMapTable16 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable16::type_id::create("AcsmMapTable16",,get_full_name());
      if(this.AcsmMapTable16.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable16.cg_bits.option.name = {get_name(), ".", "AcsmMapTable16_bits"};
      this.AcsmMapTable16.configure(this, null, "");
      this.AcsmMapTable16.build();
      this.default_map.add_reg(this.AcsmMapTable16, `UVM_REG_ADDR_WIDTH'h210, "RW", 0);
		this.AcsmMapTable16_AcsmMapTableVal32 = this.AcsmMapTable16.AcsmMapTableVal32;
		this.AcsmMapTableVal32 = this.AcsmMapTable16.AcsmMapTableVal32;
		this.AcsmMapTable16_AcsmMapTableVal33 = this.AcsmMapTable16.AcsmMapTableVal33;
		this.AcsmMapTableVal33 = this.AcsmMapTable16.AcsmMapTableVal33;
      this.AcsmMapTable17 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable17::type_id::create("AcsmMapTable17",,get_full_name());
      if(this.AcsmMapTable17.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable17.cg_bits.option.name = {get_name(), ".", "AcsmMapTable17_bits"};
      this.AcsmMapTable17.configure(this, null, "");
      this.AcsmMapTable17.build();
      this.default_map.add_reg(this.AcsmMapTable17, `UVM_REG_ADDR_WIDTH'h211, "RW", 0);
		this.AcsmMapTable17_AcsmMapTableVal34 = this.AcsmMapTable17.AcsmMapTableVal34;
		this.AcsmMapTableVal34 = this.AcsmMapTable17.AcsmMapTableVal34;
		this.AcsmMapTable17_AcsmMapTableVal35 = this.AcsmMapTable17.AcsmMapTableVal35;
		this.AcsmMapTableVal35 = this.AcsmMapTable17.AcsmMapTableVal35;
      this.AcsmMapTable18 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable18::type_id::create("AcsmMapTable18",,get_full_name());
      if(this.AcsmMapTable18.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable18.cg_bits.option.name = {get_name(), ".", "AcsmMapTable18_bits"};
      this.AcsmMapTable18.configure(this, null, "");
      this.AcsmMapTable18.build();
      this.default_map.add_reg(this.AcsmMapTable18, `UVM_REG_ADDR_WIDTH'h212, "RW", 0);
		this.AcsmMapTable18_AcsmMapTableVal36 = this.AcsmMapTable18.AcsmMapTableVal36;
		this.AcsmMapTableVal36 = this.AcsmMapTable18.AcsmMapTableVal36;
		this.AcsmMapTable18_AcsmMapTableVal37 = this.AcsmMapTable18.AcsmMapTableVal37;
		this.AcsmMapTableVal37 = this.AcsmMapTable18.AcsmMapTableVal37;
      this.AcsmMapTable19 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable19::type_id::create("AcsmMapTable19",,get_full_name());
      if(this.AcsmMapTable19.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable19.cg_bits.option.name = {get_name(), ".", "AcsmMapTable19_bits"};
      this.AcsmMapTable19.configure(this, null, "");
      this.AcsmMapTable19.build();
      this.default_map.add_reg(this.AcsmMapTable19, `UVM_REG_ADDR_WIDTH'h213, "RW", 0);
		this.AcsmMapTable19_AcsmMapTableVal38 = this.AcsmMapTable19.AcsmMapTableVal38;
		this.AcsmMapTableVal38 = this.AcsmMapTable19.AcsmMapTableVal38;
		this.AcsmMapTable19_AcsmMapTableVal39 = this.AcsmMapTable19.AcsmMapTableVal39;
		this.AcsmMapTableVal39 = this.AcsmMapTable19.AcsmMapTableVal39;
      this.AcsmMapTable20 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable20::type_id::create("AcsmMapTable20",,get_full_name());
      if(this.AcsmMapTable20.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable20.cg_bits.option.name = {get_name(), ".", "AcsmMapTable20_bits"};
      this.AcsmMapTable20.configure(this, null, "");
      this.AcsmMapTable20.build();
      this.default_map.add_reg(this.AcsmMapTable20, `UVM_REG_ADDR_WIDTH'h214, "RW", 0);
		this.AcsmMapTable20_AcsmMapTableVal40 = this.AcsmMapTable20.AcsmMapTableVal40;
		this.AcsmMapTableVal40 = this.AcsmMapTable20.AcsmMapTableVal40;
		this.AcsmMapTable20_AcsmMapTableVal41 = this.AcsmMapTable20.AcsmMapTableVal41;
		this.AcsmMapTableVal41 = this.AcsmMapTable20.AcsmMapTableVal41;
      this.AcsmMapTable21 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable21::type_id::create("AcsmMapTable21",,get_full_name());
      if(this.AcsmMapTable21.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable21.cg_bits.option.name = {get_name(), ".", "AcsmMapTable21_bits"};
      this.AcsmMapTable21.configure(this, null, "");
      this.AcsmMapTable21.build();
      this.default_map.add_reg(this.AcsmMapTable21, `UVM_REG_ADDR_WIDTH'h215, "RW", 0);
		this.AcsmMapTable21_AcsmMapTableVal42 = this.AcsmMapTable21.AcsmMapTableVal42;
		this.AcsmMapTableVal42 = this.AcsmMapTable21.AcsmMapTableVal42;
		this.AcsmMapTable21_AcsmMapTableVal43 = this.AcsmMapTable21.AcsmMapTableVal43;
		this.AcsmMapTableVal43 = this.AcsmMapTable21.AcsmMapTableVal43;
      this.AcsmMapTable22 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable22::type_id::create("AcsmMapTable22",,get_full_name());
      if(this.AcsmMapTable22.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable22.cg_bits.option.name = {get_name(), ".", "AcsmMapTable22_bits"};
      this.AcsmMapTable22.configure(this, null, "");
      this.AcsmMapTable22.build();
      this.default_map.add_reg(this.AcsmMapTable22, `UVM_REG_ADDR_WIDTH'h216, "RW", 0);
		this.AcsmMapTable22_AcsmMapTableVal44 = this.AcsmMapTable22.AcsmMapTableVal44;
		this.AcsmMapTableVal44 = this.AcsmMapTable22.AcsmMapTableVal44;
		this.AcsmMapTable22_AcsmMapTableVal45 = this.AcsmMapTable22.AcsmMapTableVal45;
		this.AcsmMapTableVal45 = this.AcsmMapTable22.AcsmMapTableVal45;
      this.AcsmMapTable23 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable23::type_id::create("AcsmMapTable23",,get_full_name());
      if(this.AcsmMapTable23.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable23.cg_bits.option.name = {get_name(), ".", "AcsmMapTable23_bits"};
      this.AcsmMapTable23.configure(this, null, "");
      this.AcsmMapTable23.build();
      this.default_map.add_reg(this.AcsmMapTable23, `UVM_REG_ADDR_WIDTH'h217, "RW", 0);
		this.AcsmMapTable23_AcsmMapTableVal46 = this.AcsmMapTable23.AcsmMapTableVal46;
		this.AcsmMapTableVal46 = this.AcsmMapTable23.AcsmMapTableVal46;
		this.AcsmMapTable23_AcsmMapTableVal47 = this.AcsmMapTable23.AcsmMapTableVal47;
		this.AcsmMapTableVal47 = this.AcsmMapTable23.AcsmMapTableVal47;
      this.AcsmMapTable24 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable24::type_id::create("AcsmMapTable24",,get_full_name());
      if(this.AcsmMapTable24.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable24.cg_bits.option.name = {get_name(), ".", "AcsmMapTable24_bits"};
      this.AcsmMapTable24.configure(this, null, "");
      this.AcsmMapTable24.build();
      this.default_map.add_reg(this.AcsmMapTable24, `UVM_REG_ADDR_WIDTH'h218, "RW", 0);
		this.AcsmMapTable24_AcsmMapTableVal48 = this.AcsmMapTable24.AcsmMapTableVal48;
		this.AcsmMapTableVal48 = this.AcsmMapTable24.AcsmMapTableVal48;
		this.AcsmMapTable24_AcsmMapTableVal49 = this.AcsmMapTable24.AcsmMapTableVal49;
		this.AcsmMapTableVal49 = this.AcsmMapTable24.AcsmMapTableVal49;
      this.AcsmMapTable25 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable25::type_id::create("AcsmMapTable25",,get_full_name());
      if(this.AcsmMapTable25.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable25.cg_bits.option.name = {get_name(), ".", "AcsmMapTable25_bits"};
      this.AcsmMapTable25.configure(this, null, "");
      this.AcsmMapTable25.build();
      this.default_map.add_reg(this.AcsmMapTable25, `UVM_REG_ADDR_WIDTH'h219, "RW", 0);
		this.AcsmMapTable25_AcsmMapTableVal50 = this.AcsmMapTable25.AcsmMapTableVal50;
		this.AcsmMapTableVal50 = this.AcsmMapTable25.AcsmMapTableVal50;
		this.AcsmMapTable25_AcsmMapTableVal51 = this.AcsmMapTable25.AcsmMapTableVal51;
		this.AcsmMapTableVal51 = this.AcsmMapTable25.AcsmMapTableVal51;
      this.AcsmMapTable26 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable26::type_id::create("AcsmMapTable26",,get_full_name());
      if(this.AcsmMapTable26.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable26.cg_bits.option.name = {get_name(), ".", "AcsmMapTable26_bits"};
      this.AcsmMapTable26.configure(this, null, "");
      this.AcsmMapTable26.build();
      this.default_map.add_reg(this.AcsmMapTable26, `UVM_REG_ADDR_WIDTH'h21A, "RW", 0);
		this.AcsmMapTable26_AcsmMapTableVal52 = this.AcsmMapTable26.AcsmMapTableVal52;
		this.AcsmMapTableVal52 = this.AcsmMapTable26.AcsmMapTableVal52;
		this.AcsmMapTable26_AcsmMapTableVal53 = this.AcsmMapTable26.AcsmMapTableVal53;
		this.AcsmMapTableVal53 = this.AcsmMapTable26.AcsmMapTableVal53;
      this.AcsmMapTable27 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable27::type_id::create("AcsmMapTable27",,get_full_name());
      if(this.AcsmMapTable27.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable27.cg_bits.option.name = {get_name(), ".", "AcsmMapTable27_bits"};
      this.AcsmMapTable27.configure(this, null, "");
      this.AcsmMapTable27.build();
      this.default_map.add_reg(this.AcsmMapTable27, `UVM_REG_ADDR_WIDTH'h21B, "RW", 0);
		this.AcsmMapTable27_AcsmMapTableVal54 = this.AcsmMapTable27.AcsmMapTableVal54;
		this.AcsmMapTableVal54 = this.AcsmMapTable27.AcsmMapTableVal54;
		this.AcsmMapTable27_AcsmMapTableVal55 = this.AcsmMapTable27.AcsmMapTableVal55;
		this.AcsmMapTableVal55 = this.AcsmMapTable27.AcsmMapTableVal55;
      this.AcsmMapTable28 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable28::type_id::create("AcsmMapTable28",,get_full_name());
      if(this.AcsmMapTable28.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable28.cg_bits.option.name = {get_name(), ".", "AcsmMapTable28_bits"};
      this.AcsmMapTable28.configure(this, null, "");
      this.AcsmMapTable28.build();
      this.default_map.add_reg(this.AcsmMapTable28, `UVM_REG_ADDR_WIDTH'h21C, "RW", 0);
		this.AcsmMapTable28_AcsmMapTableVal56 = this.AcsmMapTable28.AcsmMapTableVal56;
		this.AcsmMapTableVal56 = this.AcsmMapTable28.AcsmMapTableVal56;
		this.AcsmMapTable28_AcsmMapTableVal57 = this.AcsmMapTable28.AcsmMapTableVal57;
		this.AcsmMapTableVal57 = this.AcsmMapTable28.AcsmMapTableVal57;
      this.AcsmMapTable29 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable29::type_id::create("AcsmMapTable29",,get_full_name());
      if(this.AcsmMapTable29.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable29.cg_bits.option.name = {get_name(), ".", "AcsmMapTable29_bits"};
      this.AcsmMapTable29.configure(this, null, "");
      this.AcsmMapTable29.build();
      this.default_map.add_reg(this.AcsmMapTable29, `UVM_REG_ADDR_WIDTH'h21D, "RW", 0);
		this.AcsmMapTable29_AcsmMapTableVal58 = this.AcsmMapTable29.AcsmMapTableVal58;
		this.AcsmMapTableVal58 = this.AcsmMapTable29.AcsmMapTableVal58;
		this.AcsmMapTable29_AcsmMapTableVal59 = this.AcsmMapTable29.AcsmMapTableVal59;
		this.AcsmMapTableVal59 = this.AcsmMapTable29.AcsmMapTableVal59;
      this.AcsmMapTable30 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable30::type_id::create("AcsmMapTable30",,get_full_name());
      if(this.AcsmMapTable30.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable30.cg_bits.option.name = {get_name(), ".", "AcsmMapTable30_bits"};
      this.AcsmMapTable30.configure(this, null, "");
      this.AcsmMapTable30.build();
      this.default_map.add_reg(this.AcsmMapTable30, `UVM_REG_ADDR_WIDTH'h21E, "RW", 0);
		this.AcsmMapTable30_AcsmMapTableVal60 = this.AcsmMapTable30.AcsmMapTableVal60;
		this.AcsmMapTableVal60 = this.AcsmMapTable30.AcsmMapTableVal60;
		this.AcsmMapTable30_AcsmMapTableVal61 = this.AcsmMapTable30.AcsmMapTableVal61;
		this.AcsmMapTableVal61 = this.AcsmMapTable30.AcsmMapTableVal61;
      this.AcsmMapTable31 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable31::type_id::create("AcsmMapTable31",,get_full_name());
      if(this.AcsmMapTable31.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable31.cg_bits.option.name = {get_name(), ".", "AcsmMapTable31_bits"};
      this.AcsmMapTable31.configure(this, null, "");
      this.AcsmMapTable31.build();
      this.default_map.add_reg(this.AcsmMapTable31, `UVM_REG_ADDR_WIDTH'h21F, "RW", 0);
		this.AcsmMapTable31_AcsmMapTableVal62 = this.AcsmMapTable31.AcsmMapTableVal62;
		this.AcsmMapTableVal62 = this.AcsmMapTable31.AcsmMapTableVal62;
		this.AcsmMapTable31_AcsmMapTableVal63 = this.AcsmMapTable31.AcsmMapTableVal63;
		this.AcsmMapTableVal63 = this.AcsmMapTable31.AcsmMapTableVal63;
      this.AcsmMapTable32 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable32::type_id::create("AcsmMapTable32",,get_full_name());
      if(this.AcsmMapTable32.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable32.cg_bits.option.name = {get_name(), ".", "AcsmMapTable32_bits"};
      this.AcsmMapTable32.configure(this, null, "");
      this.AcsmMapTable32.build();
      this.default_map.add_reg(this.AcsmMapTable32, `UVM_REG_ADDR_WIDTH'h220, "RW", 0);
		this.AcsmMapTable32_AcsmMapTableVal64 = this.AcsmMapTable32.AcsmMapTableVal64;
		this.AcsmMapTableVal64 = this.AcsmMapTable32.AcsmMapTableVal64;
		this.AcsmMapTable32_AcsmMapTableVal65 = this.AcsmMapTable32.AcsmMapTableVal65;
		this.AcsmMapTableVal65 = this.AcsmMapTable32.AcsmMapTableVal65;
      this.AcsmMapTable33 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable33::type_id::create("AcsmMapTable33",,get_full_name());
      if(this.AcsmMapTable33.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable33.cg_bits.option.name = {get_name(), ".", "AcsmMapTable33_bits"};
      this.AcsmMapTable33.configure(this, null, "");
      this.AcsmMapTable33.build();
      this.default_map.add_reg(this.AcsmMapTable33, `UVM_REG_ADDR_WIDTH'h221, "RW", 0);
		this.AcsmMapTable33_AcsmMapTableVal66 = this.AcsmMapTable33.AcsmMapTableVal66;
		this.AcsmMapTableVal66 = this.AcsmMapTable33.AcsmMapTableVal66;
		this.AcsmMapTable33_AcsmMapTableVal67 = this.AcsmMapTable33.AcsmMapTableVal67;
		this.AcsmMapTableVal67 = this.AcsmMapTable33.AcsmMapTableVal67;
      this.AcsmMapTable34 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable34::type_id::create("AcsmMapTable34",,get_full_name());
      if(this.AcsmMapTable34.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable34.cg_bits.option.name = {get_name(), ".", "AcsmMapTable34_bits"};
      this.AcsmMapTable34.configure(this, null, "");
      this.AcsmMapTable34.build();
      this.default_map.add_reg(this.AcsmMapTable34, `UVM_REG_ADDR_WIDTH'h222, "RW", 0);
		this.AcsmMapTable34_AcsmMapTableVal68 = this.AcsmMapTable34.AcsmMapTableVal68;
		this.AcsmMapTableVal68 = this.AcsmMapTable34.AcsmMapTableVal68;
		this.AcsmMapTable34_AcsmMapTableVal69 = this.AcsmMapTable34.AcsmMapTableVal69;
		this.AcsmMapTableVal69 = this.AcsmMapTable34.AcsmMapTableVal69;
      this.AcsmMapTable35 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable35::type_id::create("AcsmMapTable35",,get_full_name());
      if(this.AcsmMapTable35.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable35.cg_bits.option.name = {get_name(), ".", "AcsmMapTable35_bits"};
      this.AcsmMapTable35.configure(this, null, "");
      this.AcsmMapTable35.build();
      this.default_map.add_reg(this.AcsmMapTable35, `UVM_REG_ADDR_WIDTH'h223, "RW", 0);
		this.AcsmMapTable35_AcsmMapTableVal70 = this.AcsmMapTable35.AcsmMapTableVal70;
		this.AcsmMapTableVal70 = this.AcsmMapTable35.AcsmMapTableVal70;
		this.AcsmMapTable35_AcsmMapTableVal71 = this.AcsmMapTable35.AcsmMapTableVal71;
		this.AcsmMapTableVal71 = this.AcsmMapTable35.AcsmMapTableVal71;
      this.AcsmMapTable36 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable36::type_id::create("AcsmMapTable36",,get_full_name());
      if(this.AcsmMapTable36.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable36.cg_bits.option.name = {get_name(), ".", "AcsmMapTable36_bits"};
      this.AcsmMapTable36.configure(this, null, "");
      this.AcsmMapTable36.build();
      this.default_map.add_reg(this.AcsmMapTable36, `UVM_REG_ADDR_WIDTH'h224, "RW", 0);
		this.AcsmMapTable36_AcsmMapTableVal72 = this.AcsmMapTable36.AcsmMapTableVal72;
		this.AcsmMapTableVal72 = this.AcsmMapTable36.AcsmMapTableVal72;
		this.AcsmMapTable36_AcsmMapTableVal73 = this.AcsmMapTable36.AcsmMapTableVal73;
		this.AcsmMapTableVal73 = this.AcsmMapTable36.AcsmMapTableVal73;
      this.AcsmMapTable37 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable37::type_id::create("AcsmMapTable37",,get_full_name());
      if(this.AcsmMapTable37.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable37.cg_bits.option.name = {get_name(), ".", "AcsmMapTable37_bits"};
      this.AcsmMapTable37.configure(this, null, "");
      this.AcsmMapTable37.build();
      this.default_map.add_reg(this.AcsmMapTable37, `UVM_REG_ADDR_WIDTH'h225, "RW", 0);
		this.AcsmMapTable37_AcsmMapTableVal74 = this.AcsmMapTable37.AcsmMapTableVal74;
		this.AcsmMapTableVal74 = this.AcsmMapTable37.AcsmMapTableVal74;
		this.AcsmMapTable37_AcsmMapTableVal75 = this.AcsmMapTable37.AcsmMapTableVal75;
		this.AcsmMapTableVal75 = this.AcsmMapTable37.AcsmMapTableVal75;
      this.AcsmMapTable38 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable38::type_id::create("AcsmMapTable38",,get_full_name());
      if(this.AcsmMapTable38.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable38.cg_bits.option.name = {get_name(), ".", "AcsmMapTable38_bits"};
      this.AcsmMapTable38.configure(this, null, "");
      this.AcsmMapTable38.build();
      this.default_map.add_reg(this.AcsmMapTable38, `UVM_REG_ADDR_WIDTH'h226, "RW", 0);
		this.AcsmMapTable38_AcsmMapTableVal76 = this.AcsmMapTable38.AcsmMapTableVal76;
		this.AcsmMapTableVal76 = this.AcsmMapTable38.AcsmMapTableVal76;
		this.AcsmMapTable38_AcsmMapTableVal77 = this.AcsmMapTable38.AcsmMapTableVal77;
		this.AcsmMapTableVal77 = this.AcsmMapTable38.AcsmMapTableVal77;
      this.AcsmMapTable39 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable39::type_id::create("AcsmMapTable39",,get_full_name());
      if(this.AcsmMapTable39.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable39.cg_bits.option.name = {get_name(), ".", "AcsmMapTable39_bits"};
      this.AcsmMapTable39.configure(this, null, "");
      this.AcsmMapTable39.build();
      this.default_map.add_reg(this.AcsmMapTable39, `UVM_REG_ADDR_WIDTH'h227, "RW", 0);
		this.AcsmMapTable39_AcsmMapTableVal78 = this.AcsmMapTable39.AcsmMapTableVal78;
		this.AcsmMapTableVal78 = this.AcsmMapTable39.AcsmMapTableVal78;
		this.AcsmMapTable39_AcsmMapTableVal79 = this.AcsmMapTable39.AcsmMapTableVal79;
		this.AcsmMapTableVal79 = this.AcsmMapTable39.AcsmMapTableVal79;
      this.AcsmMapTable40 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable40::type_id::create("AcsmMapTable40",,get_full_name());
      if(this.AcsmMapTable40.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable40.cg_bits.option.name = {get_name(), ".", "AcsmMapTable40_bits"};
      this.AcsmMapTable40.configure(this, null, "");
      this.AcsmMapTable40.build();
      this.default_map.add_reg(this.AcsmMapTable40, `UVM_REG_ADDR_WIDTH'h228, "RW", 0);
		this.AcsmMapTable40_AcsmMapTableVal80 = this.AcsmMapTable40.AcsmMapTableVal80;
		this.AcsmMapTableVal80 = this.AcsmMapTable40.AcsmMapTableVal80;
		this.AcsmMapTable40_AcsmMapTableVal81 = this.AcsmMapTable40.AcsmMapTableVal81;
		this.AcsmMapTableVal81 = this.AcsmMapTable40.AcsmMapTableVal81;
      this.AcsmMapTable41 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable41::type_id::create("AcsmMapTable41",,get_full_name());
      if(this.AcsmMapTable41.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable41.cg_bits.option.name = {get_name(), ".", "AcsmMapTable41_bits"};
      this.AcsmMapTable41.configure(this, null, "");
      this.AcsmMapTable41.build();
      this.default_map.add_reg(this.AcsmMapTable41, `UVM_REG_ADDR_WIDTH'h229, "RW", 0);
		this.AcsmMapTable41_AcsmMapTableVal82 = this.AcsmMapTable41.AcsmMapTableVal82;
		this.AcsmMapTableVal82 = this.AcsmMapTable41.AcsmMapTableVal82;
		this.AcsmMapTable41_AcsmMapTableVal83 = this.AcsmMapTable41.AcsmMapTableVal83;
		this.AcsmMapTableVal83 = this.AcsmMapTable41.AcsmMapTableVal83;
      this.AcsmMapTable42 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable42::type_id::create("AcsmMapTable42",,get_full_name());
      if(this.AcsmMapTable42.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable42.cg_bits.option.name = {get_name(), ".", "AcsmMapTable42_bits"};
      this.AcsmMapTable42.configure(this, null, "");
      this.AcsmMapTable42.build();
      this.default_map.add_reg(this.AcsmMapTable42, `UVM_REG_ADDR_WIDTH'h22A, "RW", 0);
		this.AcsmMapTable42_AcsmMapTableVal84 = this.AcsmMapTable42.AcsmMapTableVal84;
		this.AcsmMapTableVal84 = this.AcsmMapTable42.AcsmMapTableVal84;
		this.AcsmMapTable42_AcsmMapTableVal85 = this.AcsmMapTable42.AcsmMapTableVal85;
		this.AcsmMapTableVal85 = this.AcsmMapTable42.AcsmMapTableVal85;
      this.AcsmMapTable43 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable43::type_id::create("AcsmMapTable43",,get_full_name());
      if(this.AcsmMapTable43.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable43.cg_bits.option.name = {get_name(), ".", "AcsmMapTable43_bits"};
      this.AcsmMapTable43.configure(this, null, "");
      this.AcsmMapTable43.build();
      this.default_map.add_reg(this.AcsmMapTable43, `UVM_REG_ADDR_WIDTH'h22B, "RW", 0);
		this.AcsmMapTable43_AcsmMapTableVal86 = this.AcsmMapTable43.AcsmMapTableVal86;
		this.AcsmMapTableVal86 = this.AcsmMapTable43.AcsmMapTableVal86;
		this.AcsmMapTable43_AcsmMapTableVal87 = this.AcsmMapTable43.AcsmMapTableVal87;
		this.AcsmMapTableVal87 = this.AcsmMapTable43.AcsmMapTableVal87;
      this.AcsmMapTable44 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable44::type_id::create("AcsmMapTable44",,get_full_name());
      if(this.AcsmMapTable44.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable44.cg_bits.option.name = {get_name(), ".", "AcsmMapTable44_bits"};
      this.AcsmMapTable44.configure(this, null, "");
      this.AcsmMapTable44.build();
      this.default_map.add_reg(this.AcsmMapTable44, `UVM_REG_ADDR_WIDTH'h22C, "RW", 0);
		this.AcsmMapTable44_AcsmMapTableVal88 = this.AcsmMapTable44.AcsmMapTableVal88;
		this.AcsmMapTableVal88 = this.AcsmMapTable44.AcsmMapTableVal88;
		this.AcsmMapTable44_AcsmMapTableVal89 = this.AcsmMapTable44.AcsmMapTableVal89;
		this.AcsmMapTableVal89 = this.AcsmMapTable44.AcsmMapTableVal89;
      this.AcsmMapTable45 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable45::type_id::create("AcsmMapTable45",,get_full_name());
      if(this.AcsmMapTable45.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable45.cg_bits.option.name = {get_name(), ".", "AcsmMapTable45_bits"};
      this.AcsmMapTable45.configure(this, null, "");
      this.AcsmMapTable45.build();
      this.default_map.add_reg(this.AcsmMapTable45, `UVM_REG_ADDR_WIDTH'h22D, "RW", 0);
		this.AcsmMapTable45_AcsmMapTableVal90 = this.AcsmMapTable45.AcsmMapTableVal90;
		this.AcsmMapTableVal90 = this.AcsmMapTable45.AcsmMapTableVal90;
		this.AcsmMapTable45_AcsmMapTableVal91 = this.AcsmMapTable45.AcsmMapTableVal91;
		this.AcsmMapTableVal91 = this.AcsmMapTable45.AcsmMapTableVal91;
      this.AcsmMapTable46 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable46::type_id::create("AcsmMapTable46",,get_full_name());
      if(this.AcsmMapTable46.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable46.cg_bits.option.name = {get_name(), ".", "AcsmMapTable46_bits"};
      this.AcsmMapTable46.configure(this, null, "");
      this.AcsmMapTable46.build();
      this.default_map.add_reg(this.AcsmMapTable46, `UVM_REG_ADDR_WIDTH'h22E, "RW", 0);
		this.AcsmMapTable46_AcsmMapTableVal92 = this.AcsmMapTable46.AcsmMapTableVal92;
		this.AcsmMapTableVal92 = this.AcsmMapTable46.AcsmMapTableVal92;
		this.AcsmMapTable46_AcsmMapTableVal93 = this.AcsmMapTable46.AcsmMapTableVal93;
		this.AcsmMapTableVal93 = this.AcsmMapTable46.AcsmMapTableVal93;
      this.AcsmMapTable47 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable47::type_id::create("AcsmMapTable47",,get_full_name());
      if(this.AcsmMapTable47.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable47.cg_bits.option.name = {get_name(), ".", "AcsmMapTable47_bits"};
      this.AcsmMapTable47.configure(this, null, "");
      this.AcsmMapTable47.build();
      this.default_map.add_reg(this.AcsmMapTable47, `UVM_REG_ADDR_WIDTH'h22F, "RW", 0);
		this.AcsmMapTable47_AcsmMapTableVal94 = this.AcsmMapTable47.AcsmMapTableVal94;
		this.AcsmMapTableVal94 = this.AcsmMapTable47.AcsmMapTableVal94;
		this.AcsmMapTable47_AcsmMapTableVal95 = this.AcsmMapTable47.AcsmMapTableVal95;
		this.AcsmMapTableVal95 = this.AcsmMapTable47.AcsmMapTableVal95;
      this.AcsmMapTable48 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable48::type_id::create("AcsmMapTable48",,get_full_name());
      if(this.AcsmMapTable48.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable48.cg_bits.option.name = {get_name(), ".", "AcsmMapTable48_bits"};
      this.AcsmMapTable48.configure(this, null, "");
      this.AcsmMapTable48.build();
      this.default_map.add_reg(this.AcsmMapTable48, `UVM_REG_ADDR_WIDTH'h230, "RW", 0);
		this.AcsmMapTable48_AcsmMapTableVal96 = this.AcsmMapTable48.AcsmMapTableVal96;
		this.AcsmMapTableVal96 = this.AcsmMapTable48.AcsmMapTableVal96;
		this.AcsmMapTable48_AcsmMapTableVal97 = this.AcsmMapTable48.AcsmMapTableVal97;
		this.AcsmMapTableVal97 = this.AcsmMapTable48.AcsmMapTableVal97;
      this.AcsmMapTable49 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable49::type_id::create("AcsmMapTable49",,get_full_name());
      if(this.AcsmMapTable49.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable49.cg_bits.option.name = {get_name(), ".", "AcsmMapTable49_bits"};
      this.AcsmMapTable49.configure(this, null, "");
      this.AcsmMapTable49.build();
      this.default_map.add_reg(this.AcsmMapTable49, `UVM_REG_ADDR_WIDTH'h231, "RW", 0);
		this.AcsmMapTable49_AcsmMapTableVal98 = this.AcsmMapTable49.AcsmMapTableVal98;
		this.AcsmMapTableVal98 = this.AcsmMapTable49.AcsmMapTableVal98;
		this.AcsmMapTable49_AcsmMapTableVal99 = this.AcsmMapTable49.AcsmMapTableVal99;
		this.AcsmMapTableVal99 = this.AcsmMapTable49.AcsmMapTableVal99;
      this.AcsmMapTable50 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable50::type_id::create("AcsmMapTable50",,get_full_name());
      if(this.AcsmMapTable50.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable50.cg_bits.option.name = {get_name(), ".", "AcsmMapTable50_bits"};
      this.AcsmMapTable50.configure(this, null, "");
      this.AcsmMapTable50.build();
      this.default_map.add_reg(this.AcsmMapTable50, `UVM_REG_ADDR_WIDTH'h232, "RW", 0);
		this.AcsmMapTable50_AcsmMapTableVal100 = this.AcsmMapTable50.AcsmMapTableVal100;
		this.AcsmMapTableVal100 = this.AcsmMapTable50.AcsmMapTableVal100;
		this.AcsmMapTable50_AcsmMapTableVal101 = this.AcsmMapTable50.AcsmMapTableVal101;
		this.AcsmMapTableVal101 = this.AcsmMapTable50.AcsmMapTableVal101;
      this.AcsmMapTable51 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable51::type_id::create("AcsmMapTable51",,get_full_name());
      if(this.AcsmMapTable51.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable51.cg_bits.option.name = {get_name(), ".", "AcsmMapTable51_bits"};
      this.AcsmMapTable51.configure(this, null, "");
      this.AcsmMapTable51.build();
      this.default_map.add_reg(this.AcsmMapTable51, `UVM_REG_ADDR_WIDTH'h233, "RW", 0);
		this.AcsmMapTable51_AcsmMapTableVal102 = this.AcsmMapTable51.AcsmMapTableVal102;
		this.AcsmMapTableVal102 = this.AcsmMapTable51.AcsmMapTableVal102;
		this.AcsmMapTable51_AcsmMapTableVal103 = this.AcsmMapTable51.AcsmMapTableVal103;
		this.AcsmMapTableVal103 = this.AcsmMapTable51.AcsmMapTableVal103;
      this.AcsmMapTable52 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable52::type_id::create("AcsmMapTable52",,get_full_name());
      if(this.AcsmMapTable52.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable52.cg_bits.option.name = {get_name(), ".", "AcsmMapTable52_bits"};
      this.AcsmMapTable52.configure(this, null, "");
      this.AcsmMapTable52.build();
      this.default_map.add_reg(this.AcsmMapTable52, `UVM_REG_ADDR_WIDTH'h234, "RW", 0);
		this.AcsmMapTable52_AcsmMapTableVal104 = this.AcsmMapTable52.AcsmMapTableVal104;
		this.AcsmMapTableVal104 = this.AcsmMapTable52.AcsmMapTableVal104;
		this.AcsmMapTable52_AcsmMapTableVal105 = this.AcsmMapTable52.AcsmMapTableVal105;
		this.AcsmMapTableVal105 = this.AcsmMapTable52.AcsmMapTableVal105;
      this.AcsmMapTable53 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable53::type_id::create("AcsmMapTable53",,get_full_name());
      if(this.AcsmMapTable53.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable53.cg_bits.option.name = {get_name(), ".", "AcsmMapTable53_bits"};
      this.AcsmMapTable53.configure(this, null, "");
      this.AcsmMapTable53.build();
      this.default_map.add_reg(this.AcsmMapTable53, `UVM_REG_ADDR_WIDTH'h235, "RW", 0);
		this.AcsmMapTable53_AcsmMapTableVal106 = this.AcsmMapTable53.AcsmMapTableVal106;
		this.AcsmMapTableVal106 = this.AcsmMapTable53.AcsmMapTableVal106;
		this.AcsmMapTable53_AcsmMapTableVal107 = this.AcsmMapTable53.AcsmMapTableVal107;
		this.AcsmMapTableVal107 = this.AcsmMapTable53.AcsmMapTableVal107;
      this.AcsmMapTable54 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable54::type_id::create("AcsmMapTable54",,get_full_name());
      if(this.AcsmMapTable54.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable54.cg_bits.option.name = {get_name(), ".", "AcsmMapTable54_bits"};
      this.AcsmMapTable54.configure(this, null, "");
      this.AcsmMapTable54.build();
      this.default_map.add_reg(this.AcsmMapTable54, `UVM_REG_ADDR_WIDTH'h236, "RW", 0);
		this.AcsmMapTable54_AcsmMapTableVal108 = this.AcsmMapTable54.AcsmMapTableVal108;
		this.AcsmMapTableVal108 = this.AcsmMapTable54.AcsmMapTableVal108;
		this.AcsmMapTable54_AcsmMapTableVal109 = this.AcsmMapTable54.AcsmMapTableVal109;
		this.AcsmMapTableVal109 = this.AcsmMapTable54.AcsmMapTableVal109;
      this.AcsmMapTable55 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable55::type_id::create("AcsmMapTable55",,get_full_name());
      if(this.AcsmMapTable55.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable55.cg_bits.option.name = {get_name(), ".", "AcsmMapTable55_bits"};
      this.AcsmMapTable55.configure(this, null, "");
      this.AcsmMapTable55.build();
      this.default_map.add_reg(this.AcsmMapTable55, `UVM_REG_ADDR_WIDTH'h237, "RW", 0);
		this.AcsmMapTable55_AcsmMapTableVal110 = this.AcsmMapTable55.AcsmMapTableVal110;
		this.AcsmMapTableVal110 = this.AcsmMapTable55.AcsmMapTableVal110;
		this.AcsmMapTable55_AcsmMapTableVal111 = this.AcsmMapTable55.AcsmMapTableVal111;
		this.AcsmMapTableVal111 = this.AcsmMapTable55.AcsmMapTableVal111;
      this.AcsmMapTable56 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable56::type_id::create("AcsmMapTable56",,get_full_name());
      if(this.AcsmMapTable56.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable56.cg_bits.option.name = {get_name(), ".", "AcsmMapTable56_bits"};
      this.AcsmMapTable56.configure(this, null, "");
      this.AcsmMapTable56.build();
      this.default_map.add_reg(this.AcsmMapTable56, `UVM_REG_ADDR_WIDTH'h238, "RW", 0);
		this.AcsmMapTable56_AcsmMapTableVal112 = this.AcsmMapTable56.AcsmMapTableVal112;
		this.AcsmMapTableVal112 = this.AcsmMapTable56.AcsmMapTableVal112;
		this.AcsmMapTable56_AcsmMapTableVal113 = this.AcsmMapTable56.AcsmMapTableVal113;
		this.AcsmMapTableVal113 = this.AcsmMapTable56.AcsmMapTableVal113;
      this.AcsmMapTable57 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable57::type_id::create("AcsmMapTable57",,get_full_name());
      if(this.AcsmMapTable57.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable57.cg_bits.option.name = {get_name(), ".", "AcsmMapTable57_bits"};
      this.AcsmMapTable57.configure(this, null, "");
      this.AcsmMapTable57.build();
      this.default_map.add_reg(this.AcsmMapTable57, `UVM_REG_ADDR_WIDTH'h239, "RW", 0);
		this.AcsmMapTable57_AcsmMapTableVal114 = this.AcsmMapTable57.AcsmMapTableVal114;
		this.AcsmMapTableVal114 = this.AcsmMapTable57.AcsmMapTableVal114;
		this.AcsmMapTable57_AcsmMapTableVal115 = this.AcsmMapTable57.AcsmMapTableVal115;
		this.AcsmMapTableVal115 = this.AcsmMapTable57.AcsmMapTableVal115;
      this.AcsmMapTable58 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable58::type_id::create("AcsmMapTable58",,get_full_name());
      if(this.AcsmMapTable58.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable58.cg_bits.option.name = {get_name(), ".", "AcsmMapTable58_bits"};
      this.AcsmMapTable58.configure(this, null, "");
      this.AcsmMapTable58.build();
      this.default_map.add_reg(this.AcsmMapTable58, `UVM_REG_ADDR_WIDTH'h23A, "RW", 0);
		this.AcsmMapTable58_AcsmMapTableVal116 = this.AcsmMapTable58.AcsmMapTableVal116;
		this.AcsmMapTableVal116 = this.AcsmMapTable58.AcsmMapTableVal116;
		this.AcsmMapTable58_AcsmMapTableVal117 = this.AcsmMapTable58.AcsmMapTableVal117;
		this.AcsmMapTableVal117 = this.AcsmMapTable58.AcsmMapTableVal117;
      this.AcsmMapTable59 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable59::type_id::create("AcsmMapTable59",,get_full_name());
      if(this.AcsmMapTable59.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable59.cg_bits.option.name = {get_name(), ".", "AcsmMapTable59_bits"};
      this.AcsmMapTable59.configure(this, null, "");
      this.AcsmMapTable59.build();
      this.default_map.add_reg(this.AcsmMapTable59, `UVM_REG_ADDR_WIDTH'h23B, "RW", 0);
		this.AcsmMapTable59_AcsmMapTableVal118 = this.AcsmMapTable59.AcsmMapTableVal118;
		this.AcsmMapTableVal118 = this.AcsmMapTable59.AcsmMapTableVal118;
		this.AcsmMapTable59_AcsmMapTableVal119 = this.AcsmMapTable59.AcsmMapTableVal119;
		this.AcsmMapTableVal119 = this.AcsmMapTable59.AcsmMapTableVal119;
      this.AcsmMapTable60 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable60::type_id::create("AcsmMapTable60",,get_full_name());
      if(this.AcsmMapTable60.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable60.cg_bits.option.name = {get_name(), ".", "AcsmMapTable60_bits"};
      this.AcsmMapTable60.configure(this, null, "");
      this.AcsmMapTable60.build();
      this.default_map.add_reg(this.AcsmMapTable60, `UVM_REG_ADDR_WIDTH'h23C, "RW", 0);
		this.AcsmMapTable60_AcsmMapTableVal120 = this.AcsmMapTable60.AcsmMapTableVal120;
		this.AcsmMapTableVal120 = this.AcsmMapTable60.AcsmMapTableVal120;
		this.AcsmMapTable60_AcsmMapTableVal121 = this.AcsmMapTable60.AcsmMapTableVal121;
		this.AcsmMapTableVal121 = this.AcsmMapTable60.AcsmMapTableVal121;
      this.AcsmMapTable61 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable61::type_id::create("AcsmMapTable61",,get_full_name());
      if(this.AcsmMapTable61.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable61.cg_bits.option.name = {get_name(), ".", "AcsmMapTable61_bits"};
      this.AcsmMapTable61.configure(this, null, "");
      this.AcsmMapTable61.build();
      this.default_map.add_reg(this.AcsmMapTable61, `UVM_REG_ADDR_WIDTH'h23D, "RW", 0);
		this.AcsmMapTable61_AcsmMapTableVal122 = this.AcsmMapTable61.AcsmMapTableVal122;
		this.AcsmMapTableVal122 = this.AcsmMapTable61.AcsmMapTableVal122;
		this.AcsmMapTable61_AcsmMapTableVal123 = this.AcsmMapTable61.AcsmMapTableVal123;
		this.AcsmMapTableVal123 = this.AcsmMapTable61.AcsmMapTableVal123;
      this.AcsmMapTable62 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable62::type_id::create("AcsmMapTable62",,get_full_name());
      if(this.AcsmMapTable62.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable62.cg_bits.option.name = {get_name(), ".", "AcsmMapTable62_bits"};
      this.AcsmMapTable62.configure(this, null, "");
      this.AcsmMapTable62.build();
      this.default_map.add_reg(this.AcsmMapTable62, `UVM_REG_ADDR_WIDTH'h23E, "RW", 0);
		this.AcsmMapTable62_AcsmMapTableVal124 = this.AcsmMapTable62.AcsmMapTableVal124;
		this.AcsmMapTableVal124 = this.AcsmMapTable62.AcsmMapTableVal124;
		this.AcsmMapTable62_AcsmMapTableVal125 = this.AcsmMapTable62.AcsmMapTableVal125;
		this.AcsmMapTableVal125 = this.AcsmMapTable62.AcsmMapTableVal125;
      this.AcsmMapTable63 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmMapTable63::type_id::create("AcsmMapTable63",,get_full_name());
      if(this.AcsmMapTable63.has_coverage(UVM_CVR_ALL))
      	this.AcsmMapTable63.cg_bits.option.name = {get_name(), ".", "AcsmMapTable63_bits"};
      this.AcsmMapTable63.configure(this, null, "");
      this.AcsmMapTable63.build();
      this.default_map.add_reg(this.AcsmMapTable63, `UVM_REG_ADDR_WIDTH'h23F, "RW", 0);
		this.AcsmMapTable63_AcsmMapTableVal126 = this.AcsmMapTable63.AcsmMapTableVal126;
		this.AcsmMapTableVal126 = this.AcsmMapTable63.AcsmMapTableVal126;
		this.AcsmMapTable63_AcsmMapTableVal127 = this.AcsmMapTable63.AcsmMapTableVal127;
		this.AcsmMapTableVal127 = this.AcsmMapTable63.AcsmMapTableVal127;
      this.AcsmStartAddrXlatVal0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal0::type_id::create("AcsmStartAddrXlatVal0",,get_full_name());
      if(this.AcsmStartAddrXlatVal0.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal0.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal0_bits"};
      this.AcsmStartAddrXlatVal0.configure(this, null, "");
      this.AcsmStartAddrXlatVal0.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal0, `UVM_REG_ADDR_WIDTH'h324, "RW", 0);
		this.AcsmStartAddrXlatVal0_AcsmStartAddrXlatVal0 = this.AcsmStartAddrXlatVal0.AcsmStartAddrXlatVal0;
      this.AcsmStartAddrXlatVal1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal1::type_id::create("AcsmStartAddrXlatVal1",,get_full_name());
      if(this.AcsmStartAddrXlatVal1.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal1.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal1_bits"};
      this.AcsmStartAddrXlatVal1.configure(this, null, "");
      this.AcsmStartAddrXlatVal1.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal1, `UVM_REG_ADDR_WIDTH'h325, "RW", 0);
		this.AcsmStartAddrXlatVal1_AcsmStartAddrXlatVal1 = this.AcsmStartAddrXlatVal1.AcsmStartAddrXlatVal1;
      this.AcsmStartAddrXlatVal2 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal2::type_id::create("AcsmStartAddrXlatVal2",,get_full_name());
      if(this.AcsmStartAddrXlatVal2.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal2.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal2_bits"};
      this.AcsmStartAddrXlatVal2.configure(this, null, "");
      this.AcsmStartAddrXlatVal2.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal2, `UVM_REG_ADDR_WIDTH'h326, "RW", 0);
		this.AcsmStartAddrXlatVal2_AcsmStartAddrXlatVal2 = this.AcsmStartAddrXlatVal2.AcsmStartAddrXlatVal2;
      this.AcsmStartAddrXlatVal3 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal3::type_id::create("AcsmStartAddrXlatVal3",,get_full_name());
      if(this.AcsmStartAddrXlatVal3.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal3.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal3_bits"};
      this.AcsmStartAddrXlatVal3.configure(this, null, "");
      this.AcsmStartAddrXlatVal3.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal3, `UVM_REG_ADDR_WIDTH'h327, "RW", 0);
		this.AcsmStartAddrXlatVal3_AcsmStartAddrXlatVal3 = this.AcsmStartAddrXlatVal3.AcsmStartAddrXlatVal3;
      this.AcsmStartAddrXlatVal4 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal4::type_id::create("AcsmStartAddrXlatVal4",,get_full_name());
      if(this.AcsmStartAddrXlatVal4.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal4.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal4_bits"};
      this.AcsmStartAddrXlatVal4.configure(this, null, "");
      this.AcsmStartAddrXlatVal4.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal4, `UVM_REG_ADDR_WIDTH'h328, "RW", 0);
		this.AcsmStartAddrXlatVal4_AcsmStartAddrXlatVal4 = this.AcsmStartAddrXlatVal4.AcsmStartAddrXlatVal4;
      this.AcsmStartAddrXlatVal5 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal5::type_id::create("AcsmStartAddrXlatVal5",,get_full_name());
      if(this.AcsmStartAddrXlatVal5.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal5.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal5_bits"};
      this.AcsmStartAddrXlatVal5.configure(this, null, "");
      this.AcsmStartAddrXlatVal5.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal5, `UVM_REG_ADDR_WIDTH'h329, "RW", 0);
		this.AcsmStartAddrXlatVal5_AcsmStartAddrXlatVal5 = this.AcsmStartAddrXlatVal5.AcsmStartAddrXlatVal5;
      this.AcsmStartAddrXlatVal6 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal6::type_id::create("AcsmStartAddrXlatVal6",,get_full_name());
      if(this.AcsmStartAddrXlatVal6.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal6.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal6_bits"};
      this.AcsmStartAddrXlatVal6.configure(this, null, "");
      this.AcsmStartAddrXlatVal6.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal6, `UVM_REG_ADDR_WIDTH'h32A, "RW", 0);
		this.AcsmStartAddrXlatVal6_AcsmStartAddrXlatVal6 = this.AcsmStartAddrXlatVal6.AcsmStartAddrXlatVal6;
      this.AcsmStartAddrXlatVal7 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal7::type_id::create("AcsmStartAddrXlatVal7",,get_full_name());
      if(this.AcsmStartAddrXlatVal7.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal7.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal7_bits"};
      this.AcsmStartAddrXlatVal7.configure(this, null, "");
      this.AcsmStartAddrXlatVal7.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal7, `UVM_REG_ADDR_WIDTH'h32B, "RW", 0);
		this.AcsmStartAddrXlatVal7_AcsmStartAddrXlatVal7 = this.AcsmStartAddrXlatVal7.AcsmStartAddrXlatVal7;
      this.AcsmStartAddrXlatVal8 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal8::type_id::create("AcsmStartAddrXlatVal8",,get_full_name());
      if(this.AcsmStartAddrXlatVal8.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal8.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal8_bits"};
      this.AcsmStartAddrXlatVal8.configure(this, null, "");
      this.AcsmStartAddrXlatVal8.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal8, `UVM_REG_ADDR_WIDTH'h32C, "RW", 0);
		this.AcsmStartAddrXlatVal8_AcsmStartAddrXlatVal8 = this.AcsmStartAddrXlatVal8.AcsmStartAddrXlatVal8;
      this.AcsmStartAddrXlatVal9 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal9::type_id::create("AcsmStartAddrXlatVal9",,get_full_name());
      if(this.AcsmStartAddrXlatVal9.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal9.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal9_bits"};
      this.AcsmStartAddrXlatVal9.configure(this, null, "");
      this.AcsmStartAddrXlatVal9.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal9, `UVM_REG_ADDR_WIDTH'h32D, "RW", 0);
		this.AcsmStartAddrXlatVal9_AcsmStartAddrXlatVal9 = this.AcsmStartAddrXlatVal9.AcsmStartAddrXlatVal9;
      this.AcsmStartAddrXlatVal10 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal10::type_id::create("AcsmStartAddrXlatVal10",,get_full_name());
      if(this.AcsmStartAddrXlatVal10.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal10.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal10_bits"};
      this.AcsmStartAddrXlatVal10.configure(this, null, "");
      this.AcsmStartAddrXlatVal10.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal10, `UVM_REG_ADDR_WIDTH'h32E, "RW", 0);
		this.AcsmStartAddrXlatVal10_AcsmStartAddrXlatVal10 = this.AcsmStartAddrXlatVal10.AcsmStartAddrXlatVal10;
      this.AcsmStartAddrXlatVal11 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal11::type_id::create("AcsmStartAddrXlatVal11",,get_full_name());
      if(this.AcsmStartAddrXlatVal11.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal11.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal11_bits"};
      this.AcsmStartAddrXlatVal11.configure(this, null, "");
      this.AcsmStartAddrXlatVal11.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal11, `UVM_REG_ADDR_WIDTH'h32F, "RW", 0);
		this.AcsmStartAddrXlatVal11_AcsmStartAddrXlatVal11 = this.AcsmStartAddrXlatVal11.AcsmStartAddrXlatVal11;
      this.AcsmStartAddrXlatVal12 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal12::type_id::create("AcsmStartAddrXlatVal12",,get_full_name());
      if(this.AcsmStartAddrXlatVal12.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal12.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal12_bits"};
      this.AcsmStartAddrXlatVal12.configure(this, null, "");
      this.AcsmStartAddrXlatVal12.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal12, `UVM_REG_ADDR_WIDTH'h330, "RW", 0);
		this.AcsmStartAddrXlatVal12_AcsmStartAddrXlatVal12 = this.AcsmStartAddrXlatVal12.AcsmStartAddrXlatVal12;
      this.AcsmStartAddrXlatVal13 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal13::type_id::create("AcsmStartAddrXlatVal13",,get_full_name());
      if(this.AcsmStartAddrXlatVal13.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal13.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal13_bits"};
      this.AcsmStartAddrXlatVal13.configure(this, null, "");
      this.AcsmStartAddrXlatVal13.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal13, `UVM_REG_ADDR_WIDTH'h331, "RW", 0);
		this.AcsmStartAddrXlatVal13_AcsmStartAddrXlatVal13 = this.AcsmStartAddrXlatVal13.AcsmStartAddrXlatVal13;
      this.AcsmStartAddrXlatVal14 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal14::type_id::create("AcsmStartAddrXlatVal14",,get_full_name());
      if(this.AcsmStartAddrXlatVal14.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal14.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal14_bits"};
      this.AcsmStartAddrXlatVal14.configure(this, null, "");
      this.AcsmStartAddrXlatVal14.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal14, `UVM_REG_ADDR_WIDTH'h332, "RW", 0);
		this.AcsmStartAddrXlatVal14_AcsmStartAddrXlatVal14 = this.AcsmStartAddrXlatVal14.AcsmStartAddrXlatVal14;
      this.AcsmStartAddrXlatVal15 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal15::type_id::create("AcsmStartAddrXlatVal15",,get_full_name());
      if(this.AcsmStartAddrXlatVal15.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal15.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal15_bits"};
      this.AcsmStartAddrXlatVal15.configure(this, null, "");
      this.AcsmStartAddrXlatVal15.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal15, `UVM_REG_ADDR_WIDTH'h333, "RW", 0);
		this.AcsmStartAddrXlatVal15_AcsmStartAddrXlatVal15 = this.AcsmStartAddrXlatVal15.AcsmStartAddrXlatVal15;
      this.AcsmStartAddrXlatVal16 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal16::type_id::create("AcsmStartAddrXlatVal16",,get_full_name());
      if(this.AcsmStartAddrXlatVal16.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal16.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal16_bits"};
      this.AcsmStartAddrXlatVal16.configure(this, null, "");
      this.AcsmStartAddrXlatVal16.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal16, `UVM_REG_ADDR_WIDTH'h334, "RW", 0);
		this.AcsmStartAddrXlatVal16_AcsmStartAddrXlatVal16 = this.AcsmStartAddrXlatVal16.AcsmStartAddrXlatVal16;
      this.AcsmStartAddrXlatVal17 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal17::type_id::create("AcsmStartAddrXlatVal17",,get_full_name());
      if(this.AcsmStartAddrXlatVal17.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal17.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal17_bits"};
      this.AcsmStartAddrXlatVal17.configure(this, null, "");
      this.AcsmStartAddrXlatVal17.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal17, `UVM_REG_ADDR_WIDTH'h335, "RW", 0);
		this.AcsmStartAddrXlatVal17_AcsmStartAddrXlatVal17 = this.AcsmStartAddrXlatVal17.AcsmStartAddrXlatVal17;
      this.AcsmStartAddrXlatVal18 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal18::type_id::create("AcsmStartAddrXlatVal18",,get_full_name());
      if(this.AcsmStartAddrXlatVal18.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal18.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal18_bits"};
      this.AcsmStartAddrXlatVal18.configure(this, null, "");
      this.AcsmStartAddrXlatVal18.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal18, `UVM_REG_ADDR_WIDTH'h336, "RW", 0);
		this.AcsmStartAddrXlatVal18_AcsmStartAddrXlatVal18 = this.AcsmStartAddrXlatVal18.AcsmStartAddrXlatVal18;
      this.AcsmStartAddrXlatVal19 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal19::type_id::create("AcsmStartAddrXlatVal19",,get_full_name());
      if(this.AcsmStartAddrXlatVal19.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal19.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal19_bits"};
      this.AcsmStartAddrXlatVal19.configure(this, null, "");
      this.AcsmStartAddrXlatVal19.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal19, `UVM_REG_ADDR_WIDTH'h337, "RW", 0);
		this.AcsmStartAddrXlatVal19_AcsmStartAddrXlatVal19 = this.AcsmStartAddrXlatVal19.AcsmStartAddrXlatVal19;
      this.AcsmStartAddrXlatVal20 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal20::type_id::create("AcsmStartAddrXlatVal20",,get_full_name());
      if(this.AcsmStartAddrXlatVal20.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal20.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal20_bits"};
      this.AcsmStartAddrXlatVal20.configure(this, null, "");
      this.AcsmStartAddrXlatVal20.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal20, `UVM_REG_ADDR_WIDTH'h338, "RW", 0);
		this.AcsmStartAddrXlatVal20_AcsmStartAddrXlatVal20 = this.AcsmStartAddrXlatVal20.AcsmStartAddrXlatVal20;
      this.AcsmStartAddrXlatVal21 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal21::type_id::create("AcsmStartAddrXlatVal21",,get_full_name());
      if(this.AcsmStartAddrXlatVal21.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal21.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal21_bits"};
      this.AcsmStartAddrXlatVal21.configure(this, null, "");
      this.AcsmStartAddrXlatVal21.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal21, `UVM_REG_ADDR_WIDTH'h339, "RW", 0);
		this.AcsmStartAddrXlatVal21_AcsmStartAddrXlatVal21 = this.AcsmStartAddrXlatVal21.AcsmStartAddrXlatVal21;
      this.AcsmStartAddrXlatVal22 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal22::type_id::create("AcsmStartAddrXlatVal22",,get_full_name());
      if(this.AcsmStartAddrXlatVal22.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal22.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal22_bits"};
      this.AcsmStartAddrXlatVal22.configure(this, null, "");
      this.AcsmStartAddrXlatVal22.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal22, `UVM_REG_ADDR_WIDTH'h33A, "RW", 0);
		this.AcsmStartAddrXlatVal22_AcsmStartAddrXlatVal22 = this.AcsmStartAddrXlatVal22.AcsmStartAddrXlatVal22;
      this.AcsmStartAddrXlatVal23 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal23::type_id::create("AcsmStartAddrXlatVal23",,get_full_name());
      if(this.AcsmStartAddrXlatVal23.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal23.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal23_bits"};
      this.AcsmStartAddrXlatVal23.configure(this, null, "");
      this.AcsmStartAddrXlatVal23.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal23, `UVM_REG_ADDR_WIDTH'h33B, "RW", 0);
		this.AcsmStartAddrXlatVal23_AcsmStartAddrXlatVal23 = this.AcsmStartAddrXlatVal23.AcsmStartAddrXlatVal23;
      this.AcsmStartAddrXlatVal24 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal24::type_id::create("AcsmStartAddrXlatVal24",,get_full_name());
      if(this.AcsmStartAddrXlatVal24.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal24.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal24_bits"};
      this.AcsmStartAddrXlatVal24.configure(this, null, "");
      this.AcsmStartAddrXlatVal24.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal24, `UVM_REG_ADDR_WIDTH'h33C, "RW", 0);
		this.AcsmStartAddrXlatVal24_AcsmStartAddrXlatVal24 = this.AcsmStartAddrXlatVal24.AcsmStartAddrXlatVal24;
      this.AcsmStartAddrXlatVal25 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal25::type_id::create("AcsmStartAddrXlatVal25",,get_full_name());
      if(this.AcsmStartAddrXlatVal25.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal25.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal25_bits"};
      this.AcsmStartAddrXlatVal25.configure(this, null, "");
      this.AcsmStartAddrXlatVal25.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal25, `UVM_REG_ADDR_WIDTH'h33D, "RW", 0);
		this.AcsmStartAddrXlatVal25_AcsmStartAddrXlatVal25 = this.AcsmStartAddrXlatVal25.AcsmStartAddrXlatVal25;
      this.AcsmStartAddrXlatVal26 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal26::type_id::create("AcsmStartAddrXlatVal26",,get_full_name());
      if(this.AcsmStartAddrXlatVal26.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal26.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal26_bits"};
      this.AcsmStartAddrXlatVal26.configure(this, null, "");
      this.AcsmStartAddrXlatVal26.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal26, `UVM_REG_ADDR_WIDTH'h33E, "RW", 0);
		this.AcsmStartAddrXlatVal26_AcsmStartAddrXlatVal26 = this.AcsmStartAddrXlatVal26.AcsmStartAddrXlatVal26;
      this.AcsmStartAddrXlatVal27 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal27::type_id::create("AcsmStartAddrXlatVal27",,get_full_name());
      if(this.AcsmStartAddrXlatVal27.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal27.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal27_bits"};
      this.AcsmStartAddrXlatVal27.configure(this, null, "");
      this.AcsmStartAddrXlatVal27.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal27, `UVM_REG_ADDR_WIDTH'h33F, "RW", 0);
		this.AcsmStartAddrXlatVal27_AcsmStartAddrXlatVal27 = this.AcsmStartAddrXlatVal27.AcsmStartAddrXlatVal27;
      this.AcsmStartAddrXlatVal28 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal28::type_id::create("AcsmStartAddrXlatVal28",,get_full_name());
      if(this.AcsmStartAddrXlatVal28.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal28.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal28_bits"};
      this.AcsmStartAddrXlatVal28.configure(this, null, "");
      this.AcsmStartAddrXlatVal28.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal28, `UVM_REG_ADDR_WIDTH'h340, "RW", 0);
		this.AcsmStartAddrXlatVal28_AcsmStartAddrXlatVal28 = this.AcsmStartAddrXlatVal28.AcsmStartAddrXlatVal28;
      this.AcsmStartAddrXlatVal29 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal29::type_id::create("AcsmStartAddrXlatVal29",,get_full_name());
      if(this.AcsmStartAddrXlatVal29.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal29.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal29_bits"};
      this.AcsmStartAddrXlatVal29.configure(this, null, "");
      this.AcsmStartAddrXlatVal29.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal29, `UVM_REG_ADDR_WIDTH'h341, "RW", 0);
		this.AcsmStartAddrXlatVal29_AcsmStartAddrXlatVal29 = this.AcsmStartAddrXlatVal29.AcsmStartAddrXlatVal29;
      this.AcsmStartAddrXlatVal30 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal30::type_id::create("AcsmStartAddrXlatVal30",,get_full_name());
      if(this.AcsmStartAddrXlatVal30.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal30.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal30_bits"};
      this.AcsmStartAddrXlatVal30.configure(this, null, "");
      this.AcsmStartAddrXlatVal30.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal30, `UVM_REG_ADDR_WIDTH'h342, "RW", 0);
		this.AcsmStartAddrXlatVal30_AcsmStartAddrXlatVal30 = this.AcsmStartAddrXlatVal30.AcsmStartAddrXlatVal30;
      this.AcsmStartAddrXlatVal31 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal31::type_id::create("AcsmStartAddrXlatVal31",,get_full_name());
      if(this.AcsmStartAddrXlatVal31.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal31.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal31_bits"};
      this.AcsmStartAddrXlatVal31.configure(this, null, "");
      this.AcsmStartAddrXlatVal31.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal31, `UVM_REG_ADDR_WIDTH'h343, "RW", 0);
		this.AcsmStartAddrXlatVal31_AcsmStartAddrXlatVal31 = this.AcsmStartAddrXlatVal31.AcsmStartAddrXlatVal31;
      this.AcsmStartAddrXlatVal32 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal32::type_id::create("AcsmStartAddrXlatVal32",,get_full_name());
      if(this.AcsmStartAddrXlatVal32.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal32.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal32_bits"};
      this.AcsmStartAddrXlatVal32.configure(this, null, "");
      this.AcsmStartAddrXlatVal32.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal32, `UVM_REG_ADDR_WIDTH'h344, "RW", 0);
		this.AcsmStartAddrXlatVal32_AcsmStartAddrXlatVal32 = this.AcsmStartAddrXlatVal32.AcsmStartAddrXlatVal32;
      this.AcsmStartAddrXlatVal33 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal33::type_id::create("AcsmStartAddrXlatVal33",,get_full_name());
      if(this.AcsmStartAddrXlatVal33.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal33.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal33_bits"};
      this.AcsmStartAddrXlatVal33.configure(this, null, "");
      this.AcsmStartAddrXlatVal33.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal33, `UVM_REG_ADDR_WIDTH'h345, "RW", 0);
		this.AcsmStartAddrXlatVal33_AcsmStartAddrXlatVal33 = this.AcsmStartAddrXlatVal33.AcsmStartAddrXlatVal33;
      this.AcsmStartAddrXlatVal34 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal34::type_id::create("AcsmStartAddrXlatVal34",,get_full_name());
      if(this.AcsmStartAddrXlatVal34.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal34.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal34_bits"};
      this.AcsmStartAddrXlatVal34.configure(this, null, "");
      this.AcsmStartAddrXlatVal34.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal34, `UVM_REG_ADDR_WIDTH'h346, "RW", 0);
		this.AcsmStartAddrXlatVal34_AcsmStartAddrXlatVal34 = this.AcsmStartAddrXlatVal34.AcsmStartAddrXlatVal34;
      this.AcsmStartAddrXlatVal35 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal35::type_id::create("AcsmStartAddrXlatVal35",,get_full_name());
      if(this.AcsmStartAddrXlatVal35.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal35.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal35_bits"};
      this.AcsmStartAddrXlatVal35.configure(this, null, "");
      this.AcsmStartAddrXlatVal35.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal35, `UVM_REG_ADDR_WIDTH'h347, "RW", 0);
		this.AcsmStartAddrXlatVal35_AcsmStartAddrXlatVal35 = this.AcsmStartAddrXlatVal35.AcsmStartAddrXlatVal35;
      this.AcsmStartAddrXlatVal36 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal36::type_id::create("AcsmStartAddrXlatVal36",,get_full_name());
      if(this.AcsmStartAddrXlatVal36.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal36.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal36_bits"};
      this.AcsmStartAddrXlatVal36.configure(this, null, "");
      this.AcsmStartAddrXlatVal36.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal36, `UVM_REG_ADDR_WIDTH'h348, "RW", 0);
		this.AcsmStartAddrXlatVal36_AcsmStartAddrXlatVal36 = this.AcsmStartAddrXlatVal36.AcsmStartAddrXlatVal36;
      this.AcsmStartAddrXlatVal37 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal37::type_id::create("AcsmStartAddrXlatVal37",,get_full_name());
      if(this.AcsmStartAddrXlatVal37.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal37.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal37_bits"};
      this.AcsmStartAddrXlatVal37.configure(this, null, "");
      this.AcsmStartAddrXlatVal37.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal37, `UVM_REG_ADDR_WIDTH'h349, "RW", 0);
		this.AcsmStartAddrXlatVal37_AcsmStartAddrXlatVal37 = this.AcsmStartAddrXlatVal37.AcsmStartAddrXlatVal37;
      this.AcsmStartAddrXlatVal38 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal38::type_id::create("AcsmStartAddrXlatVal38",,get_full_name());
      if(this.AcsmStartAddrXlatVal38.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal38.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal38_bits"};
      this.AcsmStartAddrXlatVal38.configure(this, null, "");
      this.AcsmStartAddrXlatVal38.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal38, `UVM_REG_ADDR_WIDTH'h34A, "RW", 0);
		this.AcsmStartAddrXlatVal38_AcsmStartAddrXlatVal38 = this.AcsmStartAddrXlatVal38.AcsmStartAddrXlatVal38;
      this.AcsmStartAddrXlatVal39 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal39::type_id::create("AcsmStartAddrXlatVal39",,get_full_name());
      if(this.AcsmStartAddrXlatVal39.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal39.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal39_bits"};
      this.AcsmStartAddrXlatVal39.configure(this, null, "");
      this.AcsmStartAddrXlatVal39.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal39, `UVM_REG_ADDR_WIDTH'h34B, "RW", 0);
		this.AcsmStartAddrXlatVal39_AcsmStartAddrXlatVal39 = this.AcsmStartAddrXlatVal39.AcsmStartAddrXlatVal39;
      this.AcsmStartAddrXlatVal40 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal40::type_id::create("AcsmStartAddrXlatVal40",,get_full_name());
      if(this.AcsmStartAddrXlatVal40.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal40.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal40_bits"};
      this.AcsmStartAddrXlatVal40.configure(this, null, "");
      this.AcsmStartAddrXlatVal40.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal40, `UVM_REG_ADDR_WIDTH'h34C, "RW", 0);
		this.AcsmStartAddrXlatVal40_AcsmStartAddrXlatVal40 = this.AcsmStartAddrXlatVal40.AcsmStartAddrXlatVal40;
      this.AcsmStartAddrXlatVal41 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal41::type_id::create("AcsmStartAddrXlatVal41",,get_full_name());
      if(this.AcsmStartAddrXlatVal41.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal41.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal41_bits"};
      this.AcsmStartAddrXlatVal41.configure(this, null, "");
      this.AcsmStartAddrXlatVal41.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal41, `UVM_REG_ADDR_WIDTH'h34D, "RW", 0);
		this.AcsmStartAddrXlatVal41_AcsmStartAddrXlatVal41 = this.AcsmStartAddrXlatVal41.AcsmStartAddrXlatVal41;
      this.AcsmStartAddrXlatVal42 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal42::type_id::create("AcsmStartAddrXlatVal42",,get_full_name());
      if(this.AcsmStartAddrXlatVal42.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal42.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal42_bits"};
      this.AcsmStartAddrXlatVal42.configure(this, null, "");
      this.AcsmStartAddrXlatVal42.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal42, `UVM_REG_ADDR_WIDTH'h34E, "RW", 0);
		this.AcsmStartAddrXlatVal42_AcsmStartAddrXlatVal42 = this.AcsmStartAddrXlatVal42.AcsmStartAddrXlatVal42;
      this.AcsmStartAddrXlatVal43 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal43::type_id::create("AcsmStartAddrXlatVal43",,get_full_name());
      if(this.AcsmStartAddrXlatVal43.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal43.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal43_bits"};
      this.AcsmStartAddrXlatVal43.configure(this, null, "");
      this.AcsmStartAddrXlatVal43.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal43, `UVM_REG_ADDR_WIDTH'h34F, "RW", 0);
		this.AcsmStartAddrXlatVal43_AcsmStartAddrXlatVal43 = this.AcsmStartAddrXlatVal43.AcsmStartAddrXlatVal43;
      this.AcsmStartAddrXlatVal44 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal44::type_id::create("AcsmStartAddrXlatVal44",,get_full_name());
      if(this.AcsmStartAddrXlatVal44.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal44.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal44_bits"};
      this.AcsmStartAddrXlatVal44.configure(this, null, "");
      this.AcsmStartAddrXlatVal44.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal44, `UVM_REG_ADDR_WIDTH'h350, "RW", 0);
		this.AcsmStartAddrXlatVal44_AcsmStartAddrXlatVal44 = this.AcsmStartAddrXlatVal44.AcsmStartAddrXlatVal44;
      this.AcsmStartAddrXlatVal45 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal45::type_id::create("AcsmStartAddrXlatVal45",,get_full_name());
      if(this.AcsmStartAddrXlatVal45.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal45.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal45_bits"};
      this.AcsmStartAddrXlatVal45.configure(this, null, "");
      this.AcsmStartAddrXlatVal45.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal45, `UVM_REG_ADDR_WIDTH'h351, "RW", 0);
		this.AcsmStartAddrXlatVal45_AcsmStartAddrXlatVal45 = this.AcsmStartAddrXlatVal45.AcsmStartAddrXlatVal45;
      this.AcsmStartAddrXlatVal46 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal46::type_id::create("AcsmStartAddrXlatVal46",,get_full_name());
      if(this.AcsmStartAddrXlatVal46.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal46.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal46_bits"};
      this.AcsmStartAddrXlatVal46.configure(this, null, "");
      this.AcsmStartAddrXlatVal46.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal46, `UVM_REG_ADDR_WIDTH'h352, "RW", 0);
		this.AcsmStartAddrXlatVal46_AcsmStartAddrXlatVal46 = this.AcsmStartAddrXlatVal46.AcsmStartAddrXlatVal46;
      this.AcsmStartAddrXlatVal47 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal47::type_id::create("AcsmStartAddrXlatVal47",,get_full_name());
      if(this.AcsmStartAddrXlatVal47.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal47.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal47_bits"};
      this.AcsmStartAddrXlatVal47.configure(this, null, "");
      this.AcsmStartAddrXlatVal47.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal47, `UVM_REG_ADDR_WIDTH'h353, "RW", 0);
		this.AcsmStartAddrXlatVal47_AcsmStartAddrXlatVal47 = this.AcsmStartAddrXlatVal47.AcsmStartAddrXlatVal47;
      this.AcsmStartAddrXlatVal48 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal48::type_id::create("AcsmStartAddrXlatVal48",,get_full_name());
      if(this.AcsmStartAddrXlatVal48.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal48.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal48_bits"};
      this.AcsmStartAddrXlatVal48.configure(this, null, "");
      this.AcsmStartAddrXlatVal48.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal48, `UVM_REG_ADDR_WIDTH'h354, "RW", 0);
		this.AcsmStartAddrXlatVal48_AcsmStartAddrXlatVal48 = this.AcsmStartAddrXlatVal48.AcsmStartAddrXlatVal48;
      this.AcsmStartAddrXlatVal49 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal49::type_id::create("AcsmStartAddrXlatVal49",,get_full_name());
      if(this.AcsmStartAddrXlatVal49.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal49.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal49_bits"};
      this.AcsmStartAddrXlatVal49.configure(this, null, "");
      this.AcsmStartAddrXlatVal49.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal49, `UVM_REG_ADDR_WIDTH'h355, "RW", 0);
		this.AcsmStartAddrXlatVal49_AcsmStartAddrXlatVal49 = this.AcsmStartAddrXlatVal49.AcsmStartAddrXlatVal49;
      this.AcsmStartAddrXlatVal50 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal50::type_id::create("AcsmStartAddrXlatVal50",,get_full_name());
      if(this.AcsmStartAddrXlatVal50.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal50.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal50_bits"};
      this.AcsmStartAddrXlatVal50.configure(this, null, "");
      this.AcsmStartAddrXlatVal50.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal50, `UVM_REG_ADDR_WIDTH'h356, "RW", 0);
		this.AcsmStartAddrXlatVal50_AcsmStartAddrXlatVal50 = this.AcsmStartAddrXlatVal50.AcsmStartAddrXlatVal50;
      this.AcsmStartAddrXlatVal51 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal51::type_id::create("AcsmStartAddrXlatVal51",,get_full_name());
      if(this.AcsmStartAddrXlatVal51.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal51.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal51_bits"};
      this.AcsmStartAddrXlatVal51.configure(this, null, "");
      this.AcsmStartAddrXlatVal51.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal51, `UVM_REG_ADDR_WIDTH'h357, "RW", 0);
		this.AcsmStartAddrXlatVal51_AcsmStartAddrXlatVal51 = this.AcsmStartAddrXlatVal51.AcsmStartAddrXlatVal51;
      this.AcsmStartAddrXlatVal52 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal52::type_id::create("AcsmStartAddrXlatVal52",,get_full_name());
      if(this.AcsmStartAddrXlatVal52.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal52.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal52_bits"};
      this.AcsmStartAddrXlatVal52.configure(this, null, "");
      this.AcsmStartAddrXlatVal52.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal52, `UVM_REG_ADDR_WIDTH'h358, "RW", 0);
		this.AcsmStartAddrXlatVal52_AcsmStartAddrXlatVal52 = this.AcsmStartAddrXlatVal52.AcsmStartAddrXlatVal52;
      this.AcsmStartAddrXlatVal53 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal53::type_id::create("AcsmStartAddrXlatVal53",,get_full_name());
      if(this.AcsmStartAddrXlatVal53.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal53.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal53_bits"};
      this.AcsmStartAddrXlatVal53.configure(this, null, "");
      this.AcsmStartAddrXlatVal53.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal53, `UVM_REG_ADDR_WIDTH'h359, "RW", 0);
		this.AcsmStartAddrXlatVal53_AcsmStartAddrXlatVal53 = this.AcsmStartAddrXlatVal53.AcsmStartAddrXlatVal53;
      this.AcsmStartAddrXlatVal54 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal54::type_id::create("AcsmStartAddrXlatVal54",,get_full_name());
      if(this.AcsmStartAddrXlatVal54.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal54.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal54_bits"};
      this.AcsmStartAddrXlatVal54.configure(this, null, "");
      this.AcsmStartAddrXlatVal54.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal54, `UVM_REG_ADDR_WIDTH'h35A, "RW", 0);
		this.AcsmStartAddrXlatVal54_AcsmStartAddrXlatVal54 = this.AcsmStartAddrXlatVal54.AcsmStartAddrXlatVal54;
      this.AcsmStartAddrXlatVal55 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal55::type_id::create("AcsmStartAddrXlatVal55",,get_full_name());
      if(this.AcsmStartAddrXlatVal55.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal55.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal55_bits"};
      this.AcsmStartAddrXlatVal55.configure(this, null, "");
      this.AcsmStartAddrXlatVal55.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal55, `UVM_REG_ADDR_WIDTH'h35B, "RW", 0);
		this.AcsmStartAddrXlatVal55_AcsmStartAddrXlatVal55 = this.AcsmStartAddrXlatVal55.AcsmStartAddrXlatVal55;
      this.AcsmStartAddrXlatVal56 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal56::type_id::create("AcsmStartAddrXlatVal56",,get_full_name());
      if(this.AcsmStartAddrXlatVal56.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal56.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal56_bits"};
      this.AcsmStartAddrXlatVal56.configure(this, null, "");
      this.AcsmStartAddrXlatVal56.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal56, `UVM_REG_ADDR_WIDTH'h35C, "RW", 0);
		this.AcsmStartAddrXlatVal56_AcsmStartAddrXlatVal56 = this.AcsmStartAddrXlatVal56.AcsmStartAddrXlatVal56;
      this.AcsmStartAddrXlatVal57 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal57::type_id::create("AcsmStartAddrXlatVal57",,get_full_name());
      if(this.AcsmStartAddrXlatVal57.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal57.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal57_bits"};
      this.AcsmStartAddrXlatVal57.configure(this, null, "");
      this.AcsmStartAddrXlatVal57.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal57, `UVM_REG_ADDR_WIDTH'h35D, "RW", 0);
		this.AcsmStartAddrXlatVal57_AcsmStartAddrXlatVal57 = this.AcsmStartAddrXlatVal57.AcsmStartAddrXlatVal57;
      this.AcsmStartAddrXlatVal58 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal58::type_id::create("AcsmStartAddrXlatVal58",,get_full_name());
      if(this.AcsmStartAddrXlatVal58.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal58.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal58_bits"};
      this.AcsmStartAddrXlatVal58.configure(this, null, "");
      this.AcsmStartAddrXlatVal58.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal58, `UVM_REG_ADDR_WIDTH'h35E, "RW", 0);
		this.AcsmStartAddrXlatVal58_AcsmStartAddrXlatVal58 = this.AcsmStartAddrXlatVal58.AcsmStartAddrXlatVal58;
      this.AcsmStartAddrXlatVal59 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal59::type_id::create("AcsmStartAddrXlatVal59",,get_full_name());
      if(this.AcsmStartAddrXlatVal59.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal59.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal59_bits"};
      this.AcsmStartAddrXlatVal59.configure(this, null, "");
      this.AcsmStartAddrXlatVal59.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal59, `UVM_REG_ADDR_WIDTH'h35F, "RW", 0);
		this.AcsmStartAddrXlatVal59_AcsmStartAddrXlatVal59 = this.AcsmStartAddrXlatVal59.AcsmStartAddrXlatVal59;
      this.AcsmStartAddrXlatVal60 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal60::type_id::create("AcsmStartAddrXlatVal60",,get_full_name());
      if(this.AcsmStartAddrXlatVal60.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal60.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal60_bits"};
      this.AcsmStartAddrXlatVal60.configure(this, null, "");
      this.AcsmStartAddrXlatVal60.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal60, `UVM_REG_ADDR_WIDTH'h360, "RW", 0);
		this.AcsmStartAddrXlatVal60_AcsmStartAddrXlatVal60 = this.AcsmStartAddrXlatVal60.AcsmStartAddrXlatVal60;
      this.AcsmStartAddrXlatVal61 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal61::type_id::create("AcsmStartAddrXlatVal61",,get_full_name());
      if(this.AcsmStartAddrXlatVal61.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal61.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal61_bits"};
      this.AcsmStartAddrXlatVal61.configure(this, null, "");
      this.AcsmStartAddrXlatVal61.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal61, `UVM_REG_ADDR_WIDTH'h361, "RW", 0);
		this.AcsmStartAddrXlatVal61_AcsmStartAddrXlatVal61 = this.AcsmStartAddrXlatVal61.AcsmStartAddrXlatVal61;
      this.AcsmStartAddrXlatVal62 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal62::type_id::create("AcsmStartAddrXlatVal62",,get_full_name());
      if(this.AcsmStartAddrXlatVal62.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal62.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal62_bits"};
      this.AcsmStartAddrXlatVal62.configure(this, null, "");
      this.AcsmStartAddrXlatVal62.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal62, `UVM_REG_ADDR_WIDTH'h362, "RW", 0);
		this.AcsmStartAddrXlatVal62_AcsmStartAddrXlatVal62 = this.AcsmStartAddrXlatVal62.AcsmStartAddrXlatVal62;
      this.AcsmStartAddrXlatVal63 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStartAddrXlatVal63::type_id::create("AcsmStartAddrXlatVal63",,get_full_name());
      if(this.AcsmStartAddrXlatVal63.has_coverage(UVM_CVR_ALL))
      	this.AcsmStartAddrXlatVal63.cg_bits.option.name = {get_name(), ".", "AcsmStartAddrXlatVal63_bits"};
      this.AcsmStartAddrXlatVal63.configure(this, null, "");
      this.AcsmStartAddrXlatVal63.build();
      this.default_map.add_reg(this.AcsmStartAddrXlatVal63, `UVM_REG_ADDR_WIDTH'h363, "RW", 0);
		this.AcsmStartAddrXlatVal63_AcsmStartAddrXlatVal63 = this.AcsmStartAddrXlatVal63.AcsmStartAddrXlatVal63;
      this.AcsmStopAddrXlatVal0 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal0::type_id::create("AcsmStopAddrXlatVal0",,get_full_name());
      if(this.AcsmStopAddrXlatVal0.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal0.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal0_bits"};
      this.AcsmStopAddrXlatVal0.configure(this, null, "");
      this.AcsmStopAddrXlatVal0.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal0, `UVM_REG_ADDR_WIDTH'h38B, "RW", 0);
		this.AcsmStopAddrXlatVal0_AcsmStopAddrXlatVal0 = this.AcsmStopAddrXlatVal0.AcsmStopAddrXlatVal0;
      this.AcsmStopAddrXlatVal1 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal1::type_id::create("AcsmStopAddrXlatVal1",,get_full_name());
      if(this.AcsmStopAddrXlatVal1.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal1.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal1_bits"};
      this.AcsmStopAddrXlatVal1.configure(this, null, "");
      this.AcsmStopAddrXlatVal1.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal1, `UVM_REG_ADDR_WIDTH'h38C, "RW", 0);
		this.AcsmStopAddrXlatVal1_AcsmStopAddrXlatVal1 = this.AcsmStopAddrXlatVal1.AcsmStopAddrXlatVal1;
      this.AcsmStopAddrXlatVal2 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal2::type_id::create("AcsmStopAddrXlatVal2",,get_full_name());
      if(this.AcsmStopAddrXlatVal2.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal2.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal2_bits"};
      this.AcsmStopAddrXlatVal2.configure(this, null, "");
      this.AcsmStopAddrXlatVal2.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal2, `UVM_REG_ADDR_WIDTH'h38D, "RW", 0);
		this.AcsmStopAddrXlatVal2_AcsmStopAddrXlatVal2 = this.AcsmStopAddrXlatVal2.AcsmStopAddrXlatVal2;
      this.AcsmStopAddrXlatVal3 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal3::type_id::create("AcsmStopAddrXlatVal3",,get_full_name());
      if(this.AcsmStopAddrXlatVal3.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal3.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal3_bits"};
      this.AcsmStopAddrXlatVal3.configure(this, null, "");
      this.AcsmStopAddrXlatVal3.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal3, `UVM_REG_ADDR_WIDTH'h38E, "RW", 0);
		this.AcsmStopAddrXlatVal3_AcsmStopAddrXlatVal3 = this.AcsmStopAddrXlatVal3.AcsmStopAddrXlatVal3;
      this.AcsmStopAddrXlatVal4 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal4::type_id::create("AcsmStopAddrXlatVal4",,get_full_name());
      if(this.AcsmStopAddrXlatVal4.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal4.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal4_bits"};
      this.AcsmStopAddrXlatVal4.configure(this, null, "");
      this.AcsmStopAddrXlatVal4.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal4, `UVM_REG_ADDR_WIDTH'h38F, "RW", 0);
		this.AcsmStopAddrXlatVal4_AcsmStopAddrXlatVal4 = this.AcsmStopAddrXlatVal4.AcsmStopAddrXlatVal4;
      this.AcsmStopAddrXlatVal5 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal5::type_id::create("AcsmStopAddrXlatVal5",,get_full_name());
      if(this.AcsmStopAddrXlatVal5.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal5.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal5_bits"};
      this.AcsmStopAddrXlatVal5.configure(this, null, "");
      this.AcsmStopAddrXlatVal5.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal5, `UVM_REG_ADDR_WIDTH'h390, "RW", 0);
		this.AcsmStopAddrXlatVal5_AcsmStopAddrXlatVal5 = this.AcsmStopAddrXlatVal5.AcsmStopAddrXlatVal5;
      this.AcsmStopAddrXlatVal6 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal6::type_id::create("AcsmStopAddrXlatVal6",,get_full_name());
      if(this.AcsmStopAddrXlatVal6.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal6.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal6_bits"};
      this.AcsmStopAddrXlatVal6.configure(this, null, "");
      this.AcsmStopAddrXlatVal6.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal6, `UVM_REG_ADDR_WIDTH'h391, "RW", 0);
		this.AcsmStopAddrXlatVal6_AcsmStopAddrXlatVal6 = this.AcsmStopAddrXlatVal6.AcsmStopAddrXlatVal6;
      this.AcsmStopAddrXlatVal7 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal7::type_id::create("AcsmStopAddrXlatVal7",,get_full_name());
      if(this.AcsmStopAddrXlatVal7.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal7.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal7_bits"};
      this.AcsmStopAddrXlatVal7.configure(this, null, "");
      this.AcsmStopAddrXlatVal7.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal7, `UVM_REG_ADDR_WIDTH'h392, "RW", 0);
		this.AcsmStopAddrXlatVal7_AcsmStopAddrXlatVal7 = this.AcsmStopAddrXlatVal7.AcsmStopAddrXlatVal7;
      this.AcsmStopAddrXlatVal8 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal8::type_id::create("AcsmStopAddrXlatVal8",,get_full_name());
      if(this.AcsmStopAddrXlatVal8.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal8.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal8_bits"};
      this.AcsmStopAddrXlatVal8.configure(this, null, "");
      this.AcsmStopAddrXlatVal8.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal8, `UVM_REG_ADDR_WIDTH'h393, "RW", 0);
		this.AcsmStopAddrXlatVal8_AcsmStopAddrXlatVal8 = this.AcsmStopAddrXlatVal8.AcsmStopAddrXlatVal8;
      this.AcsmStopAddrXlatVal9 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal9::type_id::create("AcsmStopAddrXlatVal9",,get_full_name());
      if(this.AcsmStopAddrXlatVal9.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal9.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal9_bits"};
      this.AcsmStopAddrXlatVal9.configure(this, null, "");
      this.AcsmStopAddrXlatVal9.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal9, `UVM_REG_ADDR_WIDTH'h394, "RW", 0);
		this.AcsmStopAddrXlatVal9_AcsmStopAddrXlatVal9 = this.AcsmStopAddrXlatVal9.AcsmStopAddrXlatVal9;
      this.AcsmStopAddrXlatVal10 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal10::type_id::create("AcsmStopAddrXlatVal10",,get_full_name());
      if(this.AcsmStopAddrXlatVal10.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal10.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal10_bits"};
      this.AcsmStopAddrXlatVal10.configure(this, null, "");
      this.AcsmStopAddrXlatVal10.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal10, `UVM_REG_ADDR_WIDTH'h395, "RW", 0);
		this.AcsmStopAddrXlatVal10_AcsmStopAddrXlatVal10 = this.AcsmStopAddrXlatVal10.AcsmStopAddrXlatVal10;
      this.AcsmStopAddrXlatVal11 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal11::type_id::create("AcsmStopAddrXlatVal11",,get_full_name());
      if(this.AcsmStopAddrXlatVal11.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal11.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal11_bits"};
      this.AcsmStopAddrXlatVal11.configure(this, null, "");
      this.AcsmStopAddrXlatVal11.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal11, `UVM_REG_ADDR_WIDTH'h396, "RW", 0);
		this.AcsmStopAddrXlatVal11_AcsmStopAddrXlatVal11 = this.AcsmStopAddrXlatVal11.AcsmStopAddrXlatVal11;
      this.AcsmStopAddrXlatVal12 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal12::type_id::create("AcsmStopAddrXlatVal12",,get_full_name());
      if(this.AcsmStopAddrXlatVal12.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal12.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal12_bits"};
      this.AcsmStopAddrXlatVal12.configure(this, null, "");
      this.AcsmStopAddrXlatVal12.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal12, `UVM_REG_ADDR_WIDTH'h397, "RW", 0);
		this.AcsmStopAddrXlatVal12_AcsmStopAddrXlatVal12 = this.AcsmStopAddrXlatVal12.AcsmStopAddrXlatVal12;
      this.AcsmStopAddrXlatVal13 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal13::type_id::create("AcsmStopAddrXlatVal13",,get_full_name());
      if(this.AcsmStopAddrXlatVal13.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal13.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal13_bits"};
      this.AcsmStopAddrXlatVal13.configure(this, null, "");
      this.AcsmStopAddrXlatVal13.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal13, `UVM_REG_ADDR_WIDTH'h398, "RW", 0);
		this.AcsmStopAddrXlatVal13_AcsmStopAddrXlatVal13 = this.AcsmStopAddrXlatVal13.AcsmStopAddrXlatVal13;
      this.AcsmStopAddrXlatVal14 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal14::type_id::create("AcsmStopAddrXlatVal14",,get_full_name());
      if(this.AcsmStopAddrXlatVal14.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal14.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal14_bits"};
      this.AcsmStopAddrXlatVal14.configure(this, null, "");
      this.AcsmStopAddrXlatVal14.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal14, `UVM_REG_ADDR_WIDTH'h399, "RW", 0);
		this.AcsmStopAddrXlatVal14_AcsmStopAddrXlatVal14 = this.AcsmStopAddrXlatVal14.AcsmStopAddrXlatVal14;
      this.AcsmStopAddrXlatVal15 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal15::type_id::create("AcsmStopAddrXlatVal15",,get_full_name());
      if(this.AcsmStopAddrXlatVal15.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal15.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal15_bits"};
      this.AcsmStopAddrXlatVal15.configure(this, null, "");
      this.AcsmStopAddrXlatVal15.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal15, `UVM_REG_ADDR_WIDTH'h39A, "RW", 0);
		this.AcsmStopAddrXlatVal15_AcsmStopAddrXlatVal15 = this.AcsmStopAddrXlatVal15.AcsmStopAddrXlatVal15;
      this.AcsmStopAddrXlatVal16 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal16::type_id::create("AcsmStopAddrXlatVal16",,get_full_name());
      if(this.AcsmStopAddrXlatVal16.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal16.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal16_bits"};
      this.AcsmStopAddrXlatVal16.configure(this, null, "");
      this.AcsmStopAddrXlatVal16.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal16, `UVM_REG_ADDR_WIDTH'h39B, "RW", 0);
		this.AcsmStopAddrXlatVal16_AcsmStopAddrXlatVal16 = this.AcsmStopAddrXlatVal16.AcsmStopAddrXlatVal16;
      this.AcsmStopAddrXlatVal17 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal17::type_id::create("AcsmStopAddrXlatVal17",,get_full_name());
      if(this.AcsmStopAddrXlatVal17.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal17.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal17_bits"};
      this.AcsmStopAddrXlatVal17.configure(this, null, "");
      this.AcsmStopAddrXlatVal17.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal17, `UVM_REG_ADDR_WIDTH'h39C, "RW", 0);
		this.AcsmStopAddrXlatVal17_AcsmStopAddrXlatVal17 = this.AcsmStopAddrXlatVal17.AcsmStopAddrXlatVal17;
      this.AcsmStopAddrXlatVal18 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal18::type_id::create("AcsmStopAddrXlatVal18",,get_full_name());
      if(this.AcsmStopAddrXlatVal18.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal18.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal18_bits"};
      this.AcsmStopAddrXlatVal18.configure(this, null, "");
      this.AcsmStopAddrXlatVal18.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal18, `UVM_REG_ADDR_WIDTH'h39D, "RW", 0);
		this.AcsmStopAddrXlatVal18_AcsmStopAddrXlatVal18 = this.AcsmStopAddrXlatVal18.AcsmStopAddrXlatVal18;
      this.AcsmStopAddrXlatVal19 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal19::type_id::create("AcsmStopAddrXlatVal19",,get_full_name());
      if(this.AcsmStopAddrXlatVal19.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal19.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal19_bits"};
      this.AcsmStopAddrXlatVal19.configure(this, null, "");
      this.AcsmStopAddrXlatVal19.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal19, `UVM_REG_ADDR_WIDTH'h39E, "RW", 0);
		this.AcsmStopAddrXlatVal19_AcsmStopAddrXlatVal19 = this.AcsmStopAddrXlatVal19.AcsmStopAddrXlatVal19;
      this.AcsmStopAddrXlatVal20 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal20::type_id::create("AcsmStopAddrXlatVal20",,get_full_name());
      if(this.AcsmStopAddrXlatVal20.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal20.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal20_bits"};
      this.AcsmStopAddrXlatVal20.configure(this, null, "");
      this.AcsmStopAddrXlatVal20.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal20, `UVM_REG_ADDR_WIDTH'h39F, "RW", 0);
		this.AcsmStopAddrXlatVal20_AcsmStopAddrXlatVal20 = this.AcsmStopAddrXlatVal20.AcsmStopAddrXlatVal20;
      this.AcsmStopAddrXlatVal21 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal21::type_id::create("AcsmStopAddrXlatVal21",,get_full_name());
      if(this.AcsmStopAddrXlatVal21.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal21.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal21_bits"};
      this.AcsmStopAddrXlatVal21.configure(this, null, "");
      this.AcsmStopAddrXlatVal21.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal21, `UVM_REG_ADDR_WIDTH'h3A0, "RW", 0);
		this.AcsmStopAddrXlatVal21_AcsmStopAddrXlatVal21 = this.AcsmStopAddrXlatVal21.AcsmStopAddrXlatVal21;
      this.AcsmStopAddrXlatVal22 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal22::type_id::create("AcsmStopAddrXlatVal22",,get_full_name());
      if(this.AcsmStopAddrXlatVal22.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal22.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal22_bits"};
      this.AcsmStopAddrXlatVal22.configure(this, null, "");
      this.AcsmStopAddrXlatVal22.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal22, `UVM_REG_ADDR_WIDTH'h3A1, "RW", 0);
		this.AcsmStopAddrXlatVal22_AcsmStopAddrXlatVal22 = this.AcsmStopAddrXlatVal22.AcsmStopAddrXlatVal22;
      this.AcsmStopAddrXlatVal23 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal23::type_id::create("AcsmStopAddrXlatVal23",,get_full_name());
      if(this.AcsmStopAddrXlatVal23.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal23.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal23_bits"};
      this.AcsmStopAddrXlatVal23.configure(this, null, "");
      this.AcsmStopAddrXlatVal23.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal23, `UVM_REG_ADDR_WIDTH'h3A2, "RW", 0);
		this.AcsmStopAddrXlatVal23_AcsmStopAddrXlatVal23 = this.AcsmStopAddrXlatVal23.AcsmStopAddrXlatVal23;
      this.AcsmStopAddrXlatVal24 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal24::type_id::create("AcsmStopAddrXlatVal24",,get_full_name());
      if(this.AcsmStopAddrXlatVal24.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal24.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal24_bits"};
      this.AcsmStopAddrXlatVal24.configure(this, null, "");
      this.AcsmStopAddrXlatVal24.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal24, `UVM_REG_ADDR_WIDTH'h3A3, "RW", 0);
		this.AcsmStopAddrXlatVal24_AcsmStopAddrXlatVal24 = this.AcsmStopAddrXlatVal24.AcsmStopAddrXlatVal24;
      this.AcsmStopAddrXlatVal25 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal25::type_id::create("AcsmStopAddrXlatVal25",,get_full_name());
      if(this.AcsmStopAddrXlatVal25.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal25.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal25_bits"};
      this.AcsmStopAddrXlatVal25.configure(this, null, "");
      this.AcsmStopAddrXlatVal25.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal25, `UVM_REG_ADDR_WIDTH'h3A4, "RW", 0);
		this.AcsmStopAddrXlatVal25_AcsmStopAddrXlatVal25 = this.AcsmStopAddrXlatVal25.AcsmStopAddrXlatVal25;
      this.AcsmStopAddrXlatVal26 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal26::type_id::create("AcsmStopAddrXlatVal26",,get_full_name());
      if(this.AcsmStopAddrXlatVal26.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal26.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal26_bits"};
      this.AcsmStopAddrXlatVal26.configure(this, null, "");
      this.AcsmStopAddrXlatVal26.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal26, `UVM_REG_ADDR_WIDTH'h3A5, "RW", 0);
		this.AcsmStopAddrXlatVal26_AcsmStopAddrXlatVal26 = this.AcsmStopAddrXlatVal26.AcsmStopAddrXlatVal26;
      this.AcsmStopAddrXlatVal27 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal27::type_id::create("AcsmStopAddrXlatVal27",,get_full_name());
      if(this.AcsmStopAddrXlatVal27.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal27.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal27_bits"};
      this.AcsmStopAddrXlatVal27.configure(this, null, "");
      this.AcsmStopAddrXlatVal27.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal27, `UVM_REG_ADDR_WIDTH'h3A6, "RW", 0);
		this.AcsmStopAddrXlatVal27_AcsmStopAddrXlatVal27 = this.AcsmStopAddrXlatVal27.AcsmStopAddrXlatVal27;
      this.AcsmStopAddrXlatVal28 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal28::type_id::create("AcsmStopAddrXlatVal28",,get_full_name());
      if(this.AcsmStopAddrXlatVal28.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal28.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal28_bits"};
      this.AcsmStopAddrXlatVal28.configure(this, null, "");
      this.AcsmStopAddrXlatVal28.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal28, `UVM_REG_ADDR_WIDTH'h3A7, "RW", 0);
		this.AcsmStopAddrXlatVal28_AcsmStopAddrXlatVal28 = this.AcsmStopAddrXlatVal28.AcsmStopAddrXlatVal28;
      this.AcsmStopAddrXlatVal29 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal29::type_id::create("AcsmStopAddrXlatVal29",,get_full_name());
      if(this.AcsmStopAddrXlatVal29.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal29.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal29_bits"};
      this.AcsmStopAddrXlatVal29.configure(this, null, "");
      this.AcsmStopAddrXlatVal29.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal29, `UVM_REG_ADDR_WIDTH'h3A8, "RW", 0);
		this.AcsmStopAddrXlatVal29_AcsmStopAddrXlatVal29 = this.AcsmStopAddrXlatVal29.AcsmStopAddrXlatVal29;
      this.AcsmStopAddrXlatVal30 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal30::type_id::create("AcsmStopAddrXlatVal30",,get_full_name());
      if(this.AcsmStopAddrXlatVal30.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal30.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal30_bits"};
      this.AcsmStopAddrXlatVal30.configure(this, null, "");
      this.AcsmStopAddrXlatVal30.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal30, `UVM_REG_ADDR_WIDTH'h3A9, "RW", 0);
		this.AcsmStopAddrXlatVal30_AcsmStopAddrXlatVal30 = this.AcsmStopAddrXlatVal30.AcsmStopAddrXlatVal30;
      this.AcsmStopAddrXlatVal31 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal31::type_id::create("AcsmStopAddrXlatVal31",,get_full_name());
      if(this.AcsmStopAddrXlatVal31.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal31.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal31_bits"};
      this.AcsmStopAddrXlatVal31.configure(this, null, "");
      this.AcsmStopAddrXlatVal31.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal31, `UVM_REG_ADDR_WIDTH'h3AA, "RW", 0);
		this.AcsmStopAddrXlatVal31_AcsmStopAddrXlatVal31 = this.AcsmStopAddrXlatVal31.AcsmStopAddrXlatVal31;
      this.AcsmStopAddrXlatVal32 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal32::type_id::create("AcsmStopAddrXlatVal32",,get_full_name());
      if(this.AcsmStopAddrXlatVal32.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal32.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal32_bits"};
      this.AcsmStopAddrXlatVal32.configure(this, null, "");
      this.AcsmStopAddrXlatVal32.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal32, `UVM_REG_ADDR_WIDTH'h3AB, "RW", 0);
		this.AcsmStopAddrXlatVal32_AcsmStopAddrXlatVal32 = this.AcsmStopAddrXlatVal32.AcsmStopAddrXlatVal32;
      this.AcsmStopAddrXlatVal33 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal33::type_id::create("AcsmStopAddrXlatVal33",,get_full_name());
      if(this.AcsmStopAddrXlatVal33.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal33.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal33_bits"};
      this.AcsmStopAddrXlatVal33.configure(this, null, "");
      this.AcsmStopAddrXlatVal33.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal33, `UVM_REG_ADDR_WIDTH'h3AC, "RW", 0);
		this.AcsmStopAddrXlatVal33_AcsmStopAddrXlatVal33 = this.AcsmStopAddrXlatVal33.AcsmStopAddrXlatVal33;
      this.AcsmStopAddrXlatVal34 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal34::type_id::create("AcsmStopAddrXlatVal34",,get_full_name());
      if(this.AcsmStopAddrXlatVal34.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal34.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal34_bits"};
      this.AcsmStopAddrXlatVal34.configure(this, null, "");
      this.AcsmStopAddrXlatVal34.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal34, `UVM_REG_ADDR_WIDTH'h3AD, "RW", 0);
		this.AcsmStopAddrXlatVal34_AcsmStopAddrXlatVal34 = this.AcsmStopAddrXlatVal34.AcsmStopAddrXlatVal34;
      this.AcsmStopAddrXlatVal35 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal35::type_id::create("AcsmStopAddrXlatVal35",,get_full_name());
      if(this.AcsmStopAddrXlatVal35.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal35.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal35_bits"};
      this.AcsmStopAddrXlatVal35.configure(this, null, "");
      this.AcsmStopAddrXlatVal35.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal35, `UVM_REG_ADDR_WIDTH'h3AE, "RW", 0);
		this.AcsmStopAddrXlatVal35_AcsmStopAddrXlatVal35 = this.AcsmStopAddrXlatVal35.AcsmStopAddrXlatVal35;
      this.AcsmStopAddrXlatVal36 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal36::type_id::create("AcsmStopAddrXlatVal36",,get_full_name());
      if(this.AcsmStopAddrXlatVal36.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal36.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal36_bits"};
      this.AcsmStopAddrXlatVal36.configure(this, null, "");
      this.AcsmStopAddrXlatVal36.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal36, `UVM_REG_ADDR_WIDTH'h3AF, "RW", 0);
		this.AcsmStopAddrXlatVal36_AcsmStopAddrXlatVal36 = this.AcsmStopAddrXlatVal36.AcsmStopAddrXlatVal36;
      this.AcsmStopAddrXlatVal37 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal37::type_id::create("AcsmStopAddrXlatVal37",,get_full_name());
      if(this.AcsmStopAddrXlatVal37.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal37.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal37_bits"};
      this.AcsmStopAddrXlatVal37.configure(this, null, "");
      this.AcsmStopAddrXlatVal37.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal37, `UVM_REG_ADDR_WIDTH'h3B0, "RW", 0);
		this.AcsmStopAddrXlatVal37_AcsmStopAddrXlatVal37 = this.AcsmStopAddrXlatVal37.AcsmStopAddrXlatVal37;
      this.AcsmStopAddrXlatVal38 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal38::type_id::create("AcsmStopAddrXlatVal38",,get_full_name());
      if(this.AcsmStopAddrXlatVal38.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal38.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal38_bits"};
      this.AcsmStopAddrXlatVal38.configure(this, null, "");
      this.AcsmStopAddrXlatVal38.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal38, `UVM_REG_ADDR_WIDTH'h3B1, "RW", 0);
		this.AcsmStopAddrXlatVal38_AcsmStopAddrXlatVal38 = this.AcsmStopAddrXlatVal38.AcsmStopAddrXlatVal38;
      this.AcsmStopAddrXlatVal39 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal39::type_id::create("AcsmStopAddrXlatVal39",,get_full_name());
      if(this.AcsmStopAddrXlatVal39.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal39.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal39_bits"};
      this.AcsmStopAddrXlatVal39.configure(this, null, "");
      this.AcsmStopAddrXlatVal39.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal39, `UVM_REG_ADDR_WIDTH'h3B2, "RW", 0);
		this.AcsmStopAddrXlatVal39_AcsmStopAddrXlatVal39 = this.AcsmStopAddrXlatVal39.AcsmStopAddrXlatVal39;
      this.AcsmStopAddrXlatVal40 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal40::type_id::create("AcsmStopAddrXlatVal40",,get_full_name());
      if(this.AcsmStopAddrXlatVal40.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal40.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal40_bits"};
      this.AcsmStopAddrXlatVal40.configure(this, null, "");
      this.AcsmStopAddrXlatVal40.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal40, `UVM_REG_ADDR_WIDTH'h3B3, "RW", 0);
		this.AcsmStopAddrXlatVal40_AcsmStopAddrXlatVal40 = this.AcsmStopAddrXlatVal40.AcsmStopAddrXlatVal40;
      this.AcsmStopAddrXlatVal41 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal41::type_id::create("AcsmStopAddrXlatVal41",,get_full_name());
      if(this.AcsmStopAddrXlatVal41.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal41.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal41_bits"};
      this.AcsmStopAddrXlatVal41.configure(this, null, "");
      this.AcsmStopAddrXlatVal41.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal41, `UVM_REG_ADDR_WIDTH'h3B4, "RW", 0);
		this.AcsmStopAddrXlatVal41_AcsmStopAddrXlatVal41 = this.AcsmStopAddrXlatVal41.AcsmStopAddrXlatVal41;
      this.AcsmStopAddrXlatVal42 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal42::type_id::create("AcsmStopAddrXlatVal42",,get_full_name());
      if(this.AcsmStopAddrXlatVal42.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal42.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal42_bits"};
      this.AcsmStopAddrXlatVal42.configure(this, null, "");
      this.AcsmStopAddrXlatVal42.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal42, `UVM_REG_ADDR_WIDTH'h3B5, "RW", 0);
		this.AcsmStopAddrXlatVal42_AcsmStopAddrXlatVal42 = this.AcsmStopAddrXlatVal42.AcsmStopAddrXlatVal42;
      this.AcsmStopAddrXlatVal43 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal43::type_id::create("AcsmStopAddrXlatVal43",,get_full_name());
      if(this.AcsmStopAddrXlatVal43.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal43.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal43_bits"};
      this.AcsmStopAddrXlatVal43.configure(this, null, "");
      this.AcsmStopAddrXlatVal43.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal43, `UVM_REG_ADDR_WIDTH'h3B6, "RW", 0);
		this.AcsmStopAddrXlatVal43_AcsmStopAddrXlatVal43 = this.AcsmStopAddrXlatVal43.AcsmStopAddrXlatVal43;
      this.AcsmStopAddrXlatVal44 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal44::type_id::create("AcsmStopAddrXlatVal44",,get_full_name());
      if(this.AcsmStopAddrXlatVal44.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal44.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal44_bits"};
      this.AcsmStopAddrXlatVal44.configure(this, null, "");
      this.AcsmStopAddrXlatVal44.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal44, `UVM_REG_ADDR_WIDTH'h3B7, "RW", 0);
		this.AcsmStopAddrXlatVal44_AcsmStopAddrXlatVal44 = this.AcsmStopAddrXlatVal44.AcsmStopAddrXlatVal44;
      this.AcsmStopAddrXlatVal45 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal45::type_id::create("AcsmStopAddrXlatVal45",,get_full_name());
      if(this.AcsmStopAddrXlatVal45.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal45.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal45_bits"};
      this.AcsmStopAddrXlatVal45.configure(this, null, "");
      this.AcsmStopAddrXlatVal45.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal45, `UVM_REG_ADDR_WIDTH'h3B8, "RW", 0);
		this.AcsmStopAddrXlatVal45_AcsmStopAddrXlatVal45 = this.AcsmStopAddrXlatVal45.AcsmStopAddrXlatVal45;
      this.AcsmStopAddrXlatVal46 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal46::type_id::create("AcsmStopAddrXlatVal46",,get_full_name());
      if(this.AcsmStopAddrXlatVal46.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal46.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal46_bits"};
      this.AcsmStopAddrXlatVal46.configure(this, null, "");
      this.AcsmStopAddrXlatVal46.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal46, `UVM_REG_ADDR_WIDTH'h3B9, "RW", 0);
		this.AcsmStopAddrXlatVal46_AcsmStopAddrXlatVal46 = this.AcsmStopAddrXlatVal46.AcsmStopAddrXlatVal46;
      this.AcsmStopAddrXlatVal47 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal47::type_id::create("AcsmStopAddrXlatVal47",,get_full_name());
      if(this.AcsmStopAddrXlatVal47.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal47.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal47_bits"};
      this.AcsmStopAddrXlatVal47.configure(this, null, "");
      this.AcsmStopAddrXlatVal47.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal47, `UVM_REG_ADDR_WIDTH'h3BA, "RW", 0);
		this.AcsmStopAddrXlatVal47_AcsmStopAddrXlatVal47 = this.AcsmStopAddrXlatVal47.AcsmStopAddrXlatVal47;
      this.AcsmStopAddrXlatVal48 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal48::type_id::create("AcsmStopAddrXlatVal48",,get_full_name());
      if(this.AcsmStopAddrXlatVal48.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal48.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal48_bits"};
      this.AcsmStopAddrXlatVal48.configure(this, null, "");
      this.AcsmStopAddrXlatVal48.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal48, `UVM_REG_ADDR_WIDTH'h3BB, "RW", 0);
		this.AcsmStopAddrXlatVal48_AcsmStopAddrXlatVal48 = this.AcsmStopAddrXlatVal48.AcsmStopAddrXlatVal48;
      this.AcsmStopAddrXlatVal49 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal49::type_id::create("AcsmStopAddrXlatVal49",,get_full_name());
      if(this.AcsmStopAddrXlatVal49.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal49.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal49_bits"};
      this.AcsmStopAddrXlatVal49.configure(this, null, "");
      this.AcsmStopAddrXlatVal49.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal49, `UVM_REG_ADDR_WIDTH'h3BC, "RW", 0);
		this.AcsmStopAddrXlatVal49_AcsmStopAddrXlatVal49 = this.AcsmStopAddrXlatVal49.AcsmStopAddrXlatVal49;
      this.AcsmStopAddrXlatVal50 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal50::type_id::create("AcsmStopAddrXlatVal50",,get_full_name());
      if(this.AcsmStopAddrXlatVal50.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal50.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal50_bits"};
      this.AcsmStopAddrXlatVal50.configure(this, null, "");
      this.AcsmStopAddrXlatVal50.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal50, `UVM_REG_ADDR_WIDTH'h3BD, "RW", 0);
		this.AcsmStopAddrXlatVal50_AcsmStopAddrXlatVal50 = this.AcsmStopAddrXlatVal50.AcsmStopAddrXlatVal50;
      this.AcsmStopAddrXlatVal51 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal51::type_id::create("AcsmStopAddrXlatVal51",,get_full_name());
      if(this.AcsmStopAddrXlatVal51.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal51.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal51_bits"};
      this.AcsmStopAddrXlatVal51.configure(this, null, "");
      this.AcsmStopAddrXlatVal51.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal51, `UVM_REG_ADDR_WIDTH'h3BE, "RW", 0);
		this.AcsmStopAddrXlatVal51_AcsmStopAddrXlatVal51 = this.AcsmStopAddrXlatVal51.AcsmStopAddrXlatVal51;
      this.AcsmStopAddrXlatVal52 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal52::type_id::create("AcsmStopAddrXlatVal52",,get_full_name());
      if(this.AcsmStopAddrXlatVal52.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal52.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal52_bits"};
      this.AcsmStopAddrXlatVal52.configure(this, null, "");
      this.AcsmStopAddrXlatVal52.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal52, `UVM_REG_ADDR_WIDTH'h3BF, "RW", 0);
		this.AcsmStopAddrXlatVal52_AcsmStopAddrXlatVal52 = this.AcsmStopAddrXlatVal52.AcsmStopAddrXlatVal52;
      this.AcsmStopAddrXlatVal53 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal53::type_id::create("AcsmStopAddrXlatVal53",,get_full_name());
      if(this.AcsmStopAddrXlatVal53.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal53.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal53_bits"};
      this.AcsmStopAddrXlatVal53.configure(this, null, "");
      this.AcsmStopAddrXlatVal53.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal53, `UVM_REG_ADDR_WIDTH'h3C0, "RW", 0);
		this.AcsmStopAddrXlatVal53_AcsmStopAddrXlatVal53 = this.AcsmStopAddrXlatVal53.AcsmStopAddrXlatVal53;
      this.AcsmStopAddrXlatVal54 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal54::type_id::create("AcsmStopAddrXlatVal54",,get_full_name());
      if(this.AcsmStopAddrXlatVal54.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal54.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal54_bits"};
      this.AcsmStopAddrXlatVal54.configure(this, null, "");
      this.AcsmStopAddrXlatVal54.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal54, `UVM_REG_ADDR_WIDTH'h3C1, "RW", 0);
		this.AcsmStopAddrXlatVal54_AcsmStopAddrXlatVal54 = this.AcsmStopAddrXlatVal54.AcsmStopAddrXlatVal54;
      this.AcsmStopAddrXlatVal55 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal55::type_id::create("AcsmStopAddrXlatVal55",,get_full_name());
      if(this.AcsmStopAddrXlatVal55.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal55.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal55_bits"};
      this.AcsmStopAddrXlatVal55.configure(this, null, "");
      this.AcsmStopAddrXlatVal55.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal55, `UVM_REG_ADDR_WIDTH'h3C2, "RW", 0);
		this.AcsmStopAddrXlatVal55_AcsmStopAddrXlatVal55 = this.AcsmStopAddrXlatVal55.AcsmStopAddrXlatVal55;
      this.AcsmStopAddrXlatVal56 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal56::type_id::create("AcsmStopAddrXlatVal56",,get_full_name());
      if(this.AcsmStopAddrXlatVal56.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal56.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal56_bits"};
      this.AcsmStopAddrXlatVal56.configure(this, null, "");
      this.AcsmStopAddrXlatVal56.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal56, `UVM_REG_ADDR_WIDTH'h3C3, "RW", 0);
		this.AcsmStopAddrXlatVal56_AcsmStopAddrXlatVal56 = this.AcsmStopAddrXlatVal56.AcsmStopAddrXlatVal56;
      this.AcsmStopAddrXlatVal57 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal57::type_id::create("AcsmStopAddrXlatVal57",,get_full_name());
      if(this.AcsmStopAddrXlatVal57.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal57.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal57_bits"};
      this.AcsmStopAddrXlatVal57.configure(this, null, "");
      this.AcsmStopAddrXlatVal57.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal57, `UVM_REG_ADDR_WIDTH'h3C4, "RW", 0);
		this.AcsmStopAddrXlatVal57_AcsmStopAddrXlatVal57 = this.AcsmStopAddrXlatVal57.AcsmStopAddrXlatVal57;
      this.AcsmStopAddrXlatVal58 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal58::type_id::create("AcsmStopAddrXlatVal58",,get_full_name());
      if(this.AcsmStopAddrXlatVal58.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal58.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal58_bits"};
      this.AcsmStopAddrXlatVal58.configure(this, null, "");
      this.AcsmStopAddrXlatVal58.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal58, `UVM_REG_ADDR_WIDTH'h3C5, "RW", 0);
		this.AcsmStopAddrXlatVal58_AcsmStopAddrXlatVal58 = this.AcsmStopAddrXlatVal58.AcsmStopAddrXlatVal58;
      this.AcsmStopAddrXlatVal59 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal59::type_id::create("AcsmStopAddrXlatVal59",,get_full_name());
      if(this.AcsmStopAddrXlatVal59.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal59.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal59_bits"};
      this.AcsmStopAddrXlatVal59.configure(this, null, "");
      this.AcsmStopAddrXlatVal59.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal59, `UVM_REG_ADDR_WIDTH'h3C6, "RW", 0);
		this.AcsmStopAddrXlatVal59_AcsmStopAddrXlatVal59 = this.AcsmStopAddrXlatVal59.AcsmStopAddrXlatVal59;
      this.AcsmStopAddrXlatVal60 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal60::type_id::create("AcsmStopAddrXlatVal60",,get_full_name());
      if(this.AcsmStopAddrXlatVal60.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal60.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal60_bits"};
      this.AcsmStopAddrXlatVal60.configure(this, null, "");
      this.AcsmStopAddrXlatVal60.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal60, `UVM_REG_ADDR_WIDTH'h3C7, "RW", 0);
		this.AcsmStopAddrXlatVal60_AcsmStopAddrXlatVal60 = this.AcsmStopAddrXlatVal60.AcsmStopAddrXlatVal60;
      this.AcsmStopAddrXlatVal61 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal61::type_id::create("AcsmStopAddrXlatVal61",,get_full_name());
      if(this.AcsmStopAddrXlatVal61.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal61.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal61_bits"};
      this.AcsmStopAddrXlatVal61.configure(this, null, "");
      this.AcsmStopAddrXlatVal61.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal61, `UVM_REG_ADDR_WIDTH'h3C8, "RW", 0);
		this.AcsmStopAddrXlatVal61_AcsmStopAddrXlatVal61 = this.AcsmStopAddrXlatVal61.AcsmStopAddrXlatVal61;
      this.AcsmStopAddrXlatVal62 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal62::type_id::create("AcsmStopAddrXlatVal62",,get_full_name());
      if(this.AcsmStopAddrXlatVal62.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal62.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal62_bits"};
      this.AcsmStopAddrXlatVal62.configure(this, null, "");
      this.AcsmStopAddrXlatVal62.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal62, `UVM_REG_ADDR_WIDTH'h3C9, "RW", 0);
		this.AcsmStopAddrXlatVal62_AcsmStopAddrXlatVal62 = this.AcsmStopAddrXlatVal62.AcsmStopAddrXlatVal62;
      this.AcsmStopAddrXlatVal63 = ral_reg_DWC_DDRPHYA_PPGC0_p0_AcsmStopAddrXlatVal63::type_id::create("AcsmStopAddrXlatVal63",,get_full_name());
      if(this.AcsmStopAddrXlatVal63.has_coverage(UVM_CVR_ALL))
      	this.AcsmStopAddrXlatVal63.cg_bits.option.name = {get_name(), ".", "AcsmStopAddrXlatVal63_bits"};
      this.AcsmStopAddrXlatVal63.configure(this, null, "");
      this.AcsmStopAddrXlatVal63.build();
      this.default_map.add_reg(this.AcsmStopAddrXlatVal63, `UVM_REG_ADDR_WIDTH'h3CA, "RW", 0);
		this.AcsmStopAddrXlatVal63_AcsmStopAddrXlatVal63 = this.AcsmStopAddrXlatVal63.AcsmStopAddrXlatVal63;
   endfunction : build

	`uvm_object_utils(ral_block_DWC_DDRPHYA_PPGC0_p0)


function void sample(uvm_reg_addr_t offset,
                     bit            is_read,
                     uvm_reg_map    map);
  if (get_coverage(UVM_CVR_ADDR_MAP)) begin
    m_offset = offset;
    cg_addr.sample();
  end
endfunction
endclass : ral_block_DWC_DDRPHYA_PPGC0_p0


endpackage
`endif
