// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: imc_bank behavioral model.
//
// Authors: Roel Uytterhoeven, Bram Rooseleer
// Owner: Bram Rooseleer <bram.rooseleer@axelera.ai>

`timescale 1ns/1ps

module imc_bank
import imc_bank_pkg::*;
(
  // Common interface
  input	  wire                                  clock,
  input	  wire                                  rst_n,
  input	  wire [IMC_NB_TOTAL_COLS_PER_BANK-2:0] repair_setting,
  input	  wire                                  update_repair_setting,

  // Write interface
  input   wire                                  write_enable,         // weight write enable bit for this block
  input   wire [IMC_ROW_PW-1:0]                 write_row,            // row select address
  input   wire [IMC_WEIGHT_SET_PW-1:0]          write_wss,            // weight set select for weight writing (should never equal compute_wss when w_en is active)
  input   wire [IMC_DATA_W-1:0]                 write_values_0,       // weight values to be written
  input   wire [IMC_DATA_W-1:0]                 write_values_1,
  input   wire [IMC_DATA_W-1:0]                 write_values_2,
  input   wire [IMC_DATA_W-1:0]                 write_values_3,
  input   wire [IMC_DATA_W-1:0]                 write_values_4,
  input   wire [IMC_DATA_W-1:0]                 write_values_5,
  input   wire [IMC_DATA_W-1:0]                 write_values_6,
  input   wire [IMC_DATA_W-1:0]                 write_values_7,
  input   wire [IMC_DATA_W-1:0]                 write_values_8,
  input   wire [IMC_DATA_W-1:0]                 write_values_9,
  input   wire [IMC_DATA_W-1:0]                 write_values_10,
  input   wire [IMC_DATA_W-1:0]                 write_values_11,
  input   wire [IMC_DATA_W-1:0]                 write_values_12,
  input   wire [IMC_DATA_W-1:0]                 write_values_13,
  input   wire [IMC_DATA_W-1:0]                 write_values_14,
  input   wire [IMC_DATA_W-1:0]                 write_values_15,
  input   wire [IMC_DATA_W-1:0]                 write_values_16,
  input   wire [IMC_DATA_W-1:0]                 write_values_17,
  input   wire [IMC_DATA_W-1:0]                 write_values_18,
  input   wire [IMC_DATA_W-1:0]                 write_values_19,
  input   wire [IMC_DATA_W-1:0]                 write_values_20,
  input   wire [IMC_DATA_W-1:0]                 write_values_21,
  input   wire [IMC_DATA_W-1:0]                 write_values_22,
  input   wire [IMC_DATA_W-1:0]                 write_values_23,
  input   wire [IMC_DATA_W-1:0]                 write_values_24,
  input   wire [IMC_DATA_W-1:0]                 write_values_25,
  input   wire [IMC_DATA_W-1:0]                 write_values_26,
  input   wire [IMC_DATA_W-1:0]                 write_values_27,
  input   wire [IMC_DATA_W-1:0]                 write_values_28,
  input   wire [IMC_DATA_W-1:0]                 write_values_29,
  input   wire [IMC_DATA_W-1:0]                 write_values_30,
  input   wire [IMC_DATA_W-1:0]                 write_values_31,
  input   wire [IMC_DATA_W-1:0]                 write_values_32,

  // Compute interface
  input   wire                                  compute_enable,
  input   wire [IMC_NB_ROWS-1:0]                compute_inp,            // compute input vector of 1 bit elements
  input   wire [IMC_WEIGHT_SET_PW-1:0]          compute_wss,            // compute weight set select (should never equal write_wss when w_en is active)
  input   wire [IMC_BLOCK_ENABLE_W-1:0]         compute_block_enable,   // compute block enable. If all blocks enables are disabled (0) then the imc operation equals zero.
  input   wire [1:0]                            compute_weight_format,  // determines how weights should be interpreted (00: unsigned, 01: 4 bit signed, 10: 8 bit signed, 11: 16 bit signed)
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_0,          // Partial accumulation result
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_1,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_2,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_3,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_4,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_5,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_6,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_7,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_8,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_9,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_10,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_11,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_12,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_13,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_14,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_15,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_16,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_17,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_18,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_19,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_20,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_21,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_22,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_23,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_24,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_25,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_26,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_27,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_28,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_29,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_30,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_31,
  output  wire [IMC_OUT_DATA_W-1:0]             compute_out_32
);

    // Quick sanity check on parameters
    // * interface port sizes are hardcoded due to timing annotations
    // * multidimensional interface ports are split (also hardcoded)
    // * logical limitations

    // synopsys translate_off
    initial begin
      assert(IMC_DATA_W == 4);
      assert(1 << IMC_COLUMNS_W > IMC_NB_TOTAL_COLS_PER_BANK)
      assert(IMC_OUT_DATA_W == 15);
      assert(IMC_NB_TOTAL_COLS_PER_BANK == 33);
      assert(IMC_NB_ROWS == 576);
      assert(IMC_ROW_PW == 10);
      assert(IMC_WEIGHT_SET_PW == 2);
      assert(IMC_NB_DELAY_CYCLES > 1);
      assert(IMC_BLOCK_GATING_GRANULARITY == 32);
      assert(IMC_BLOCK_ENABLE_W == 18);
    end
    // synopsys translate_on


    // Bring expanded inputs back to 2d arrays. Expansion is required for lib and lef syntax
    logic [IMC_DATA_W-1:0]      write_values [0:IMC_NB_TOTAL_COLS_PER_BANK-1];
    logic [IMC_OUT_DATA_W-1:0]  compute_out  [0:IMC_NB_TOTAL_COLS_PER_BANK-1];

    assign compute_out_0 = compute_out[0];
    assign compute_out_1 = compute_out[1];
    assign compute_out_2 = compute_out[2];
    assign compute_out_3 = compute_out[3];
    assign compute_out_4 = compute_out[4];
    assign compute_out_5 = compute_out[5];
    assign compute_out_6 = compute_out[6];
    assign compute_out_7 = compute_out[7];
    assign compute_out_8 = compute_out[8];
    assign compute_out_9 = compute_out[9];
    assign compute_out_10 = compute_out[10];
    assign compute_out_11 = compute_out[11];
    assign compute_out_12 = compute_out[12];
    assign compute_out_13 = compute_out[13];
    assign compute_out_14 = compute_out[14];
    assign compute_out_15 = compute_out[15];
    assign compute_out_16 = compute_out[16];
    assign compute_out_17 = compute_out[17];
    assign compute_out_18 = compute_out[18];
    assign compute_out_19 = compute_out[19];
    assign compute_out_20 = compute_out[20];
    assign compute_out_21 = compute_out[21];
    assign compute_out_22 = compute_out[22];
    assign compute_out_23 = compute_out[23];
    assign compute_out_24 = compute_out[24];
    assign compute_out_25 = compute_out[25];
    assign compute_out_26 = compute_out[26];
    assign compute_out_27 = compute_out[27];
    assign compute_out_28 = compute_out[28];
    assign compute_out_29 = compute_out[29];
    assign compute_out_30 = compute_out[30];
    assign compute_out_31 = compute_out[31];
    assign compute_out_32 = compute_out[32];
    assign write_values[0] = write_values_0;
    assign write_values[1] = write_values_1;
    assign write_values[2] = write_values_2;
    assign write_values[3] = write_values_3;
    assign write_values[4] = write_values_4;
    assign write_values[5] = write_values_5;
    assign write_values[6] = write_values_6;
    assign write_values[7] = write_values_7;
    assign write_values[8] = write_values_8;
    assign write_values[9] = write_values_9;
    assign write_values[10] = write_values_10;
    assign write_values[11] = write_values_11;
    assign write_values[12] = write_values_12;
    assign write_values[13] = write_values_13;
    assign write_values[14] = write_values_14;
    assign write_values[15] = write_values_15;
    assign write_values[16] = write_values_16;
    assign write_values[17] = write_values_17;
    assign write_values[18] = write_values_18;
    assign write_values[19] = write_values_19;
    assign write_values[20] = write_values_20;
    assign write_values[21] = write_values_21;
    assign write_values[22] = write_values_22;
    assign write_values[23] = write_values_23;
    assign write_values[24] = write_values_24;
    assign write_values[25] = write_values_25;
    assign write_values[26] = write_values_26;
    assign write_values[27] = write_values_27;
    assign write_values[28] = write_values_28;
    assign write_values[29] = write_values_29;
    assign write_values[30] = write_values_30;
    assign write_values[31] = write_values_31;
    assign write_values[32] = write_values_32;


      ////////////////////////
     // Internal registers //
    ////////////////////////

    // Instantiation of the compute input registers
    logic [IMC_NB_ROWS-1:0] compute_inp_q;
    logic [IMC_WEIGHT_SET_PW-1:0] compute_wss_q;
    logic [IMC_BLOCK_ENABLE_W-1:0] compute_block_enable_q;
    logic [1:0] compute_weight_format_q;
    logic compute_enable_q;

    // Instantiation of the write input registers
    logic [IMC_WEIGHT_SET_PW-1:0] write_wss_q;
    logic write_enable_q;

    // Instantiation of the weight storage elements
    // for Veloce:
    // pragma attribute WEIGHTS logic_block 1
    logic [IMC_DATA_W-1:0] WEIGHTS [0:IMC_NB_WEIGHT_SETS-1][0:IMC_NB_ROWS-1][0:IMC_NB_TOTAL_COLS_PER_BANK-1];

    // Instantiation of the repair settings registers
    logic [IMC_NB_TOTAL_COLS_PER_BANK-2:0] REPAIR;

    // Instantiation of the output pipeline
    logic signed [IMC_OUT_DATA_W-1:0] OUT [0:IMC_NB_TOTAL_COLS_PER_BANK-1][0:IMC_NB_DELAY_CYCLES-2];


      ///////////
     // Reset //
    ///////////

    bit reset_used_reg;
    wire reset_used = reset_used_reg === 1'b1;
    always @(negedge rst_n) begin
        reset_used_reg <= 1'b1;
    end


      ////////////////////////////
     // Update repair settings //
    ////////////////////////////

    always_ff @(posedge clock or negedge rst_n) begin
      // When update_repair_setting, store the repair_setting input vector
      // weights and pipeline should also be invalidated
      if(!rst_n) begin
        REPAIR <= 0;
      end else if(update_repair_setting) begin
        REPAIR <= repair_setting;
        assert($onehot0(-repair_setting));
      end
    end
    //one-hot bus indicating which column is skipped
    wire [IMC_NB_TOTAL_COLS_PER_BANK-1:0] unused_column;
    assign unused_column = -{1'b1, REPAIR};


      //////////////////////
     // Write conflicts  //
    //////////////////////

    logic concurrent_compute_write_conflict;
    always @(posedge clock)
      concurrent_compute_write_conflict <= write_enable & compute_enable & (compute_wss == write_wss);

    logic pipeline_stall_write_conflict;
    always @(posedge clock) begin
      write_wss_q <= write_wss;
      write_enable_q <= write_enable;
      compute_enable_q <= compute_enable;
      if(write_enable & !compute_enable & (compute_wss_q == write_wss))
        pipeline_stall_write_conflict <= 1;
      else if(compute_enable)
        pipeline_stall_write_conflict <= 0;
    end

    wss_collision: assert property(
      @(posedge clock) disable iff($isunknown(write_wss) || $isunknown(compute_wss))
        write_enable && compute_enable |-> (write_wss != compute_wss)
    ) else $warning("write_wss %b equals compute_wss %b when write_enable and compute_enable active. Output corrupted at time %d", write_wss, compute_wss, $time);


      /////////////////////
     // Write operation //
    /////////////////////

    always_ff @(posedge clock or negedge rst_n) begin
      // When write_enable, write the entire weight vector to the correct row of weights
      if(!rst_n || update_repair_setting) begin
        foreach(WEIGHTS[w,r,c]) begin
          `ifndef IMC_DISABLE_RESET_WEIGHTS
            WEIGHTS[w][r][c] <= 4'bxxxx;
          `endif
        end
      end else if(write_enable) begin
        foreach(write_values[i]) begin
          WEIGHTS[write_wss][write_row][i] <= write_values[i];
        end
      end
    end

      ///////////////////////
     // Compute operation //
    ///////////////////////

    // Ensure no compute operation is started before reset
    compute_before_reset: assert property(
      @(posedge clock)
        compute_enable |-> reset_used
    ) else $warning("compute operation stared before reset at time %d", $time);

    // Last pipeline stage is presented towards the outside.
    always_comb
      foreach(compute_out[c]) compute_out[c] = OUT[c][IMC_NB_DELAY_CYCLES-2];

    // Compute logic
    function [IMC_COLUMNS_W-1:0] relative_column;
      input [IMC_COLUMNS_W-1:0] column;
      relative_column = column - {1'b1, REPAIR}[column];
    endfunction

    function automatic sign;
      input [IMC_COLUMNS_W-1:0] column;
      case(compute_weight_format_q)
        2'b00: sign = 1'b0;
        2'b01: sign = 1'b1;
        2'b10: sign = relative_column(column)%2 == 1;
        2'b11: sign = relative_column(column)%4 == 3;
      endcase
    endfunction

    function automatic signed [14:0] column_sum;
      input [IMC_COLUMNS_W-1:0] column;
      if(unused_column[column]) begin
        // 'broken' column
        column_sum = 15'hxxxx;
      end else if(!reset_used) begin
        // compute started before reset, correct results cannot be guaranteed (also covered by assert)
        column_sum = 15'hxxxx;
      end else if(!$onehot0(-repair_setting)) begin
        // invalid repair settings (also covered by assert)
        column_sum = 15'hxxxx;
      end else if(concurrent_compute_write_conflict) begin
        // simultaneous compute and write on same weight set (also covered by assert)
        column_sum = 15'hxxxx;
      end
      `ifndef IMC_STALL_CONFLICT_MIMIC_IMPLEMENTATION
      else if(pipeline_stall_write_conflict) begin
        // write happened on stalled compute results
        column_sum = 15'hxxxx;
      end
      `endif
      else begin
        column_sum = 0;
        for(int r=0; r<IMC_NB_ROWS; r++) begin
          column_sum = column_sum + (
            (sign(column) ? (WEIGHTS[compute_wss_q][r][column] + 8)%16 - 8 : WEIGHTS[compute_wss_q][r][column]) &
            ({15{compute_block_enable_q[r/IMC_BLOCK_GATING_GRANULARITY] & compute_inp_q[r]}}));
        end
      end
    endfunction

    // When compute_enable, advance the pipeline and enter new compute results
    always_ff @(posedge clock or negedge rst_n) begin
      if(!rst_n || update_repair_setting) begin
        foreach(OUT[c,p])
          OUT[c][p] <= 15'hxxxx;
        compute_inp_q <= {576{1'bx}};
        compute_wss_q <= 2'bxx;
        compute_block_enable_q <= {18{1'bx}};
        compute_weight_format_q <= 2'bxx;
      end else if(compute_enable) begin
        compute_inp_q <= compute_inp;
        compute_wss_q <= compute_wss;
        compute_block_enable_q <= compute_block_enable;
        compute_weight_format_q <= compute_weight_format;
        // operation per column
        for(int c = 0; c < IMC_NB_TOTAL_COLS_PER_BANK; c++) begin
          OUT[c][0] <= column_sum(c);
          for(int p = 1; p < IMC_NB_DELAY_CYCLES-1; p++)
            OUT[c][p] <= OUT[c][p-1];
        end
      end
    end


      ////////////////////////
     // Timing annotations //
    ////////////////////////

    `ifdef IMC_SPECIFY
    reg notif;
    specify
      specparam
        trise=0,
        tfall=0,
        tpck=0.495,
        tnck=0.495,
        tckp=1.240,
        tdef=0.150;
      (posedge clock *> compute_out_0) = (trise,tfall);
      (posedge clock *> compute_out_1) = (trise,tfall);
      (posedge clock *> compute_out_2) = (trise,tfall);
      (posedge clock *> compute_out_3) = (trise,tfall);
      (posedge clock *> compute_out_4) = (trise,tfall);
      (posedge clock *> compute_out_5) = (trise,tfall);
      (posedge clock *> compute_out_6) = (trise,tfall);
      (posedge clock *> compute_out_7) = (trise,tfall);
      (posedge clock *> compute_out_8) = (trise,tfall);
      (posedge clock *> compute_out_9) = (trise,tfall);
      (posedge clock *> compute_out_10) = (trise,tfall);
      (posedge clock *> compute_out_11) = (trise,tfall);
      (posedge clock *> compute_out_12) = (trise,tfall);
      (posedge clock *> compute_out_13) = (trise,tfall);
      (posedge clock *> compute_out_14) = (trise,tfall);
      (posedge clock *> compute_out_15) = (trise,tfall);
      (posedge clock *> compute_out_16) = (trise,tfall);
      (posedge clock *> compute_out_17) = (trise,tfall);
      (posedge clock *> compute_out_18) = (trise,tfall);
      (posedge clock *> compute_out_19) = (trise,tfall);
      (posedge clock *> compute_out_20) = (trise,tfall);
      (posedge clock *> compute_out_21) = (trise,tfall);
      (posedge clock *> compute_out_22) = (trise,tfall);
      (posedge clock *> compute_out_23) = (trise,tfall);
      (posedge clock *> compute_out_24) = (trise,tfall);
      (posedge clock *> compute_out_25) = (trise,tfall);
      (posedge clock *> compute_out_26) = (trise,tfall);
      (posedge clock *> compute_out_27) = (trise,tfall);
      (posedge clock *> compute_out_28) = (trise,tfall);
      (posedge clock *> compute_out_29) = (trise,tfall);
      (posedge clock *> compute_out_30) = (trise,tfall);
      (posedge clock *> compute_out_31) = (trise,tfall);
      (posedge clock *> compute_out_32) = (trise,tfall);
      $width(posedge clock, tpck, 0, notif);
      $width(negedge clock, tnck, 0, notif);
      $period(posedge clock, tckp, notif);
      $period(negedge clock, tckp, notif);

      $setuphold(posedge clock, posedge update_repair_setting, tdef, tdef, notif);
      $setuphold(posedge clock, negedge update_repair_setting, tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[4], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[4], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[5], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[5], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[6], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[6], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[7], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[7], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[8], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[8], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[9], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[9], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[10], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[10], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[11], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[11], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[12], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[12], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[13], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[13], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[14], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[14], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[15], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[15], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[16], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[16], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[17], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[17], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[18], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[18], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[19], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[19], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[20], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[20], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[21], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[21], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[22], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[22], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[23], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[23], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[24], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[24], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[25], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[25], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[26], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[26], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[27], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[27], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[28], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[28], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[29], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[29], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[30], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[30], tdef, tdef, notif);
      $setuphold(posedge clock, posedge repair_setting[31], tdef, tdef, notif);
      $setuphold(posedge clock, negedge repair_setting[31], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[4], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[4], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[5], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[5], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[6], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[6], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[7], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[7], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[8], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[8], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[9], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[9], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[10], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[10], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[11], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[11], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[12], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[12], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[13], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[13], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[14], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[14], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[15], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[15], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[16], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[16], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_block_enable[17], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_block_enable[17], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_enable, tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_enable, tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[4], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[4], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[5], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[5], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[6], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[6], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[7], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[7], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[8], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[8], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[9], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[9], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[10], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[10], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[11], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[11], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[12], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[12], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[13], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[13], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[14], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[14], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[15], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[15], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[16], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[16], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[17], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[17], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[18], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[18], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[19], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[19], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[20], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[20], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[21], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[21], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[22], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[22], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[23], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[23], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[24], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[24], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[25], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[25], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[26], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[26], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[27], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[27], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[28], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[28], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[29], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[29], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[30], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[30], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[31], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[31], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[32], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[32], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[33], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[33], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[34], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[34], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[35], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[35], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[36], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[36], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[37], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[37], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[38], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[38], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[39], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[39], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[40], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[40], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[41], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[41], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[42], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[42], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[43], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[43], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[44], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[44], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[45], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[45], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[46], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[46], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[47], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[47], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[48], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[48], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[49], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[49], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[50], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[50], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[51], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[51], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[52], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[52], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[53], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[53], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[54], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[54], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[55], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[55], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[56], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[56], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[57], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[57], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[58], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[58], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[59], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[59], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[60], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[60], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[61], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[61], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[62], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[62], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[63], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[63], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[64], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[64], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[65], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[65], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[66], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[66], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[67], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[67], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[68], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[68], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[69], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[69], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[70], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[70], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[71], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[71], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[72], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[72], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[73], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[73], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[74], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[74], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[75], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[75], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[76], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[76], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[77], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[77], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[78], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[78], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[79], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[79], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[80], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[80], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[81], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[81], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[82], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[82], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[83], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[83], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[84], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[84], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[85], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[85], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[86], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[86], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[87], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[87], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[88], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[88], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[89], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[89], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[90], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[90], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[91], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[91], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[92], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[92], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[93], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[93], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[94], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[94], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[95], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[95], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[96], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[96], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[97], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[97], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[98], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[98], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[99], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[99], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[100], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[100], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[101], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[101], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[102], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[102], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[103], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[103], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[104], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[104], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[105], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[105], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[106], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[106], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[107], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[107], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[108], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[108], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[109], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[109], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[110], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[110], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[111], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[111], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[112], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[112], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[113], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[113], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[114], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[114], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[115], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[115], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[116], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[116], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[117], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[117], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[118], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[118], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[119], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[119], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[120], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[120], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[121], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[121], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[122], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[122], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[123], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[123], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[124], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[124], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[125], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[125], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[126], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[126], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[127], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[127], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[128], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[128], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[129], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[129], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[130], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[130], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[131], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[131], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[132], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[132], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[133], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[133], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[134], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[134], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[135], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[135], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[136], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[136], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[137], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[137], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[138], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[138], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[139], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[139], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[140], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[140], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[141], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[141], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[142], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[142], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[143], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[143], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[144], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[144], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[145], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[145], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[146], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[146], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[147], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[147], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[148], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[148], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[149], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[149], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[150], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[150], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[151], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[151], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[152], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[152], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[153], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[153], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[154], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[154], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[155], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[155], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[156], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[156], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[157], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[157], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[158], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[158], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[159], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[159], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[160], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[160], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[161], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[161], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[162], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[162], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[163], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[163], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[164], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[164], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[165], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[165], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[166], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[166], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[167], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[167], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[168], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[168], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[169], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[169], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[170], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[170], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[171], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[171], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[172], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[172], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[173], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[173], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[174], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[174], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[175], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[175], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[176], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[176], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[177], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[177], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[178], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[178], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[179], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[179], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[180], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[180], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[181], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[181], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[182], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[182], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[183], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[183], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[184], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[184], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[185], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[185], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[186], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[186], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[187], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[187], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[188], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[188], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[189], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[189], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[190], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[190], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[191], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[191], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[192], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[192], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[193], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[193], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[194], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[194], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[195], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[195], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[196], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[196], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[197], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[197], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[198], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[198], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[199], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[199], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[200], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[200], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[201], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[201], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[202], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[202], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[203], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[203], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[204], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[204], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[205], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[205], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[206], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[206], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[207], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[207], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[208], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[208], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[209], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[209], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[210], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[210], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[211], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[211], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[212], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[212], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[213], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[213], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[214], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[214], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[215], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[215], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[216], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[216], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[217], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[217], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[218], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[218], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[219], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[219], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[220], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[220], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[221], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[221], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[222], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[222], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[223], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[223], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[224], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[224], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[225], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[225], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[226], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[226], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[227], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[227], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[228], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[228], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[229], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[229], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[230], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[230], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[231], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[231], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[232], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[232], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[233], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[233], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[234], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[234], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[235], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[235], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[236], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[236], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[237], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[237], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[238], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[238], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[239], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[239], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[240], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[240], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[241], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[241], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[242], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[242], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[243], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[243], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[244], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[244], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[245], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[245], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[246], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[246], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[247], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[247], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[248], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[248], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[249], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[249], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[250], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[250], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[251], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[251], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[252], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[252], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[253], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[253], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[254], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[254], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[255], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[255], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[256], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[256], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[257], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[257], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[258], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[258], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[259], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[259], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[260], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[260], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[261], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[261], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[262], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[262], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[263], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[263], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[264], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[264], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[265], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[265], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[266], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[266], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[267], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[267], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[268], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[268], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[269], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[269], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[270], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[270], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[271], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[271], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[272], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[272], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[273], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[273], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[274], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[274], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[275], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[275], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[276], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[276], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[277], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[277], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[278], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[278], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[279], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[279], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[280], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[280], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[281], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[281], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[282], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[282], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[283], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[283], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[284], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[284], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[285], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[285], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[286], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[286], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[287], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[287], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[288], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[288], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[289], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[289], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[290], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[290], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[291], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[291], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[292], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[292], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[293], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[293], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[294], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[294], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[295], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[295], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[296], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[296], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[297], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[297], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[298], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[298], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[299], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[299], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[300], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[300], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[301], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[301], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[302], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[302], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[303], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[303], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[304], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[304], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[305], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[305], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[306], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[306], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[307], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[307], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[308], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[308], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[309], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[309], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[310], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[310], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[311], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[311], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[312], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[312], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[313], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[313], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[314], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[314], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[315], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[315], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[316], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[316], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[317], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[317], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[318], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[318], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[319], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[319], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[320], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[320], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[321], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[321], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[322], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[322], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[323], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[323], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[324], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[324], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[325], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[325], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[326], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[326], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[327], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[327], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[328], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[328], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[329], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[329], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[330], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[330], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[331], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[331], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[332], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[332], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[333], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[333], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[334], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[334], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[335], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[335], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[336], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[336], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[337], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[337], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[338], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[338], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[339], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[339], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[340], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[340], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[341], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[341], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[342], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[342], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[343], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[343], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[344], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[344], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[345], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[345], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[346], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[346], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[347], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[347], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[348], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[348], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[349], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[349], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[350], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[350], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[351], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[351], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[352], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[352], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[353], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[353], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[354], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[354], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[355], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[355], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[356], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[356], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[357], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[357], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[358], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[358], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[359], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[359], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[360], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[360], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[361], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[361], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[362], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[362], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[363], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[363], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[364], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[364], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[365], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[365], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[366], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[366], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[367], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[367], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[368], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[368], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[369], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[369], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[370], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[370], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[371], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[371], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[372], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[372], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[373], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[373], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[374], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[374], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[375], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[375], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[376], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[376], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[377], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[377], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[378], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[378], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[379], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[379], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[380], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[380], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[381], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[381], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[382], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[382], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[383], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[383], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[384], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[384], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[385], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[385], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[386], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[386], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[387], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[387], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[388], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[388], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[389], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[389], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[390], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[390], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[391], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[391], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[392], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[392], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[393], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[393], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[394], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[394], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[395], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[395], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[396], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[396], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[397], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[397], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[398], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[398], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[399], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[399], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[400], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[400], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[401], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[401], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[402], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[402], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[403], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[403], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[404], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[404], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[405], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[405], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[406], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[406], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[407], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[407], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[408], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[408], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[409], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[409], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[410], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[410], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[411], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[411], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[412], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[412], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[413], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[413], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[414], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[414], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[415], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[415], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[416], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[416], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[417], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[417], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[418], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[418], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[419], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[419], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[420], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[420], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[421], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[421], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[422], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[422], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[423], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[423], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[424], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[424], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[425], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[425], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[426], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[426], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[427], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[427], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[428], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[428], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[429], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[429], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[430], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[430], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[431], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[431], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[432], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[432], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[433], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[433], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[434], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[434], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[435], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[435], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[436], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[436], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[437], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[437], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[438], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[438], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[439], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[439], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[440], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[440], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[441], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[441], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[442], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[442], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[443], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[443], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[444], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[444], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[445], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[445], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[446], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[446], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[447], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[447], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[448], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[448], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[449], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[449], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[450], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[450], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[451], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[451], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[452], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[452], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[453], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[453], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[454], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[454], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[455], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[455], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[456], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[456], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[457], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[457], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[458], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[458], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[459], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[459], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[460], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[460], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[461], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[461], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[462], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[462], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[463], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[463], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[464], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[464], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[465], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[465], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[466], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[466], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[467], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[467], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[468], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[468], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[469], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[469], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[470], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[470], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[471], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[471], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[472], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[472], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[473], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[473], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[474], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[474], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[475], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[475], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[476], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[476], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[477], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[477], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[478], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[478], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[479], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[479], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[480], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[480], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[481], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[481], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[482], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[482], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[483], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[483], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[484], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[484], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[485], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[485], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[486], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[486], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[487], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[487], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[488], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[488], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[489], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[489], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[490], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[490], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[491], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[491], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[492], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[492], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[493], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[493], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[494], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[494], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[495], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[495], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[496], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[496], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[497], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[497], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[498], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[498], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[499], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[499], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[500], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[500], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[501], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[501], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[502], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[502], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[503], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[503], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[504], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[504], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[505], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[505], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[506], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[506], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[507], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[507], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[508], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[508], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[509], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[509], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[510], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[510], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[511], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[511], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[512], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[512], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[513], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[513], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[514], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[514], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[515], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[515], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[516], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[516], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[517], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[517], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[518], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[518], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[519], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[519], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[520], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[520], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[521], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[521], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[522], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[522], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[523], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[523], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[524], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[524], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[525], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[525], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[526], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[526], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[527], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[527], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[528], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[528], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[529], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[529], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[530], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[530], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[531], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[531], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[532], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[532], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[533], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[533], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[534], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[534], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[535], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[535], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[536], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[536], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[537], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[537], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[538], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[538], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[539], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[539], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[540], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[540], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[541], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[541], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[542], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[542], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[543], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[543], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[544], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[544], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[545], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[545], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[546], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[546], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[547], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[547], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[548], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[548], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[549], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[549], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[550], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[550], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[551], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[551], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[552], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[552], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[553], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[553], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[554], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[554], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[555], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[555], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[556], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[556], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[557], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[557], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[558], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[558], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[559], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[559], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[560], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[560], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[561], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[561], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[562], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[562], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[563], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[563], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[564], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[564], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[565], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[565], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[566], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[566], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[567], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[567], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[568], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[568], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[569], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[569], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[570], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[570], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[571], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[571], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[572], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[572], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[573], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[573], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[574], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[574], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_inp[575], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_inp[575], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_weight_format[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_weight_format[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_weight_format[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_weight_format[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_wss[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_wss[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge compute_wss[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge compute_wss[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_enable, tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_enable, tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[4], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[4], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[5], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[5], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[6], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[6], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[7], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[7], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[8], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[8], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_row[9], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_row[9], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_0[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_0[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_0[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_0[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_0[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_0[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_0[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_0[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_1[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_1[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_1[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_1[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_1[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_1[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_1[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_1[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_2[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_2[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_2[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_2[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_2[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_2[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_2[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_2[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_3[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_3[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_3[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_3[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_3[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_3[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_3[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_3[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_4[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_4[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_4[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_4[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_4[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_4[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_4[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_4[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_5[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_5[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_5[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_5[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_5[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_5[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_5[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_5[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_6[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_6[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_6[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_6[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_6[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_6[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_6[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_6[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_7[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_7[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_7[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_7[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_7[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_7[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_7[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_7[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_8[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_8[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_8[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_8[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_8[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_8[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_8[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_8[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_9[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_9[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_9[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_9[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_9[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_9[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_9[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_9[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_10[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_10[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_10[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_10[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_10[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_10[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_10[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_10[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_11[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_11[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_11[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_11[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_11[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_11[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_11[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_11[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_12[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_12[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_12[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_12[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_12[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_12[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_12[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_12[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_13[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_13[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_13[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_13[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_13[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_13[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_13[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_13[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_14[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_14[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_14[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_14[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_14[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_14[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_14[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_14[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_15[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_15[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_15[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_15[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_15[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_15[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_15[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_15[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_16[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_16[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_16[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_16[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_16[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_16[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_16[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_16[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_17[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_17[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_17[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_17[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_17[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_17[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_17[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_17[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_18[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_18[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_18[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_18[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_18[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_18[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_18[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_18[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_19[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_19[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_19[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_19[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_19[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_19[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_19[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_19[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_20[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_20[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_20[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_20[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_20[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_20[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_20[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_20[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_21[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_21[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_21[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_21[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_21[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_21[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_21[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_21[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_22[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_22[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_22[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_22[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_22[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_22[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_22[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_22[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_23[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_23[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_23[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_23[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_23[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_23[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_23[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_23[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_24[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_24[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_24[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_24[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_24[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_24[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_24[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_24[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_25[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_25[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_25[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_25[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_25[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_25[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_25[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_25[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_26[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_26[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_26[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_26[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_26[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_26[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_26[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_26[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_27[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_27[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_27[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_27[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_27[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_27[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_27[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_27[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_28[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_28[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_28[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_28[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_28[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_28[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_28[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_28[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_29[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_29[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_29[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_29[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_29[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_29[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_29[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_29[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_30[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_30[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_30[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_30[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_30[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_30[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_30[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_30[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_31[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_31[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_31[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_31[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_31[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_31[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_31[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_31[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_32[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_32[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_32[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_32[1], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_32[2], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_32[2], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_values_32[3], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_values_32[3], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_wss[0], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_wss[0], tdef, tdef, notif);
      $setuphold(posedge clock, posedge write_wss[1], tdef, tdef, notif);
      $setuphold(posedge clock, negedge write_wss[1], tdef, tdef, notif);
    endspecify

    `endif

endmodule
