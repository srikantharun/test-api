// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: Manuel Oliveira <manuel.oliveira@axelera.ai>

/// Bind SVA in imc_bank
///

bind imc_bank imc_bank_sva u_imc_bank_sva (.*);
