// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: {{ cookiecutter.author_full_name }} <{{ cookiecutter.author_email }}>

/// TODO:__one_line_summary_of_{{ cookiecutter.block_name }}__
///
module {{ cookiecutter.block_name }} (
  /// Clock, positive edge triggered
  input  wire i_clk,
  /// Asynchronous reset, active low
  input  wire i_rst_n,


);


endmodule
