// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024



`ifndef GUARD__TREK_TLM_ADAPTER__SV
`define GUARD__TREK_TLM_ADAPTER__SV


`ifndef TREK_TLM_ADAPTER_VIP_BASE_TYPE
`define TREK_TLM_ADAPTER_VIP_BASE_TYPE uvm_pkg::uvm_sequence_item
`endif

// Users specialize this class to provide a conversion between the TLM
// transaction datatypes used by Trek5 and the datatypes used by their
// VIPs.
//
// Note that this class is virtual. You MUST extend it to use it.
//
// This class does not have any dependencies on UVM, although the
// datatypes used to parameterize it may (or may not).
//
virtual class trek_tlm_adapter#(
    type VIP_REQ  = `TREK_TLM_ADAPTER_VIP_BASE_TYPE,
    type VIP_RSP  = VIP_REQ,
    type TREK_REQ = int,
    type TREK_RSP = TREK_REQ);

  TREK_REQ  m_req;  // Composing a response may require the request.
  string    m_name;

  function new(string name = "trek_tlm_adapter");
    m_name = name;
  endfunction

  function string get_name();
    return m_name;
  endfunction

  // Convert the datatype sent by Trek to the datatype used by the VIP.
  //
  pure virtual function VIP_REQ  trek2req(TREK_REQ t);

  // Convert the VIP response datatype to the type expected by Trek.
  //
  pure virtual function TREK_RSP rsp2trek(VIP_RSP t);

endclass: trek_tlm_adapter

`endif // GUARD__TREK_TLM_ADAPTER__SV
