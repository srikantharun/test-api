// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024


`define DELAY_CLK   hdl_top.clk
`define DELAY_INIT  hdl_top.rst_n

`ifndef GUARD__TREK_UVM__SV
`define GUARD__TREK_UVM__SV

`define TREK_C2T_MBOX_SIZE (2 * 8)  // two words of 8-bytes each

// This module contains the method that the user calls to start TrekSoC.
// It also contains methods that are called by TrekSoc, to indicate that
// transaction data is available, and to issue messages in a consistent manner.
module trek_uvm();
`ifdef VERILATOR
`include "trek_dpi.sv"
  typedef enum {UVM_NONE   = 0,   // This typedef is copied from 
                UVM_LOW    = 100, //   "uvm_object_globals.svh"
                UVM_MEDIUM = 200, // Please see the copyright
                UVM_HIGH   = 300, //   in that file...
                UVM_FULL   = 400,
                UVM_DEBUG  = 500} uvm_verbosity;
`else // ~VERILATOR
  import uvm_pkg::*;

  import trek_dpi_pkg::*;
  import trek_uvm_pkg::*;
`endif // VERILATOR

  // mailbox addresses
  bit                       trek_started  = 1'b0;
  bit                       trek_finished = 1'b0;
  longint unsigned          c2t_mboxes_base;
  int unsigned              sdv_threads;
  longint unsigned          seed;
`ifndef VERILATOR
  trek_mbox_wrapper         mbox_wrapper;
`endif

  import "DPI-C" context function int trek_uvm_start_tbx(
      input string            tbx_file,
      output longint unsigned c2t_mboxes_base,
      output int unsigned     sdv_threads,
      output longint unsigned seed,
      input int unsigned      run_mode);

  import "DPI-C" context function int trek_solver_begin(
    input longint unsigned seed = 64'h0,
    input int is_reactive = 1);
  import "DPI-C" context function int trek_solver_end();

  import "DPI-C" context function int trek_entry(
    input string entryAction);
  import "DPI-C" context function int trek_reactive_entry(
    input string entryAction);

 //  export "DPI-C" function trek_tlm_avail_callback;
 //  export "DPI-C" function trek_end_of_test_callback;
 //  export "DPI-C" function trek_get_time;

 //  export "DPI-C" function trek_info_callback;
 //  export "DPI-C" function trek_warn_callback;
 //  export "DPI-C" function trek_error_callback;
 //  export "DPI-C" function trek_fatal_callback;

 //  export "DPI-C" function trek_backdoor_read64;
 //  export "DPI-C" function trek_backdoor_write64;
`ifndef VERILATOR
  mailbox#(longint unsigned)  trek_mbox_event;
`endif

  // *** IMPORTANT ***
  // You must define the methods "trek_backdoor_read64()" and
  // "trek_backdoor_write64()" void functions for your system
  // and put them in a file with this name so the compiler
  // fetches it here! They need to appear in this "scope".
`include "trek_user_backdoor.sv"

`ifndef VERILATOR
  initial begin: mbox_watcher
    mbox_wrapper = new("mbox_wrapper");
    uvm_config_db#(trek_mbox_wrapper)::set(
       uvm_root::get(), "*", "mbox_wrapper", mbox_wrapper);
    fork
      forever begin: loop
        longint unsigned  addr;
        mbox_wrapper.mbox_event.get(addr);
        if (trek_is_c2t_event_addr(addr)) begin: hit
          trek_poll_mbox();
        end
      end
    join_none
  end
`endif // ~VERILATOR

  function automatic void trek_poll_mbox();
    if (trek_started == 1'b0)  // cannot poll before Trek has started
      return;
    for (int unsigned thread_id=0; thread_id<sdv_threads; thread_id++) begin
      longint unsigned data_addr, data, valid_addr, valid;
      data_addr = c2t_mboxes_base + (thread_id * `TREK_C2T_MBOX_SIZE);

      valid_addr = data_addr + 8;
      trek_backdoor_read64(valid_addr, valid, 0 /* debug */);
      if (valid != 64'h0) begin: maibox_has_data
        trek_backdoor_read64(data_addr, data, 0 /* debug */);
        trek_info_callback(
          $sformatf("trek_poll_mbox(): trek_c2t_message [thread=%02d]: read='h%0h",
                    thread_id, data),
          UVM_FULL);
        void'(trek_c2t_message($time, thread_id, data));  ///@todo check return status?
        trek_backdoor_write64(valid_addr, 0, 0 /* debug */);
      end
    end
  endfunction: trek_poll_mbox

  // Try to start TrekSoc at time zero whenever this module is instanitated.
  // Unless you pass a +TREK_TBX_FILE=whatever.tbx, this should be benign.
  // In Verilator, you must call "start_tbx()" manually...
`ifndef VERILATOR
  initial begin: always_try_to_start_trek
    string here;
    $sformat(here, "%m");
    if (trek_uvm_pkg::trek_uvm_module_instance.len()) begin: check
      trek_fatal_callback($sformatf(
         {"Multiple instances of the 'trek_uvm' module detected\n  ",
          trek_uvm_pkg::trek_uvm_module_instance, "\n  ", here}));
    end
    trek_uvm_pkg::trek_uvm_module_instance = here;
    start_tbx();
  end
`endif // ~VERILATOR

  // The User calls this method when their test bench is booted and ready
  // for TrekSoC to start. It ultimately wants a "trekbox events file", which
  // can be obtained on the call to this method, passed on the simulator
  // command line, or fetched from the uvm configuration database.
  task start_tbx();
    int     retval;
    string  tbxFile;
    string  entryAction;
`ifndef VERILATOR
    uvm_event e;
     
    // Start Trek in NON-REACTIVE-mode.
    if ($value$plusargs("TREK_ENTRY=%s", entryAction)) begin: non_reactive_mode
      e = trek_uvm_events::get("_trek_end_of_test");

      trek_info_callback($sformatf(
        "trek: Starting with +TREK_ENTRY=%s", entryAction),
        UVM_NONE);
      retval = trek_solver_begin({$urandom(), $urandom()}, 0);
      if (retval != 0) begin: e1
        trek_fatal_callback("trek_solver_begin() has returned non-zero.");
      end

      retval = trek_reactive_entry(entryAction);
      if (retval != 0) begin: e2
        trek_fatal_callback("trek_reactive_entry() has returned non-zero.");
      end

      trek_started <= 1'b1;
      trek_uvm_pkg::trek_started = 1'b1;

      e.wait_on(); // Block here and wait for data from Trek
      e.reset();
      if (!trek_uvm_events::end_of_test()) begin
         trek_fatal_callback("trek_reactive_entry() has returned but end_of_test() not set");
      end

      retval = trek_solver_end();
      if (retval != 0) begin: e3
        trek_fatal_callback("trek_solver_end() has returned non-zero.");
      end

      trek_uvm_events::clear();
    end: non_reactive_mode

    // Start Trek in TBX-mode.
    if ($value$plusargs("TREK_TBX_FILE=%s", tbxFile)) begin: tbx_mode

      trek_info_callback({"trek: Starting with +TREK_TBX_FILE=", tbxFile},
        UVM_NONE);

`ifndef VERILATOR
      trek_info_callback(
        "trek: Waiting for user to call trek_uvm_events::do_backdoor_init()...",
        UVM_LOW);
      // Wait here for the user to indicate that it is safe to begin
      // backdoor loading of memory.  Verilator doesn't wait, but requires
      // the user to manually call start_tbx() after time zero when safe.
      begin: wait_here
        uvm_event  e;
        e = trek_uvm_events::get("_trek_backdoor_init");
        e.wait_on();
        //e.reset();
      end
      trek_info_callback(
        "trek: ... got call to trek_uvm_events::do_backdoor_init()",
        UVM_LOW);
`endif // ~VERILATOR

      retval = trek_uvm_start_tbx(tbxFile,
                                  c2t_mboxes_base,
                                  sdv_threads,
                                  seed,
                                  0);
      if (retval != 0) begin: trek_cannot_start
        trek_fatal_callback(
          $sformatf("trek_uvm_start_tbx(\"%s\") has returned %0d.",
                    tbxFile, retval));
      end
      // NBA to quiet Verilator lint when called from sequential procedure
      trek_started <= 1'b1;
`ifndef VERILATOR
      trek_uvm_pkg::trek_started = 1'b1;
`endif
    end: tbx_mode

    // Start Trek in REACTIVE-mode.
    if ($value$plusargs("TREK_REACTIVE_ENTRY=%s", entryAction)) begin: reactive_mode
      e = trek_uvm_events::get("_trek_end_of_test");

      trek_info_callback($sformatf(
        "trek: Starting with +TREK_REACTIVE_ENTRY=%s", entryAction),
        UVM_NONE);

      fork begin
        retval = trek_solver_begin({$urandom(), $urandom()}, 1);
        if (retval != 0) begin: e1
          trek_fatal_callback("trek_solver_begin() has returned non-zero.");
        end

`ifndef VERILATOR
      trek_info_callback(
        "trek: Waiting for user to call trek_uvm_events::do_backdoor_init()...",
        UVM_LOW);
      // Wait here for the user to indicate that it is safe to begin
      // backdoor loading of memory.  Verilator doesn't wait, but requires
      // the user to manually call start_tbx() after time zero when safe.
      begin: wait_here
        uvm_event  e;
        e = trek_uvm_events::get("_trek_backdoor_init");
        e.wait_on();
        //e.reset();
      end
      trek_info_callback(
        "trek: ... got call to trek_uvm_events::do_backdoor_init()",
        UVM_LOW);
`endif

        retval = trek_reactive_entry(entryAction);
        if (retval != 0) begin: e2
          trek_fatal_callback("trek_reactive_entry() has returned non-zero.");
        end

        trek_started <= 1'b1;
        trek_uvm_pkg::trek_started = 1'b1;

        e.wait_on(); // Block here and wait for data from Trek
        e.reset();
        if (!trek_uvm_events::end_of_test()) begin
           trek_fatal_callback("trek_reactive_entry() has returned but end_of_test() not set");
        end

        retval = trek_solver_end();
        if (retval != 0) begin: e3
          trek_fatal_callback("trek_solver_end() has returned non-zero.");
        end
      end join_none // fork begin
       
    end: reactive_mode
`endif // VERILATOR
     
     // wait for any reactive calls 
     wait fork;

  endtask: start_tbx

  function static bit trek_is_c2t_event_addr(input longint unsigned address);
    return ((trek_started == 1'b1) &&
            ((address >= c2t_mboxes_base) &&
             (address < (c2t_mboxes_base + (sdv_threads * `TREK_C2T_MBOX_SIZE)))));
  endfunction : trek_is_c2t_event_addr

  // TrekSoC calls this method to inform the test bench that a transaction
  // is available for the 'testbench port' with the given "tb_path".
  function static void trek_tlm_avail_callback(input string tb_path = "UNKNOWN");
`ifdef VERILATOR
    // At this moment, VERILATOR only supports pure-SDV tests...
    trek_info_callback({"trek_tlm_avail_callback(", tb_path ,") called."}, UVM_HIGH);
`else // ~VERILATOR
    uvm_event e;

    // This call to get() will build a new event or return an existing one.
    e = trek_uvm_events::get(tb_path);

    if (e.is_on() && (trek_dpi_pkg::trek_done() == 0)) begin: slow_tb
      trek_fatal_callback(
        {"trek_tlm_avail_callback: Unserviced tb_path: ", tb_path});
    end

    trek_info_callback($sformatf(
        "trek_tlm_avail_callback: Notifying tb_path '%s' (%0d waiters)",
        tb_path, e.get_num_waiters()),
      UVM_FULL);

    e.trigger(); // Wake up all waiters. Stay "on" until the event is "reset()".
`endif // ~VERILATOR
  endfunction: trek_tlm_avail_callback

  function static void trek_end_of_test_callback();
    trek_finished = 1'b1;
`ifdef VERILATOR
    trek_info_callback("trek_end_of_test_callback() called, but unimplemented!", UVM_LOW);
`else
    trek_uvm_pkg::trek_finished = 1'b1;
    trek_uvm_events::set_end_of_test();
`endif
  endfunction

  // What time is it in this module scope?
  function static longint unsigned trek_get_time();
    return $time;
  endfunction

`ifndef TREK_DEFAULT_INFO_VERBOSITY
`define TREK_DEFAULT_INFO_VERBOSITY UVM_LOW
`endif

  // Issue an informational message.
  function static void trek_info_callback(input string s,
                                   uvm_verbosity v = `TREK_DEFAULT_INFO_VERBOSITY);
`ifdef VERILATOR
    $display("INFO(%0d): %s", $stime, s);
`else
    uvm_report_info("trek", s, v
      `ifdef UVM_POST_VERSION_1_1
        , .context_name("trek_uvm")
      `endif
    );
`endif
  endfunction

  // Issue a warning message.
  function static void trek_warn_callback(input string s);
`ifdef VERILATOR
    $display("WARNING(%0d): %s", $stime, s);
`else
    uvm_report_warning("trek", s
     `ifdef UVM_POST_VERSION_1_1
       , .context_name("trek_uvm")
     `endif
    );
`endif
  endfunction

  // Issue an error message.
  function static void trek_error_callback(input string s);
`ifdef VERILATOR
    $display("ERROR(%0d): %s", $stime, s);
`else
    uvm_report_error("trek", s
      `ifdef UVM_POST_VERSION_1_1
        , .context_name("trek_uvm")
      `endif
    );
`endif
  endfunction

  // Issue a fatal error message.
  function static void trek_fatal_callback(input string s);
`ifdef VERILATOR
    $display("FATAL(%0d): %s", $stime, s);
    $finish(0);
`else
    uvm_report_fatal("trek", s
      `ifdef UVM_POST_VERSION_1_1
        , .context_name("trek_uvm")
      `endif
    );
`endif
  endfunction

endmodule: trek_uvm

`endif // GUARD__TREK_UVM__SV
