// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_h_east
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_h_east (
    input  logic [686:0]  i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head,
    output logic          o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld,
    output logic [108:0]  o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head,
    output logic          o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld,
    output logic [108:0]  o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld,
    input  logic [146:0]  i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head,
    output logic          o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld,
    input  logic [146:0]  i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head,
    output logic          o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld,
    input  logic [182:0]  i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head,
    output logic          o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld,
    output logic [182:0]  o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld,
    output logic [686:0]  o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data,
    output logic          o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head,
    input  logic          i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail,
    output logic          o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld,
    input  logic [108:0]  i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld,
    output logic [146:0]  o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data,
    output logic          o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head,
    input  logic          i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy,
    output logic          o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail,
    output logic          o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld,
    input  logic [686:0]  i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld,
    output logic [182:0]  o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data,
    output logic          o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head,
    input  logic          i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail,
    output logic          o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld,
    input  logic [182:0]  i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld,
    output logic [686:0]  o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld,
    input  logic [108:0]  i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld,
    output logic [686:0]  o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld,
    input  logic [108:0]  i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld,
    output logic [146:0]  o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld,
    input  logic [686:0]  i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld,
    output logic [146:0]  o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld,
    input  logic [686:0]  i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld,
    output logic [182:0]  o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld,
    input  logic [182:0]  i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data,
    input  logic          i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head,
    output logic          o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy,
    input  logic          i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail,
    input  logic          i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld,
    output logic [108:0]  o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data,
    output logic          o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head,
    input  logic          i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy,
    output logic          o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail,
    output logic          o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld,
    input  logic [146:0]  i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data,
    input  logic          i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head,
    output logic          o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy,
    input  logic          i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail,
    input  logic          i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld,
    output logic [686:0]  o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data,
    output logic          o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head,
    input  logic          i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy,
    output logic          o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail,
    output logic          o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld,
    input  logic [182:0]  i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data,
    input  logic          i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head,
    output logic          o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy,
    input  logic          i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail,
    input  logic          i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld,
    output logic [182:0]  o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data,
    output logic          o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head,
    input  logic          i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy,
    output logic          o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail,
    output logic          o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld,
    input  wire           i_noc_clk,
    input  wire           i_noc_rst_n,
    input  logic          scan_en
);

    noc_art_h_east u_noc_art_h_east (
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Data(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data),
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Head(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head),
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Data(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Head(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Data(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Head(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Data(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Head(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Data(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Head(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Rdy(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Tail(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Vld(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Data(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Head(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Rdy(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Tail(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Vld(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Data(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Head(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Rdy(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Tail(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Vld(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Data(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Head(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Rdy(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Tail(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Vld(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Data(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Head(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Rdy(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Tail(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Vld(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Data(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Head(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Rdy(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Tail(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Vld(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Data(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Head(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Rdy(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Tail(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Vld(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Data(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Head(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Rdy(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Tail(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Vld(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Data(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Head(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Rdy(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Tail(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Vld(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Data(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Head(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Rdy(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Tail(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Vld(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Data(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Head(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Rdy(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Tail(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Vld(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Data(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Head(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Rdy(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Tail(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Vld(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Data(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Head(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Rdy(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Tail(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Vld(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Data(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Head(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Rdy(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Tail(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Vld(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Data(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Head(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Rdy(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Tail(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Vld(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Data(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Head(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Rdy(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Tail(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Vld(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Data(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Head(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Rdy(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Tail(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Vld(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Data(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Head(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Rdy(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Tail(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Vld(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Data(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Head(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Rdy(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Tail(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Vld(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Data(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Head(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Rdy(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Tail(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Vld(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Data(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Head(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Rdy(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Tail(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Vld(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Data(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Head(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Rdy(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Tail(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Vld(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Data(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Head(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Rdy(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Tail(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Vld(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Data(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Head(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Rdy(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Tail(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Vld(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld),
    .noc_clk(i_noc_clk),
    .noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
    );

endmodule
