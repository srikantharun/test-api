// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_ddr_east
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_ddr_east (
    output logic [182:0]                                 o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data,
    output logic                                         o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head,
    input  logic                                         i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy,
    output logic                                         o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail,
    output logic                                         o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld,
    input  logic [182:0]                                 i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data,
    input  logic                                         i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head,
    output logic                                         o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy,
    input  logic                                         i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail,
    input  logic                                         i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld,
    input  logic [398:0]                                 i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld,
    output logic [398:0]                                 o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld,
    input  logic [398:0]                                 i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld,
    output logic [398:0]                                 o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld,
    input  logic [398:0]                                 i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld,
    output logic [398:0]                                 o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld,
    input  logic [398:0]                                 i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld,
    output logic [398:0]                                 o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld,
    input  logic [182:0]                                 i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld,
    output logic [182:0]                                 o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head,
    input  logic                                         i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail,
    output logic                                         o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld,
    input  logic                                         i_l2_addr_mode_port_b0,
    input  logic                                         i_l2_addr_mode_port_b1,
    input  logic                                         i_l2_intr_mode_port_b0,
    input  logic                                         i_l2_intr_mode_port_b1,
    input  logic                                         i_lpddr_graph_addr_mode_port_b0,
    input  logic                                         i_lpddr_graph_addr_mode_port_b1,
    input  logic                                         i_lpddr_graph_intr_mode_port_b0,
    input  logic                                         i_lpddr_graph_intr_mode_port_b1,
    input  wire                                          i_lpddr_ppp_0_aon_clk,
    input  wire                                          i_lpddr_ppp_0_aon_rst_n,
    output logic                                         o_lpddr_ppp_0_cfg_pwr_idle_val,
    output logic                                         o_lpddr_ppp_0_cfg_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_0_cfg_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_0_clk,
    input  wire                                          i_lpddr_ppp_0_clken,
    output logic                                         o_lpddr_ppp_0_pwr_idle_val,
    output logic                                         o_lpddr_ppp_0_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_0_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_0_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t     o_lpddr_ppp_0_targ_cfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_0_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_0_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     i_lpddr_ppp_0_targ_cfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_0_targ_cfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_0_targ_cfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_0_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                   o_lpddr_ppp_0_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     o_lpddr_ppp_0_targ_cfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_0_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_0_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_0_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_0_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_0_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_0_targ_mt_axi_m_arlen,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_0_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_0_targ_mt_axi_m_arqos,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_0_targ_mt_axi_m_arsize,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_0_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_0_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_0_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_0_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_0_targ_mt_axi_m_awlen,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_0_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_0_targ_mt_axi_m_awqos,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_0_targ_mt_axi_m_awsize,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_0_targ_mt_axi_m_bid,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_0_targ_mt_axi_m_bresp,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       i_lpddr_ppp_0_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_0_targ_mt_axi_m_rid,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_rlast,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_0_targ_mt_axi_m_rresp,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       o_lpddr_ppp_0_targ_mt_axi_m_wdata,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_wlast,
    input  logic                                         i_lpddr_ppp_0_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t       o_lpddr_ppp_0_targ_mt_axi_m_wstrb,
    output logic                                         o_lpddr_ppp_0_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_lpddr_ppp_0_targ_syscfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_lpddr_ppp_0_targ_syscfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_0_targ_syscfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_0_targ_syscfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_lpddr_ppp_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_lpddr_ppp_0_targ_syscfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_0_targ_syscfg_apb_m_pwrite,
    input  wire                                          i_lpddr_ppp_1_aon_clk,
    input  wire                                          i_lpddr_ppp_1_aon_rst_n,
    output logic                                         o_lpddr_ppp_1_cfg_pwr_idle_val,
    output logic                                         o_lpddr_ppp_1_cfg_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_1_cfg_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_1_clk,
    input  wire                                          i_lpddr_ppp_1_clken,
    output logic                                         o_lpddr_ppp_1_pwr_idle_val,
    output logic                                         o_lpddr_ppp_1_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_1_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_1_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t     o_lpddr_ppp_1_targ_cfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_1_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_1_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     i_lpddr_ppp_1_targ_cfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_1_targ_cfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_1_targ_cfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_1_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                   o_lpddr_ppp_1_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     o_lpddr_ppp_1_targ_cfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_1_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_1_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_1_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_1_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_1_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_1_targ_mt_axi_m_arlen,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_1_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_1_targ_mt_axi_m_arqos,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_1_targ_mt_axi_m_arsize,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_1_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_1_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_1_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_1_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_1_targ_mt_axi_m_awlen,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_1_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_1_targ_mt_axi_m_awqos,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_1_targ_mt_axi_m_awsize,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_1_targ_mt_axi_m_bid,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_1_targ_mt_axi_m_bresp,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       i_lpddr_ppp_1_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_1_targ_mt_axi_m_rid,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_rlast,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_1_targ_mt_axi_m_rresp,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       o_lpddr_ppp_1_targ_mt_axi_m_wdata,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_wlast,
    input  logic                                         i_lpddr_ppp_1_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t       o_lpddr_ppp_1_targ_mt_axi_m_wstrb,
    output logic                                         o_lpddr_ppp_1_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_lpddr_ppp_1_targ_syscfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_lpddr_ppp_1_targ_syscfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_1_targ_syscfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_1_targ_syscfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_lpddr_ppp_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_lpddr_ppp_1_targ_syscfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_1_targ_syscfg_apb_m_pwrite,
    input  wire                                          i_lpddr_ppp_2_aon_clk,
    input  wire                                          i_lpddr_ppp_2_aon_rst_n,
    output logic                                         o_lpddr_ppp_2_cfg_pwr_idle_val,
    output logic                                         o_lpddr_ppp_2_cfg_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_2_cfg_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_2_clk,
    input  wire                                          i_lpddr_ppp_2_clken,
    output logic                                         o_lpddr_ppp_2_pwr_idle_val,
    output logic                                         o_lpddr_ppp_2_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_2_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_2_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t     o_lpddr_ppp_2_targ_cfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_2_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_2_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     i_lpddr_ppp_2_targ_cfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_2_targ_cfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_2_targ_cfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_2_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                   o_lpddr_ppp_2_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     o_lpddr_ppp_2_targ_cfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_2_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_2_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_2_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_2_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_2_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_2_targ_mt_axi_m_arlen,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_2_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_2_targ_mt_axi_m_arqos,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_2_targ_mt_axi_m_arsize,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_2_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_2_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_2_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_2_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_2_targ_mt_axi_m_awlen,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_2_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_2_targ_mt_axi_m_awqos,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_2_targ_mt_axi_m_awsize,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_2_targ_mt_axi_m_bid,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_2_targ_mt_axi_m_bresp,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       i_lpddr_ppp_2_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_2_targ_mt_axi_m_rid,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_rlast,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_2_targ_mt_axi_m_rresp,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       o_lpddr_ppp_2_targ_mt_axi_m_wdata,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_wlast,
    input  logic                                         i_lpddr_ppp_2_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t       o_lpddr_ppp_2_targ_mt_axi_m_wstrb,
    output logic                                         o_lpddr_ppp_2_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_lpddr_ppp_2_targ_syscfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_lpddr_ppp_2_targ_syscfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_2_targ_syscfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_2_targ_syscfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_lpddr_ppp_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_lpddr_ppp_2_targ_syscfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_2_targ_syscfg_apb_m_pwrite,
    input  wire                                          i_lpddr_ppp_3_aon_clk,
    input  wire                                          i_lpddr_ppp_3_aon_rst_n,
    output logic                                         o_lpddr_ppp_3_cfg_pwr_idle_val,
    output logic                                         o_lpddr_ppp_3_cfg_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_3_cfg_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_3_clk,
    input  wire                                          i_lpddr_ppp_3_clken,
    output logic                                         o_lpddr_ppp_3_pwr_idle_val,
    output logic                                         o_lpddr_ppp_3_pwr_idle_ack,
    input  logic                                         i_lpddr_ppp_3_pwr_idle_req,
    input  wire                                          i_lpddr_ppp_3_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t     o_lpddr_ppp_3_targ_cfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_3_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_3_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     i_lpddr_ppp_3_targ_cfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_3_targ_cfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_3_targ_cfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_3_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                   o_lpddr_ppp_3_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t     o_lpddr_ppp_3_targ_cfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_3_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_3_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_3_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_3_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_3_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_3_targ_mt_axi_m_arlen,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_3_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_3_targ_mt_axi_m_arqos,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_3_targ_mt_axi_m_arsize,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_lpddr_ppp_3_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_lpddr_ppp_3_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_lpddr_ppp_3_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         o_lpddr_ppp_3_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_lpddr_ppp_3_targ_mt_axi_m_awlen,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_lpddr_ppp_3_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_lpddr_ppp_3_targ_mt_axi_m_awqos,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_lpddr_ppp_3_targ_mt_axi_m_awsize,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_3_targ_mt_axi_m_bid,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_3_targ_mt_axi_m_bresp,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       i_lpddr_ppp_3_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t         i_lpddr_ppp_3_targ_mt_axi_m_rid,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_rlast,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_lpddr_ppp_3_targ_mt_axi_m_rresp,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t       o_lpddr_ppp_3_targ_mt_axi_m_wdata,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_wlast,
    input  logic                                         i_lpddr_ppp_3_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t       o_lpddr_ppp_3_targ_mt_axi_m_wstrb,
    output logic                                         o_lpddr_ppp_3_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_lpddr_ppp_3_targ_syscfg_apb_m_paddr,
    output logic                                         o_lpddr_ppp_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_lpddr_ppp_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_lpddr_ppp_3_targ_syscfg_apb_m_prdata,
    input  logic                                         i_lpddr_ppp_3_targ_syscfg_apb_m_pready,
    output logic                                         o_lpddr_ppp_3_targ_syscfg_apb_m_psel,
    input  logic                                         i_lpddr_ppp_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_lpddr_ppp_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_lpddr_ppp_3_targ_syscfg_apb_m_pwdata,
    output logic                                         o_lpddr_ppp_3_targ_syscfg_apb_m_pwrite,
    input  logic                                         i_lpddr_ppp_addr_mode_port_b0,
    input  logic                                         i_lpddr_ppp_addr_mode_port_b1,
    input  logic                                         i_lpddr_ppp_intr_mode_port_b0,
    input  logic                                         i_lpddr_ppp_intr_mode_port_b1,
    input  wire                                          i_noc_clk,
    input  wire                                          i_noc_rst_n,
    input  logic                                         scan_en,
    input  wire                                          i_soc_periph_aon_clk,
    input  wire                                          i_soc_periph_aon_rst_n,
    input  wire                                          i_soc_periph_clk,
    input  wire                                          i_soc_periph_clken,
    input  chip_pkg::chip_axi_addr_t                     i_soc_periph_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                          i_soc_periph_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                          i_soc_periph_init_lt_axi_s_arcache,
    input  soc_periph_pkg::soc_periph_init_lt_axi_id_t   i_soc_periph_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                            i_soc_periph_init_lt_axi_s_arlen,
    input  logic                                         i_soc_periph_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                           i_soc_periph_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                            i_soc_periph_init_lt_axi_s_arqos,
    output logic                                         o_soc_periph_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                           i_soc_periph_init_lt_axi_s_arsize,
    input  logic                                         i_soc_periph_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                     i_soc_periph_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                          i_soc_periph_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                          i_soc_periph_init_lt_axi_s_awcache,
    input  soc_periph_pkg::soc_periph_init_lt_axi_id_t   i_soc_periph_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                            i_soc_periph_init_lt_axi_s_awlen,
    input  logic                                         i_soc_periph_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                           i_soc_periph_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                            i_soc_periph_init_lt_axi_s_awqos,
    output logic                                         o_soc_periph_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                           i_soc_periph_init_lt_axi_s_awsize,
    input  logic                                         i_soc_periph_init_lt_axi_s_awvalid,
    output soc_periph_pkg::soc_periph_init_lt_axi_id_t   o_soc_periph_init_lt_axi_s_bid,
    input  logic                                         i_soc_periph_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                           o_soc_periph_init_lt_axi_s_bresp,
    output logic                                         o_soc_periph_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                  o_soc_periph_init_lt_axi_s_rdata,
    output soc_periph_pkg::soc_periph_init_lt_axi_id_t   o_soc_periph_init_lt_axi_s_rid,
    output logic                                         o_soc_periph_init_lt_axi_s_rlast,
    input  logic                                         i_soc_periph_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                           o_soc_periph_init_lt_axi_s_rresp,
    output logic                                         o_soc_periph_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                  i_soc_periph_init_lt_axi_s_wdata,
    input  logic                                         i_soc_periph_init_lt_axi_s_wlast,
    output logic                                         o_soc_periph_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                 i_soc_periph_init_lt_axi_s_wstrb,
    input  logic                                         i_soc_periph_init_lt_axi_s_wvalid,
    output logic                                         o_soc_periph_pwr_idle_val,
    output logic                                         o_soc_periph_pwr_idle_ack,
    input  logic                                         i_soc_periph_pwr_idle_req,
    input  wire                                          i_soc_periph_rst_n,
    output chip_pkg::chip_axi_addr_t                     o_soc_periph_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                          o_soc_periph_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                          o_soc_periph_targ_lt_axi_m_arcache,
    output soc_periph_pkg::soc_periph_targ_lt_axi_id_t   o_soc_periph_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                            o_soc_periph_targ_lt_axi_m_arlen,
    output logic                                         o_soc_periph_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                           o_soc_periph_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                            o_soc_periph_targ_lt_axi_m_arqos,
    input  logic                                         i_soc_periph_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                           o_soc_periph_targ_lt_axi_m_arsize,
    output logic                                         o_soc_periph_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                     o_soc_periph_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                          o_soc_periph_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                          o_soc_periph_targ_lt_axi_m_awcache,
    output soc_periph_pkg::soc_periph_targ_lt_axi_id_t   o_soc_periph_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                            o_soc_periph_targ_lt_axi_m_awlen,
    output logic                                         o_soc_periph_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                           o_soc_periph_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                            o_soc_periph_targ_lt_axi_m_awqos,
    input  logic                                         i_soc_periph_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                           o_soc_periph_targ_lt_axi_m_awsize,
    output logic                                         o_soc_periph_targ_lt_axi_m_awvalid,
    input  soc_periph_pkg::soc_periph_targ_lt_axi_id_t   i_soc_periph_targ_lt_axi_m_bid,
    output logic                                         o_soc_periph_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                           i_soc_periph_targ_lt_axi_m_bresp,
    input  logic                                         i_soc_periph_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                  i_soc_periph_targ_lt_axi_m_rdata,
    input  soc_periph_pkg::soc_periph_targ_lt_axi_id_t   i_soc_periph_targ_lt_axi_m_rid,
    input  logic                                         i_soc_periph_targ_lt_axi_m_rlast,
    output logic                                         o_soc_periph_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                           i_soc_periph_targ_lt_axi_m_rresp,
    input  logic                                         i_soc_periph_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                  o_soc_periph_targ_lt_axi_m_wdata,
    output logic                                         o_soc_periph_targ_lt_axi_m_wlast,
    input  logic                                         i_soc_periph_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                 o_soc_periph_targ_lt_axi_m_wstrb,
    output logic                                         o_soc_periph_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                  o_soc_periph_targ_syscfg_apb_m_paddr,
    output logic                                         o_soc_periph_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                       o_soc_periph_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t              i_soc_periph_targ_syscfg_apb_m_prdata,
    input  logic                                         i_soc_periph_targ_syscfg_apb_m_pready,
    output logic                                         o_soc_periph_targ_syscfg_apb_m_psel,
    input  logic                                         i_soc_periph_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t              o_soc_periph_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t              o_soc_periph_targ_syscfg_apb_m_pwdata,
    output logic                                         o_soc_periph_targ_syscfg_apb_m_pwrite
);

    // Automated Address MSB fix: extra nets declaration
    logic[40:0] lpddr_ppp_0_targ_mt_axi_m_araddr_msb_fixed;
    logic[40:0] lpddr_ppp_0_targ_mt_axi_m_awaddr_msb_fixed;
    logic[40:0] lpddr_ppp_1_targ_mt_axi_m_araddr_msb_fixed;
    logic[40:0] lpddr_ppp_1_targ_mt_axi_m_awaddr_msb_fixed;
    logic[40:0] lpddr_ppp_2_targ_mt_axi_m_araddr_msb_fixed;
    logic[40:0] lpddr_ppp_2_targ_mt_axi_m_awaddr_msb_fixed;
    logic[40:0] lpddr_ppp_3_targ_mt_axi_m_araddr_msb_fixed;
    logic[40:0] lpddr_ppp_3_targ_mt_axi_m_awaddr_msb_fixed;
    logic[40:0] soc_periph_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] soc_periph_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] soc_periph_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] soc_periph_targ_lt_axi_m_awaddr_msb_fixed;

    // Automated Address MSB fix: Initiator-side assignments to extend addresses by 1 bit
    noc_common_addr_msb_setter u_addr_msb_fix_soc_periph_init_lt (
        .i_axi_araddr_40b (i_soc_periph_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (soc_periph_init_lt_axi_s_araddr_msb_fixed)
    );
    assign soc_periph_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_soc_periph_init_lt_axi_s_awaddr};

    // Automated Address MSB fix: Target-side assignments to drop unused MSB
    assign o_lpddr_ppp_0_targ_mt_axi_m_araddr = lpddr_ppp_0_targ_mt_axi_m_araddr_msb_fixed[39:0];
    assign o_lpddr_ppp_0_targ_mt_axi_m_awaddr = lpddr_ppp_0_targ_mt_axi_m_awaddr_msb_fixed[39:0];
    assign o_lpddr_ppp_1_targ_mt_axi_m_araddr = lpddr_ppp_1_targ_mt_axi_m_araddr_msb_fixed[39:0];
    assign o_lpddr_ppp_1_targ_mt_axi_m_awaddr = lpddr_ppp_1_targ_mt_axi_m_awaddr_msb_fixed[39:0];
    assign o_lpddr_ppp_2_targ_mt_axi_m_araddr = lpddr_ppp_2_targ_mt_axi_m_araddr_msb_fixed[39:0];
    assign o_lpddr_ppp_2_targ_mt_axi_m_awaddr = lpddr_ppp_2_targ_mt_axi_m_awaddr_msb_fixed[39:0];
    assign o_lpddr_ppp_3_targ_mt_axi_m_araddr = lpddr_ppp_3_targ_mt_axi_m_araddr_msb_fixed[39:0];
    assign o_lpddr_ppp_3_targ_mt_axi_m_awaddr = lpddr_ppp_3_targ_mt_axi_m_awaddr_msb_fixed[39:0];
    assign o_soc_periph_targ_lt_axi_m_araddr = soc_periph_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_soc_periph_targ_lt_axi_m_awaddr = soc_periph_targ_lt_axi_m_awaddr_msb_fixed[39:0];


    noc_art_ddr_east u_noc_art_ddr_east (
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Data(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Head(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Rdy(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Tail(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Vld(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Data(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Head(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Rdy(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Tail(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Vld(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Data(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Head(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Rdy(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Tail(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Vld(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Data(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Head(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Rdy(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Tail(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Vld(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Data(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Head(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Rdy(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Tail(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Vld(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Data(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Head(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Rdy(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Tail(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Vld(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Data(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Head(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Rdy(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Tail(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Vld(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Data(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Head(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Rdy(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Tail(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Vld(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Data(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Head(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Rdy(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Tail(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Vld(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Data(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Head(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Rdy(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Tail(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Vld(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Data(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Head(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Rdy(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Tail(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Vld(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Data(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Head(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Rdy(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Tail(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Vld(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld),
    .l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .lpddr_ppp_0_aon_clk(i_lpddr_ppp_0_aon_clk),
    .lpddr_ppp_0_aon_rst_n(i_lpddr_ppp_0_aon_rst_n),
    .lpddr_ppp_0_cfg_pwr_Idle(o_lpddr_ppp_0_cfg_pwr_idle_val),
    .lpddr_ppp_0_cfg_pwr_IdleAck(o_lpddr_ppp_0_cfg_pwr_idle_ack),
    .lpddr_ppp_0_cfg_pwr_IdleReq(i_lpddr_ppp_0_cfg_pwr_idle_req),
    .lpddr_ppp_0_clk(i_lpddr_ppp_0_clk),
    .lpddr_ppp_0_clken(i_lpddr_ppp_0_clken),
    .lpddr_ppp_0_pwr_Idle(o_lpddr_ppp_0_pwr_idle_val),
    .lpddr_ppp_0_pwr_IdleAck(o_lpddr_ppp_0_pwr_idle_ack),
    .lpddr_ppp_0_pwr_IdleReq(i_lpddr_ppp_0_pwr_idle_req),
    .lpddr_ppp_0_rst_n(i_lpddr_ppp_0_rst_n),
    .lpddr_ppp_0_targ_cfg_PAddr(o_lpddr_ppp_0_targ_cfg_apb_m_paddr),
    .lpddr_ppp_0_targ_cfg_PEnable(o_lpddr_ppp_0_targ_cfg_apb_m_penable),
    .lpddr_ppp_0_targ_cfg_PProt(o_lpddr_ppp_0_targ_cfg_apb_m_pprot),
    .lpddr_ppp_0_targ_cfg_PRData(i_lpddr_ppp_0_targ_cfg_apb_m_prdata),
    .lpddr_ppp_0_targ_cfg_PReady(i_lpddr_ppp_0_targ_cfg_apb_m_pready),
    .lpddr_ppp_0_targ_cfg_PSel(o_lpddr_ppp_0_targ_cfg_apb_m_psel),
    .lpddr_ppp_0_targ_cfg_PSlvErr(i_lpddr_ppp_0_targ_cfg_apb_m_pslverr),
    .lpddr_ppp_0_targ_cfg_PStrb(o_lpddr_ppp_0_targ_cfg_apb_m_pstrb),
    .lpddr_ppp_0_targ_cfg_PWData(o_lpddr_ppp_0_targ_cfg_apb_m_pwdata),
    .lpddr_ppp_0_targ_cfg_PWrite(o_lpddr_ppp_0_targ_cfg_apb_m_pwrite),
    .lpddr_ppp_0_targ_mt_Ar_Addr(lpddr_ppp_0_targ_mt_axi_m_araddr_msb_fixed),
    .lpddr_ppp_0_targ_mt_Ar_Burst(o_lpddr_ppp_0_targ_mt_axi_m_arburst),
    .lpddr_ppp_0_targ_mt_Ar_Cache(o_lpddr_ppp_0_targ_mt_axi_m_arcache),
    .lpddr_ppp_0_targ_mt_Ar_Id(o_lpddr_ppp_0_targ_mt_axi_m_arid),
    .lpddr_ppp_0_targ_mt_Ar_Len(o_lpddr_ppp_0_targ_mt_axi_m_arlen),
    .lpddr_ppp_0_targ_mt_Ar_Lock(o_lpddr_ppp_0_targ_mt_axi_m_arlock),
    .lpddr_ppp_0_targ_mt_Ar_Prot(o_lpddr_ppp_0_targ_mt_axi_m_arprot),
    .lpddr_ppp_0_targ_mt_Ar_Qos(o_lpddr_ppp_0_targ_mt_axi_m_arqos),
    .lpddr_ppp_0_targ_mt_Ar_Ready(i_lpddr_ppp_0_targ_mt_axi_m_arready),
    .lpddr_ppp_0_targ_mt_Ar_Size(o_lpddr_ppp_0_targ_mt_axi_m_arsize),
    .lpddr_ppp_0_targ_mt_Ar_Valid(o_lpddr_ppp_0_targ_mt_axi_m_arvalid),
    .lpddr_ppp_0_targ_mt_Aw_Addr(lpddr_ppp_0_targ_mt_axi_m_awaddr_msb_fixed),
    .lpddr_ppp_0_targ_mt_Aw_Burst(o_lpddr_ppp_0_targ_mt_axi_m_awburst),
    .lpddr_ppp_0_targ_mt_Aw_Cache(o_lpddr_ppp_0_targ_mt_axi_m_awcache),
    .lpddr_ppp_0_targ_mt_Aw_Id(o_lpddr_ppp_0_targ_mt_axi_m_awid),
    .lpddr_ppp_0_targ_mt_Aw_Len(o_lpddr_ppp_0_targ_mt_axi_m_awlen),
    .lpddr_ppp_0_targ_mt_Aw_Lock(o_lpddr_ppp_0_targ_mt_axi_m_awlock),
    .lpddr_ppp_0_targ_mt_Aw_Prot(o_lpddr_ppp_0_targ_mt_axi_m_awprot),
    .lpddr_ppp_0_targ_mt_Aw_Qos(o_lpddr_ppp_0_targ_mt_axi_m_awqos),
    .lpddr_ppp_0_targ_mt_Aw_Ready(i_lpddr_ppp_0_targ_mt_axi_m_awready),
    .lpddr_ppp_0_targ_mt_Aw_Size(o_lpddr_ppp_0_targ_mt_axi_m_awsize),
    .lpddr_ppp_0_targ_mt_Aw_Valid(o_lpddr_ppp_0_targ_mt_axi_m_awvalid),
    .lpddr_ppp_0_targ_mt_B_Id(i_lpddr_ppp_0_targ_mt_axi_m_bid),
    .lpddr_ppp_0_targ_mt_B_Ready(o_lpddr_ppp_0_targ_mt_axi_m_bready),
    .lpddr_ppp_0_targ_mt_B_Resp(i_lpddr_ppp_0_targ_mt_axi_m_bresp),
    .lpddr_ppp_0_targ_mt_B_Valid(i_lpddr_ppp_0_targ_mt_axi_m_bvalid),
    .lpddr_ppp_0_targ_mt_R_Data(i_lpddr_ppp_0_targ_mt_axi_m_rdata),
    .lpddr_ppp_0_targ_mt_R_Id(i_lpddr_ppp_0_targ_mt_axi_m_rid),
    .lpddr_ppp_0_targ_mt_R_Last(i_lpddr_ppp_0_targ_mt_axi_m_rlast),
    .lpddr_ppp_0_targ_mt_R_Ready(o_lpddr_ppp_0_targ_mt_axi_m_rready),
    .lpddr_ppp_0_targ_mt_R_Resp(i_lpddr_ppp_0_targ_mt_axi_m_rresp),
    .lpddr_ppp_0_targ_mt_R_Valid(i_lpddr_ppp_0_targ_mt_axi_m_rvalid),
    .lpddr_ppp_0_targ_mt_W_Data(o_lpddr_ppp_0_targ_mt_axi_m_wdata),
    .lpddr_ppp_0_targ_mt_W_Last(o_lpddr_ppp_0_targ_mt_axi_m_wlast),
    .lpddr_ppp_0_targ_mt_W_Ready(i_lpddr_ppp_0_targ_mt_axi_m_wready),
    .lpddr_ppp_0_targ_mt_W_Strb(o_lpddr_ppp_0_targ_mt_axi_m_wstrb),
    .lpddr_ppp_0_targ_mt_W_Valid(o_lpddr_ppp_0_targ_mt_axi_m_wvalid),
    .lpddr_ppp_0_targ_syscfg_PAddr(o_lpddr_ppp_0_targ_syscfg_apb_m_paddr),
    .lpddr_ppp_0_targ_syscfg_PEnable(o_lpddr_ppp_0_targ_syscfg_apb_m_penable),
    .lpddr_ppp_0_targ_syscfg_PProt(o_lpddr_ppp_0_targ_syscfg_apb_m_pprot),
    .lpddr_ppp_0_targ_syscfg_PRData(i_lpddr_ppp_0_targ_syscfg_apb_m_prdata),
    .lpddr_ppp_0_targ_syscfg_PReady(i_lpddr_ppp_0_targ_syscfg_apb_m_pready),
    .lpddr_ppp_0_targ_syscfg_PSel(o_lpddr_ppp_0_targ_syscfg_apb_m_psel),
    .lpddr_ppp_0_targ_syscfg_PSlvErr(i_lpddr_ppp_0_targ_syscfg_apb_m_pslverr),
    .lpddr_ppp_0_targ_syscfg_PStrb(o_lpddr_ppp_0_targ_syscfg_apb_m_pstrb),
    .lpddr_ppp_0_targ_syscfg_PWData(o_lpddr_ppp_0_targ_syscfg_apb_m_pwdata),
    .lpddr_ppp_0_targ_syscfg_PWrite(o_lpddr_ppp_0_targ_syscfg_apb_m_pwrite),
    .lpddr_ppp_1_aon_clk(i_lpddr_ppp_1_aon_clk),
    .lpddr_ppp_1_aon_rst_n(i_lpddr_ppp_1_aon_rst_n),
    .lpddr_ppp_1_cfg_pwr_Idle(o_lpddr_ppp_1_cfg_pwr_idle_val),
    .lpddr_ppp_1_cfg_pwr_IdleAck(o_lpddr_ppp_1_cfg_pwr_idle_ack),
    .lpddr_ppp_1_cfg_pwr_IdleReq(i_lpddr_ppp_1_cfg_pwr_idle_req),
    .lpddr_ppp_1_clk(i_lpddr_ppp_1_clk),
    .lpddr_ppp_1_clken(i_lpddr_ppp_1_clken),
    .lpddr_ppp_1_pwr_Idle(o_lpddr_ppp_1_pwr_idle_val),
    .lpddr_ppp_1_pwr_IdleAck(o_lpddr_ppp_1_pwr_idle_ack),
    .lpddr_ppp_1_pwr_IdleReq(i_lpddr_ppp_1_pwr_idle_req),
    .lpddr_ppp_1_rst_n(i_lpddr_ppp_1_rst_n),
    .lpddr_ppp_1_targ_cfg_PAddr(o_lpddr_ppp_1_targ_cfg_apb_m_paddr),
    .lpddr_ppp_1_targ_cfg_PEnable(o_lpddr_ppp_1_targ_cfg_apb_m_penable),
    .lpddr_ppp_1_targ_cfg_PProt(o_lpddr_ppp_1_targ_cfg_apb_m_pprot),
    .lpddr_ppp_1_targ_cfg_PRData(i_lpddr_ppp_1_targ_cfg_apb_m_prdata),
    .lpddr_ppp_1_targ_cfg_PReady(i_lpddr_ppp_1_targ_cfg_apb_m_pready),
    .lpddr_ppp_1_targ_cfg_PSel(o_lpddr_ppp_1_targ_cfg_apb_m_psel),
    .lpddr_ppp_1_targ_cfg_PSlvErr(i_lpddr_ppp_1_targ_cfg_apb_m_pslverr),
    .lpddr_ppp_1_targ_cfg_PStrb(o_lpddr_ppp_1_targ_cfg_apb_m_pstrb),
    .lpddr_ppp_1_targ_cfg_PWData(o_lpddr_ppp_1_targ_cfg_apb_m_pwdata),
    .lpddr_ppp_1_targ_cfg_PWrite(o_lpddr_ppp_1_targ_cfg_apb_m_pwrite),
    .lpddr_ppp_1_targ_mt_Ar_Addr(lpddr_ppp_1_targ_mt_axi_m_araddr_msb_fixed),
    .lpddr_ppp_1_targ_mt_Ar_Burst(o_lpddr_ppp_1_targ_mt_axi_m_arburst),
    .lpddr_ppp_1_targ_mt_Ar_Cache(o_lpddr_ppp_1_targ_mt_axi_m_arcache),
    .lpddr_ppp_1_targ_mt_Ar_Id(o_lpddr_ppp_1_targ_mt_axi_m_arid),
    .lpddr_ppp_1_targ_mt_Ar_Len(o_lpddr_ppp_1_targ_mt_axi_m_arlen),
    .lpddr_ppp_1_targ_mt_Ar_Lock(o_lpddr_ppp_1_targ_mt_axi_m_arlock),
    .lpddr_ppp_1_targ_mt_Ar_Prot(o_lpddr_ppp_1_targ_mt_axi_m_arprot),
    .lpddr_ppp_1_targ_mt_Ar_Qos(o_lpddr_ppp_1_targ_mt_axi_m_arqos),
    .lpddr_ppp_1_targ_mt_Ar_Ready(i_lpddr_ppp_1_targ_mt_axi_m_arready),
    .lpddr_ppp_1_targ_mt_Ar_Size(o_lpddr_ppp_1_targ_mt_axi_m_arsize),
    .lpddr_ppp_1_targ_mt_Ar_Valid(o_lpddr_ppp_1_targ_mt_axi_m_arvalid),
    .lpddr_ppp_1_targ_mt_Aw_Addr(lpddr_ppp_1_targ_mt_axi_m_awaddr_msb_fixed),
    .lpddr_ppp_1_targ_mt_Aw_Burst(o_lpddr_ppp_1_targ_mt_axi_m_awburst),
    .lpddr_ppp_1_targ_mt_Aw_Cache(o_lpddr_ppp_1_targ_mt_axi_m_awcache),
    .lpddr_ppp_1_targ_mt_Aw_Id(o_lpddr_ppp_1_targ_mt_axi_m_awid),
    .lpddr_ppp_1_targ_mt_Aw_Len(o_lpddr_ppp_1_targ_mt_axi_m_awlen),
    .lpddr_ppp_1_targ_mt_Aw_Lock(o_lpddr_ppp_1_targ_mt_axi_m_awlock),
    .lpddr_ppp_1_targ_mt_Aw_Prot(o_lpddr_ppp_1_targ_mt_axi_m_awprot),
    .lpddr_ppp_1_targ_mt_Aw_Qos(o_lpddr_ppp_1_targ_mt_axi_m_awqos),
    .lpddr_ppp_1_targ_mt_Aw_Ready(i_lpddr_ppp_1_targ_mt_axi_m_awready),
    .lpddr_ppp_1_targ_mt_Aw_Size(o_lpddr_ppp_1_targ_mt_axi_m_awsize),
    .lpddr_ppp_1_targ_mt_Aw_Valid(o_lpddr_ppp_1_targ_mt_axi_m_awvalid),
    .lpddr_ppp_1_targ_mt_B_Id(i_lpddr_ppp_1_targ_mt_axi_m_bid),
    .lpddr_ppp_1_targ_mt_B_Ready(o_lpddr_ppp_1_targ_mt_axi_m_bready),
    .lpddr_ppp_1_targ_mt_B_Resp(i_lpddr_ppp_1_targ_mt_axi_m_bresp),
    .lpddr_ppp_1_targ_mt_B_Valid(i_lpddr_ppp_1_targ_mt_axi_m_bvalid),
    .lpddr_ppp_1_targ_mt_R_Data(i_lpddr_ppp_1_targ_mt_axi_m_rdata),
    .lpddr_ppp_1_targ_mt_R_Id(i_lpddr_ppp_1_targ_mt_axi_m_rid),
    .lpddr_ppp_1_targ_mt_R_Last(i_lpddr_ppp_1_targ_mt_axi_m_rlast),
    .lpddr_ppp_1_targ_mt_R_Ready(o_lpddr_ppp_1_targ_mt_axi_m_rready),
    .lpddr_ppp_1_targ_mt_R_Resp(i_lpddr_ppp_1_targ_mt_axi_m_rresp),
    .lpddr_ppp_1_targ_mt_R_Valid(i_lpddr_ppp_1_targ_mt_axi_m_rvalid),
    .lpddr_ppp_1_targ_mt_W_Data(o_lpddr_ppp_1_targ_mt_axi_m_wdata),
    .lpddr_ppp_1_targ_mt_W_Last(o_lpddr_ppp_1_targ_mt_axi_m_wlast),
    .lpddr_ppp_1_targ_mt_W_Ready(i_lpddr_ppp_1_targ_mt_axi_m_wready),
    .lpddr_ppp_1_targ_mt_W_Strb(o_lpddr_ppp_1_targ_mt_axi_m_wstrb),
    .lpddr_ppp_1_targ_mt_W_Valid(o_lpddr_ppp_1_targ_mt_axi_m_wvalid),
    .lpddr_ppp_1_targ_syscfg_PAddr(o_lpddr_ppp_1_targ_syscfg_apb_m_paddr),
    .lpddr_ppp_1_targ_syscfg_PEnable(o_lpddr_ppp_1_targ_syscfg_apb_m_penable),
    .lpddr_ppp_1_targ_syscfg_PProt(o_lpddr_ppp_1_targ_syscfg_apb_m_pprot),
    .lpddr_ppp_1_targ_syscfg_PRData(i_lpddr_ppp_1_targ_syscfg_apb_m_prdata),
    .lpddr_ppp_1_targ_syscfg_PReady(i_lpddr_ppp_1_targ_syscfg_apb_m_pready),
    .lpddr_ppp_1_targ_syscfg_PSel(o_lpddr_ppp_1_targ_syscfg_apb_m_psel),
    .lpddr_ppp_1_targ_syscfg_PSlvErr(i_lpddr_ppp_1_targ_syscfg_apb_m_pslverr),
    .lpddr_ppp_1_targ_syscfg_PStrb(o_lpddr_ppp_1_targ_syscfg_apb_m_pstrb),
    .lpddr_ppp_1_targ_syscfg_PWData(o_lpddr_ppp_1_targ_syscfg_apb_m_pwdata),
    .lpddr_ppp_1_targ_syscfg_PWrite(o_lpddr_ppp_1_targ_syscfg_apb_m_pwrite),
    .lpddr_ppp_2_aon_clk(i_lpddr_ppp_2_aon_clk),
    .lpddr_ppp_2_aon_rst_n(i_lpddr_ppp_2_aon_rst_n),
    .lpddr_ppp_2_cfg_pwr_Idle(o_lpddr_ppp_2_cfg_pwr_idle_val),
    .lpddr_ppp_2_cfg_pwr_IdleAck(o_lpddr_ppp_2_cfg_pwr_idle_ack),
    .lpddr_ppp_2_cfg_pwr_IdleReq(i_lpddr_ppp_2_cfg_pwr_idle_req),
    .lpddr_ppp_2_clk(i_lpddr_ppp_2_clk),
    .lpddr_ppp_2_clken(i_lpddr_ppp_2_clken),
    .lpddr_ppp_2_pwr_Idle(o_lpddr_ppp_2_pwr_idle_val),
    .lpddr_ppp_2_pwr_IdleAck(o_lpddr_ppp_2_pwr_idle_ack),
    .lpddr_ppp_2_pwr_IdleReq(i_lpddr_ppp_2_pwr_idle_req),
    .lpddr_ppp_2_rst_n(i_lpddr_ppp_2_rst_n),
    .lpddr_ppp_2_targ_cfg_PAddr(o_lpddr_ppp_2_targ_cfg_apb_m_paddr),
    .lpddr_ppp_2_targ_cfg_PEnable(o_lpddr_ppp_2_targ_cfg_apb_m_penable),
    .lpddr_ppp_2_targ_cfg_PProt(o_lpddr_ppp_2_targ_cfg_apb_m_pprot),
    .lpddr_ppp_2_targ_cfg_PRData(i_lpddr_ppp_2_targ_cfg_apb_m_prdata),
    .lpddr_ppp_2_targ_cfg_PReady(i_lpddr_ppp_2_targ_cfg_apb_m_pready),
    .lpddr_ppp_2_targ_cfg_PSel(o_lpddr_ppp_2_targ_cfg_apb_m_psel),
    .lpddr_ppp_2_targ_cfg_PSlvErr(i_lpddr_ppp_2_targ_cfg_apb_m_pslverr),
    .lpddr_ppp_2_targ_cfg_PStrb(o_lpddr_ppp_2_targ_cfg_apb_m_pstrb),
    .lpddr_ppp_2_targ_cfg_PWData(o_lpddr_ppp_2_targ_cfg_apb_m_pwdata),
    .lpddr_ppp_2_targ_cfg_PWrite(o_lpddr_ppp_2_targ_cfg_apb_m_pwrite),
    .lpddr_ppp_2_targ_mt_Ar_Addr(lpddr_ppp_2_targ_mt_axi_m_araddr_msb_fixed),
    .lpddr_ppp_2_targ_mt_Ar_Burst(o_lpddr_ppp_2_targ_mt_axi_m_arburst),
    .lpddr_ppp_2_targ_mt_Ar_Cache(o_lpddr_ppp_2_targ_mt_axi_m_arcache),
    .lpddr_ppp_2_targ_mt_Ar_Id(o_lpddr_ppp_2_targ_mt_axi_m_arid),
    .lpddr_ppp_2_targ_mt_Ar_Len(o_lpddr_ppp_2_targ_mt_axi_m_arlen),
    .lpddr_ppp_2_targ_mt_Ar_Lock(o_lpddr_ppp_2_targ_mt_axi_m_arlock),
    .lpddr_ppp_2_targ_mt_Ar_Prot(o_lpddr_ppp_2_targ_mt_axi_m_arprot),
    .lpddr_ppp_2_targ_mt_Ar_Qos(o_lpddr_ppp_2_targ_mt_axi_m_arqos),
    .lpddr_ppp_2_targ_mt_Ar_Ready(i_lpddr_ppp_2_targ_mt_axi_m_arready),
    .lpddr_ppp_2_targ_mt_Ar_Size(o_lpddr_ppp_2_targ_mt_axi_m_arsize),
    .lpddr_ppp_2_targ_mt_Ar_Valid(o_lpddr_ppp_2_targ_mt_axi_m_arvalid),
    .lpddr_ppp_2_targ_mt_Aw_Addr(lpddr_ppp_2_targ_mt_axi_m_awaddr_msb_fixed),
    .lpddr_ppp_2_targ_mt_Aw_Burst(o_lpddr_ppp_2_targ_mt_axi_m_awburst),
    .lpddr_ppp_2_targ_mt_Aw_Cache(o_lpddr_ppp_2_targ_mt_axi_m_awcache),
    .lpddr_ppp_2_targ_mt_Aw_Id(o_lpddr_ppp_2_targ_mt_axi_m_awid),
    .lpddr_ppp_2_targ_mt_Aw_Len(o_lpddr_ppp_2_targ_mt_axi_m_awlen),
    .lpddr_ppp_2_targ_mt_Aw_Lock(o_lpddr_ppp_2_targ_mt_axi_m_awlock),
    .lpddr_ppp_2_targ_mt_Aw_Prot(o_lpddr_ppp_2_targ_mt_axi_m_awprot),
    .lpddr_ppp_2_targ_mt_Aw_Qos(o_lpddr_ppp_2_targ_mt_axi_m_awqos),
    .lpddr_ppp_2_targ_mt_Aw_Ready(i_lpddr_ppp_2_targ_mt_axi_m_awready),
    .lpddr_ppp_2_targ_mt_Aw_Size(o_lpddr_ppp_2_targ_mt_axi_m_awsize),
    .lpddr_ppp_2_targ_mt_Aw_Valid(o_lpddr_ppp_2_targ_mt_axi_m_awvalid),
    .lpddr_ppp_2_targ_mt_B_Id(i_lpddr_ppp_2_targ_mt_axi_m_bid),
    .lpddr_ppp_2_targ_mt_B_Ready(o_lpddr_ppp_2_targ_mt_axi_m_bready),
    .lpddr_ppp_2_targ_mt_B_Resp(i_lpddr_ppp_2_targ_mt_axi_m_bresp),
    .lpddr_ppp_2_targ_mt_B_Valid(i_lpddr_ppp_2_targ_mt_axi_m_bvalid),
    .lpddr_ppp_2_targ_mt_R_Data(i_lpddr_ppp_2_targ_mt_axi_m_rdata),
    .lpddr_ppp_2_targ_mt_R_Id(i_lpddr_ppp_2_targ_mt_axi_m_rid),
    .lpddr_ppp_2_targ_mt_R_Last(i_lpddr_ppp_2_targ_mt_axi_m_rlast),
    .lpddr_ppp_2_targ_mt_R_Ready(o_lpddr_ppp_2_targ_mt_axi_m_rready),
    .lpddr_ppp_2_targ_mt_R_Resp(i_lpddr_ppp_2_targ_mt_axi_m_rresp),
    .lpddr_ppp_2_targ_mt_R_Valid(i_lpddr_ppp_2_targ_mt_axi_m_rvalid),
    .lpddr_ppp_2_targ_mt_W_Data(o_lpddr_ppp_2_targ_mt_axi_m_wdata),
    .lpddr_ppp_2_targ_mt_W_Last(o_lpddr_ppp_2_targ_mt_axi_m_wlast),
    .lpddr_ppp_2_targ_mt_W_Ready(i_lpddr_ppp_2_targ_mt_axi_m_wready),
    .lpddr_ppp_2_targ_mt_W_Strb(o_lpddr_ppp_2_targ_mt_axi_m_wstrb),
    .lpddr_ppp_2_targ_mt_W_Valid(o_lpddr_ppp_2_targ_mt_axi_m_wvalid),
    .lpddr_ppp_2_targ_syscfg_PAddr(o_lpddr_ppp_2_targ_syscfg_apb_m_paddr),
    .lpddr_ppp_2_targ_syscfg_PEnable(o_lpddr_ppp_2_targ_syscfg_apb_m_penable),
    .lpddr_ppp_2_targ_syscfg_PProt(o_lpddr_ppp_2_targ_syscfg_apb_m_pprot),
    .lpddr_ppp_2_targ_syscfg_PRData(i_lpddr_ppp_2_targ_syscfg_apb_m_prdata),
    .lpddr_ppp_2_targ_syscfg_PReady(i_lpddr_ppp_2_targ_syscfg_apb_m_pready),
    .lpddr_ppp_2_targ_syscfg_PSel(o_lpddr_ppp_2_targ_syscfg_apb_m_psel),
    .lpddr_ppp_2_targ_syscfg_PSlvErr(i_lpddr_ppp_2_targ_syscfg_apb_m_pslverr),
    .lpddr_ppp_2_targ_syscfg_PStrb(o_lpddr_ppp_2_targ_syscfg_apb_m_pstrb),
    .lpddr_ppp_2_targ_syscfg_PWData(o_lpddr_ppp_2_targ_syscfg_apb_m_pwdata),
    .lpddr_ppp_2_targ_syscfg_PWrite(o_lpddr_ppp_2_targ_syscfg_apb_m_pwrite),
    .lpddr_ppp_3_aon_clk(i_lpddr_ppp_3_aon_clk),
    .lpddr_ppp_3_aon_rst_n(i_lpddr_ppp_3_aon_rst_n),
    .lpddr_ppp_3_cfg_pwr_Idle(o_lpddr_ppp_3_cfg_pwr_idle_val),
    .lpddr_ppp_3_cfg_pwr_IdleAck(o_lpddr_ppp_3_cfg_pwr_idle_ack),
    .lpddr_ppp_3_cfg_pwr_IdleReq(i_lpddr_ppp_3_cfg_pwr_idle_req),
    .lpddr_ppp_3_clk(i_lpddr_ppp_3_clk),
    .lpddr_ppp_3_clken(i_lpddr_ppp_3_clken),
    .lpddr_ppp_3_pwr_Idle(o_lpddr_ppp_3_pwr_idle_val),
    .lpddr_ppp_3_pwr_IdleAck(o_lpddr_ppp_3_pwr_idle_ack),
    .lpddr_ppp_3_pwr_IdleReq(i_lpddr_ppp_3_pwr_idle_req),
    .lpddr_ppp_3_rst_n(i_lpddr_ppp_3_rst_n),
    .lpddr_ppp_3_targ_cfg_PAddr(o_lpddr_ppp_3_targ_cfg_apb_m_paddr),
    .lpddr_ppp_3_targ_cfg_PEnable(o_lpddr_ppp_3_targ_cfg_apb_m_penable),
    .lpddr_ppp_3_targ_cfg_PProt(o_lpddr_ppp_3_targ_cfg_apb_m_pprot),
    .lpddr_ppp_3_targ_cfg_PRData(i_lpddr_ppp_3_targ_cfg_apb_m_prdata),
    .lpddr_ppp_3_targ_cfg_PReady(i_lpddr_ppp_3_targ_cfg_apb_m_pready),
    .lpddr_ppp_3_targ_cfg_PSel(o_lpddr_ppp_3_targ_cfg_apb_m_psel),
    .lpddr_ppp_3_targ_cfg_PSlvErr(i_lpddr_ppp_3_targ_cfg_apb_m_pslverr),
    .lpddr_ppp_3_targ_cfg_PStrb(o_lpddr_ppp_3_targ_cfg_apb_m_pstrb),
    .lpddr_ppp_3_targ_cfg_PWData(o_lpddr_ppp_3_targ_cfg_apb_m_pwdata),
    .lpddr_ppp_3_targ_cfg_PWrite(o_lpddr_ppp_3_targ_cfg_apb_m_pwrite),
    .lpddr_ppp_3_targ_mt_Ar_Addr(lpddr_ppp_3_targ_mt_axi_m_araddr_msb_fixed),
    .lpddr_ppp_3_targ_mt_Ar_Burst(o_lpddr_ppp_3_targ_mt_axi_m_arburst),
    .lpddr_ppp_3_targ_mt_Ar_Cache(o_lpddr_ppp_3_targ_mt_axi_m_arcache),
    .lpddr_ppp_3_targ_mt_Ar_Id(o_lpddr_ppp_3_targ_mt_axi_m_arid),
    .lpddr_ppp_3_targ_mt_Ar_Len(o_lpddr_ppp_3_targ_mt_axi_m_arlen),
    .lpddr_ppp_3_targ_mt_Ar_Lock(o_lpddr_ppp_3_targ_mt_axi_m_arlock),
    .lpddr_ppp_3_targ_mt_Ar_Prot(o_lpddr_ppp_3_targ_mt_axi_m_arprot),
    .lpddr_ppp_3_targ_mt_Ar_Qos(o_lpddr_ppp_3_targ_mt_axi_m_arqos),
    .lpddr_ppp_3_targ_mt_Ar_Ready(i_lpddr_ppp_3_targ_mt_axi_m_arready),
    .lpddr_ppp_3_targ_mt_Ar_Size(o_lpddr_ppp_3_targ_mt_axi_m_arsize),
    .lpddr_ppp_3_targ_mt_Ar_Valid(o_lpddr_ppp_3_targ_mt_axi_m_arvalid),
    .lpddr_ppp_3_targ_mt_Aw_Addr(lpddr_ppp_3_targ_mt_axi_m_awaddr_msb_fixed),
    .lpddr_ppp_3_targ_mt_Aw_Burst(o_lpddr_ppp_3_targ_mt_axi_m_awburst),
    .lpddr_ppp_3_targ_mt_Aw_Cache(o_lpddr_ppp_3_targ_mt_axi_m_awcache),
    .lpddr_ppp_3_targ_mt_Aw_Id(o_lpddr_ppp_3_targ_mt_axi_m_awid),
    .lpddr_ppp_3_targ_mt_Aw_Len(o_lpddr_ppp_3_targ_mt_axi_m_awlen),
    .lpddr_ppp_3_targ_mt_Aw_Lock(o_lpddr_ppp_3_targ_mt_axi_m_awlock),
    .lpddr_ppp_3_targ_mt_Aw_Prot(o_lpddr_ppp_3_targ_mt_axi_m_awprot),
    .lpddr_ppp_3_targ_mt_Aw_Qos(o_lpddr_ppp_3_targ_mt_axi_m_awqos),
    .lpddr_ppp_3_targ_mt_Aw_Ready(i_lpddr_ppp_3_targ_mt_axi_m_awready),
    .lpddr_ppp_3_targ_mt_Aw_Size(o_lpddr_ppp_3_targ_mt_axi_m_awsize),
    .lpddr_ppp_3_targ_mt_Aw_Valid(o_lpddr_ppp_3_targ_mt_axi_m_awvalid),
    .lpddr_ppp_3_targ_mt_B_Id(i_lpddr_ppp_3_targ_mt_axi_m_bid),
    .lpddr_ppp_3_targ_mt_B_Ready(o_lpddr_ppp_3_targ_mt_axi_m_bready),
    .lpddr_ppp_3_targ_mt_B_Resp(i_lpddr_ppp_3_targ_mt_axi_m_bresp),
    .lpddr_ppp_3_targ_mt_B_Valid(i_lpddr_ppp_3_targ_mt_axi_m_bvalid),
    .lpddr_ppp_3_targ_mt_R_Data(i_lpddr_ppp_3_targ_mt_axi_m_rdata),
    .lpddr_ppp_3_targ_mt_R_Id(i_lpddr_ppp_3_targ_mt_axi_m_rid),
    .lpddr_ppp_3_targ_mt_R_Last(i_lpddr_ppp_3_targ_mt_axi_m_rlast),
    .lpddr_ppp_3_targ_mt_R_Ready(o_lpddr_ppp_3_targ_mt_axi_m_rready),
    .lpddr_ppp_3_targ_mt_R_Resp(i_lpddr_ppp_3_targ_mt_axi_m_rresp),
    .lpddr_ppp_3_targ_mt_R_Valid(i_lpddr_ppp_3_targ_mt_axi_m_rvalid),
    .lpddr_ppp_3_targ_mt_W_Data(o_lpddr_ppp_3_targ_mt_axi_m_wdata),
    .lpddr_ppp_3_targ_mt_W_Last(o_lpddr_ppp_3_targ_mt_axi_m_wlast),
    .lpddr_ppp_3_targ_mt_W_Ready(i_lpddr_ppp_3_targ_mt_axi_m_wready),
    .lpddr_ppp_3_targ_mt_W_Strb(o_lpddr_ppp_3_targ_mt_axi_m_wstrb),
    .lpddr_ppp_3_targ_mt_W_Valid(o_lpddr_ppp_3_targ_mt_axi_m_wvalid),
    .lpddr_ppp_3_targ_syscfg_PAddr(o_lpddr_ppp_3_targ_syscfg_apb_m_paddr),
    .lpddr_ppp_3_targ_syscfg_PEnable(o_lpddr_ppp_3_targ_syscfg_apb_m_penable),
    .lpddr_ppp_3_targ_syscfg_PProt(o_lpddr_ppp_3_targ_syscfg_apb_m_pprot),
    .lpddr_ppp_3_targ_syscfg_PRData(i_lpddr_ppp_3_targ_syscfg_apb_m_prdata),
    .lpddr_ppp_3_targ_syscfg_PReady(i_lpddr_ppp_3_targ_syscfg_apb_m_pready),
    .lpddr_ppp_3_targ_syscfg_PSel(o_lpddr_ppp_3_targ_syscfg_apb_m_psel),
    .lpddr_ppp_3_targ_syscfg_PSlvErr(i_lpddr_ppp_3_targ_syscfg_apb_m_pslverr),
    .lpddr_ppp_3_targ_syscfg_PStrb(o_lpddr_ppp_3_targ_syscfg_apb_m_pstrb),
    .lpddr_ppp_3_targ_syscfg_PWData(o_lpddr_ppp_3_targ_syscfg_apb_m_pwdata),
    .lpddr_ppp_3_targ_syscfg_PWrite(o_lpddr_ppp_3_targ_syscfg_apb_m_pwrite),
    .lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .noc_clk(i_noc_clk),
    .noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en),
    .soc_periph_aon_clk(i_soc_periph_aon_clk),
    .soc_periph_aon_rst_n(i_soc_periph_aon_rst_n),
    .soc_periph_clk(i_soc_periph_clk),
    .soc_periph_clken(i_soc_periph_clken),
    .soc_periph_init_lt_Ar_Addr(soc_periph_init_lt_axi_s_araddr_msb_fixed),
    .soc_periph_init_lt_Ar_Burst(i_soc_periph_init_lt_axi_s_arburst),
    .soc_periph_init_lt_Ar_Cache(i_soc_periph_init_lt_axi_s_arcache),
    .soc_periph_init_lt_Ar_Id(i_soc_periph_init_lt_axi_s_arid),
    .soc_periph_init_lt_Ar_Len(i_soc_periph_init_lt_axi_s_arlen),
    .soc_periph_init_lt_Ar_Lock(i_soc_periph_init_lt_axi_s_arlock),
    .soc_periph_init_lt_Ar_Prot(i_soc_periph_init_lt_axi_s_arprot),
    .soc_periph_init_lt_Ar_Qos(i_soc_periph_init_lt_axi_s_arqos),
    .soc_periph_init_lt_Ar_Ready(o_soc_periph_init_lt_axi_s_arready),
    .soc_periph_init_lt_Ar_Size(i_soc_periph_init_lt_axi_s_arsize),
    .soc_periph_init_lt_Ar_Valid(i_soc_periph_init_lt_axi_s_arvalid),
    .soc_periph_init_lt_Aw_Addr(soc_periph_init_lt_axi_s_awaddr_msb_fixed),
    .soc_periph_init_lt_Aw_Burst(i_soc_periph_init_lt_axi_s_awburst),
    .soc_periph_init_lt_Aw_Cache(i_soc_periph_init_lt_axi_s_awcache),
    .soc_periph_init_lt_Aw_Id(i_soc_periph_init_lt_axi_s_awid),
    .soc_periph_init_lt_Aw_Len(i_soc_periph_init_lt_axi_s_awlen),
    .soc_periph_init_lt_Aw_Lock(i_soc_periph_init_lt_axi_s_awlock),
    .soc_periph_init_lt_Aw_Prot(i_soc_periph_init_lt_axi_s_awprot),
    .soc_periph_init_lt_Aw_Qos(i_soc_periph_init_lt_axi_s_awqos),
    .soc_periph_init_lt_Aw_Ready(o_soc_periph_init_lt_axi_s_awready),
    .soc_periph_init_lt_Aw_Size(i_soc_periph_init_lt_axi_s_awsize),
    .soc_periph_init_lt_Aw_Valid(i_soc_periph_init_lt_axi_s_awvalid),
    .soc_periph_init_lt_B_Id(o_soc_periph_init_lt_axi_s_bid),
    .soc_periph_init_lt_B_Ready(i_soc_periph_init_lt_axi_s_bready),
    .soc_periph_init_lt_B_Resp(o_soc_periph_init_lt_axi_s_bresp),
    .soc_periph_init_lt_B_Valid(o_soc_periph_init_lt_axi_s_bvalid),
    .soc_periph_init_lt_R_Data(o_soc_periph_init_lt_axi_s_rdata),
    .soc_periph_init_lt_R_Id(o_soc_periph_init_lt_axi_s_rid),
    .soc_periph_init_lt_R_Last(o_soc_periph_init_lt_axi_s_rlast),
    .soc_periph_init_lt_R_Ready(i_soc_periph_init_lt_axi_s_rready),
    .soc_periph_init_lt_R_Resp(o_soc_periph_init_lt_axi_s_rresp),
    .soc_periph_init_lt_R_Valid(o_soc_periph_init_lt_axi_s_rvalid),
    .soc_periph_init_lt_W_Data(i_soc_periph_init_lt_axi_s_wdata),
    .soc_periph_init_lt_W_Last(i_soc_periph_init_lt_axi_s_wlast),
    .soc_periph_init_lt_W_Ready(o_soc_periph_init_lt_axi_s_wready),
    .soc_periph_init_lt_W_Strb(i_soc_periph_init_lt_axi_s_wstrb),
    .soc_periph_init_lt_W_Valid(i_soc_periph_init_lt_axi_s_wvalid),
    .soc_periph_pwr_Idle(o_soc_periph_pwr_idle_val),
    .soc_periph_pwr_IdleAck(o_soc_periph_pwr_idle_ack),
    .soc_periph_pwr_IdleReq(i_soc_periph_pwr_idle_req),
    .soc_periph_rst_n(i_soc_periph_rst_n),
    .soc_periph_targ_lt_Ar_Addr(soc_periph_targ_lt_axi_m_araddr_msb_fixed),
    .soc_periph_targ_lt_Ar_Burst(o_soc_periph_targ_lt_axi_m_arburst),
    .soc_periph_targ_lt_Ar_Cache(o_soc_periph_targ_lt_axi_m_arcache),
    .soc_periph_targ_lt_Ar_Id(o_soc_periph_targ_lt_axi_m_arid),
    .soc_periph_targ_lt_Ar_Len(o_soc_periph_targ_lt_axi_m_arlen),
    .soc_periph_targ_lt_Ar_Lock(o_soc_periph_targ_lt_axi_m_arlock),
    .soc_periph_targ_lt_Ar_Prot(o_soc_periph_targ_lt_axi_m_arprot),
    .soc_periph_targ_lt_Ar_Qos(o_soc_periph_targ_lt_axi_m_arqos),
    .soc_periph_targ_lt_Ar_Ready(i_soc_periph_targ_lt_axi_m_arready),
    .soc_periph_targ_lt_Ar_Size(o_soc_periph_targ_lt_axi_m_arsize),
    .soc_periph_targ_lt_Ar_Valid(o_soc_periph_targ_lt_axi_m_arvalid),
    .soc_periph_targ_lt_Aw_Addr(soc_periph_targ_lt_axi_m_awaddr_msb_fixed),
    .soc_periph_targ_lt_Aw_Burst(o_soc_periph_targ_lt_axi_m_awburst),
    .soc_periph_targ_lt_Aw_Cache(o_soc_periph_targ_lt_axi_m_awcache),
    .soc_periph_targ_lt_Aw_Id(o_soc_periph_targ_lt_axi_m_awid),
    .soc_periph_targ_lt_Aw_Len(o_soc_periph_targ_lt_axi_m_awlen),
    .soc_periph_targ_lt_Aw_Lock(o_soc_periph_targ_lt_axi_m_awlock),
    .soc_periph_targ_lt_Aw_Prot(o_soc_periph_targ_lt_axi_m_awprot),
    .soc_periph_targ_lt_Aw_Qos(o_soc_periph_targ_lt_axi_m_awqos),
    .soc_periph_targ_lt_Aw_Ready(i_soc_periph_targ_lt_axi_m_awready),
    .soc_periph_targ_lt_Aw_Size(o_soc_periph_targ_lt_axi_m_awsize),
    .soc_periph_targ_lt_Aw_Valid(o_soc_periph_targ_lt_axi_m_awvalid),
    .soc_periph_targ_lt_B_Id(i_soc_periph_targ_lt_axi_m_bid),
    .soc_periph_targ_lt_B_Ready(o_soc_periph_targ_lt_axi_m_bready),
    .soc_periph_targ_lt_B_Resp(i_soc_periph_targ_lt_axi_m_bresp),
    .soc_periph_targ_lt_B_Valid(i_soc_periph_targ_lt_axi_m_bvalid),
    .soc_periph_targ_lt_R_Data(i_soc_periph_targ_lt_axi_m_rdata),
    .soc_periph_targ_lt_R_Id(i_soc_periph_targ_lt_axi_m_rid),
    .soc_periph_targ_lt_R_Last(i_soc_periph_targ_lt_axi_m_rlast),
    .soc_periph_targ_lt_R_Ready(o_soc_periph_targ_lt_axi_m_rready),
    .soc_periph_targ_lt_R_Resp(i_soc_periph_targ_lt_axi_m_rresp),
    .soc_periph_targ_lt_R_Valid(i_soc_periph_targ_lt_axi_m_rvalid),
    .soc_periph_targ_lt_W_Data(o_soc_periph_targ_lt_axi_m_wdata),
    .soc_periph_targ_lt_W_Last(o_soc_periph_targ_lt_axi_m_wlast),
    .soc_periph_targ_lt_W_Ready(i_soc_periph_targ_lt_axi_m_wready),
    .soc_periph_targ_lt_W_Strb(o_soc_periph_targ_lt_axi_m_wstrb),
    .soc_periph_targ_lt_W_Valid(o_soc_periph_targ_lt_axi_m_wvalid),
    .soc_periph_targ_syscfg_PAddr(o_soc_periph_targ_syscfg_apb_m_paddr),
    .soc_periph_targ_syscfg_PEnable(o_soc_periph_targ_syscfg_apb_m_penable),
    .soc_periph_targ_syscfg_PProt(o_soc_periph_targ_syscfg_apb_m_pprot),
    .soc_periph_targ_syscfg_PRData(i_soc_periph_targ_syscfg_apb_m_prdata),
    .soc_periph_targ_syscfg_PReady(i_soc_periph_targ_syscfg_apb_m_pready),
    .soc_periph_targ_syscfg_PSel(o_soc_periph_targ_syscfg_apb_m_psel),
    .soc_periph_targ_syscfg_PSlvErr(i_soc_periph_targ_syscfg_apb_m_pslverr),
    .soc_periph_targ_syscfg_PStrb(o_soc_periph_targ_syscfg_apb_m_pstrb),
    .soc_periph_targ_syscfg_PWData(o_soc_periph_targ_syscfg_apb_m_pwdata),
    .soc_periph_targ_syscfg_PWrite(o_soc_periph_targ_syscfg_apb_m_pwrite)
);

endmodule
