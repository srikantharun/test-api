// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: {{ cookiecutter.author_full_name }} <{{ cookiecutter.author_email }}>

/// Bind SVA in {{ cookiecutter.design_name }}
///

bind {{ cookiecutter.design_name }} {{ cookiecutter.design_name }}_sva u_{{ cookiecutter.design_name }}_sva (.*);
