// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description:
// UVM Incrementors
// Pre-configured numeric package
// Provide and cover interesting values for numeric variables
// Owner: abond

// Package: axe_uvm_incrementor_pkg 
package axe_uvm_numeric_pkg;
  
    `include "uvm_macros.svh"
  
    import uvm_pkg::*;
  
    `include "axe_uvm_numeric.svh"
    `include "axe_uvm_distribution.svh"
endpackage : axe_uvm_numeric_pkg
