// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: andrew dickson <andrew.dickson@axelera.ai>


// tests for the soc management IP
//

`include "reset_gen_test.svh"
`include "clock_test.svh"
`include "memory_map_test.svh"
`include "rtc_test.svh"
`include "wtd_test.svh"
`include "tms_test.svh"
`include "otp_test.svh"
`include "kse_test.svh"
`include "pctl_test.svh"
`include "debugger_test.svh"
