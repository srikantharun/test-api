// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024



package trek_dpi_pkg;

`include "trek_dpi.sv"

endpackage: trek_dpi_pkg
