// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024


`ifndef GUARD__TREK_UVM_PKG__SV
`define GUARD__TREK_UVM_PKG__SV

// This package contains low-level import/export methods that are
//   used in communication with TrekSoC via DPI.
`include "trek_dpi_pkg.sv"

// This package contains sequence items defined for this particular
//   test bench.  It also includes a straightforward sequence that
//   you might use for delivery of these items from Trek to your DUT.
//
package trek_uvm_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import trek_dpi_pkg::*;

  // Information about ports defined in the PSS model
  //
  typedef struct {
    string pss_name;
    string port_base_type;
    string port_type;
    string primary_txn_type;
    string secondary_txn_type;
    string adapter_type;
    int    built;
  } PortInformation_t;

  static bit trek_started  = 1'b0;
  static bit trek_finished = 1'b0;
  static string trek_uvm_module_instance;

  static int unsigned numPorts = 1;

  static       PortInformation_t portInfo[string] = '{
  //      tb_path               pss_name           base_type                     port_type                   primary_txn      secondary_txn              adapter_type             built
     "trek_delay_port" : '{"trek_delay_port", "trek_master_port", "trek_master_port_delay_req_delay_req", "trek_delay_req", "trek_delay_req", "trek_delay_req_delay_req_adapter", 0}
  };

  `include "trek_port_helpers.sv"

  // Infrastructure common to most UVM testbenches
  //
  `include "trek_uvm_events.sv"
  `include "trek_tlm_adapter.sv"
  `include "trek_port_base.sv"
  `include "trek_check_port.sv"
  `include "trek_get_port.sv"
  `include "trek_master_port.sv"
  `include "trek_put_port.sv"

  // Enumeration datatypes defined in the default package within the PSS model
  //


  // Transaction datatypes defined in the default package within the PSS model
  //
  `include "trek_delay_req.sv"


  // Port specializations defined in the PSS model
  //
  `include "trek_master_port_delay_req_delay_req.sv"


  // [Optional] port instances
  //
  `ifndef TREK_NO_PORT_INSTANCES
  static trek_master_port_delay_req_delay_req  trek_delay_port = new("trek_delay_port");
  `endif

  // Adapter typedefs for ports required by the PSS model
  // Your testbench should create adapters for types your sequences use.
  //
  `include "trek_delay_req_delay_req_adapter.sv"

  `include "trek_mbox_wrapper.sv"

endpackage: trek_uvm_pkg


// This module contains import/export methods that are used to
//   communication with TrekSoC.  Since it imports the "trek_uvm_pkg"
//   defined above, it goes here at the bottom of this file.
//
`ifndef TREK_NO_MODULE_IN_TREK_UVM_PKG
`include "trek_uvm.sv"
`endif


`endif // GUARD__TREK_UVM_PKG__SV
