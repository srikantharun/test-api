// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_soc
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_soc_p (
  input logic [7:0] i_apu_init_tok_ocpl_s_maddr,
  input logic i_apu_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_apu_init_tok_ocpl_s_mdata,
  output logic  o_apu_init_tok_ocpl_s_scmdaccept,
  output logic  o_apu_pwr_tok_idle_val,
  output logic  o_apu_pwr_tok_idle_ack,
  input logic  i_apu_pwr_tok_idle_req,
  output logic [7:0] o_apu_targ_tok_ocpl_m_maddr,
  output logic o_apu_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_apu_targ_tok_ocpl_m_mdata,
  input logic  i_apu_targ_tok_ocpl_m_scmdaccept,
  input logic [41:0] i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld,

    input  wire                                     i_apu_aon_clk,
    input  wire                                     i_apu_aon_rst_n,
    input  chip_pkg::chip_axi_addr_t                i_apu_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_apu_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_apu_init_lt_axi_s_arcache,
    input  logic[9:0]                               i_apu_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_apu_init_lt_axi_s_arlen,
    input  logic                                    i_apu_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_apu_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_apu_init_lt_axi_s_arqos,
    output logic                                    o_apu_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_apu_init_lt_axi_s_arsize,
    input  logic                                    i_apu_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                i_apu_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_apu_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_apu_init_lt_axi_s_awcache,
    input  logic[9:0]                               i_apu_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_apu_init_lt_axi_s_awlen,
    input  logic                                    i_apu_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_apu_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_apu_init_lt_axi_s_awqos,
    output logic                                    o_apu_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_apu_init_lt_axi_s_awsize,
    input  logic                                    i_apu_init_lt_axi_s_awvalid,
    output logic[9:0]                               o_apu_init_lt_axi_s_bid,
    input  logic                                    i_apu_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_apu_init_lt_axi_s_bresp,
    output logic                                    o_apu_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t             o_apu_init_lt_axi_s_rdata,
    output logic[9:0]                               o_apu_init_lt_axi_s_rid,
    output logic                                    o_apu_init_lt_axi_s_rlast,
    input  logic                                    i_apu_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_apu_init_lt_axi_s_rresp,
    output logic                                    o_apu_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_apu_init_lt_axi_s_wdata,
    input  logic                                    i_apu_init_lt_axi_s_wlast,
    output logic                                    o_apu_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t            i_apu_init_lt_axi_s_wstrb,
    input  logic                                    i_apu_init_lt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_apu_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_apu_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_apu_init_mt_axi_s_arcache,
    input  logic[8:0]                               i_apu_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_apu_init_mt_axi_s_arlen,
    input  logic                                    i_apu_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_apu_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_apu_init_mt_axi_s_arqos,
    output logic                                    o_apu_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_apu_init_mt_axi_s_arsize,
    input  logic                                    i_apu_init_mt_axi_s_arvalid,
    output apu_pkg::apu_axi_mt_data_t               o_apu_init_mt_axi_s_rdata,
    output logic[8:0]                               o_apu_init_mt_axi_s_rid,
    output logic                                    o_apu_init_mt_axi_s_rlast,
    input  logic                                    i_apu_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_apu_init_mt_axi_s_rresp,
    output logic                                    o_apu_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_apu_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_apu_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_apu_init_mt_axi_s_awcache,
    input  logic[8:0]                               i_apu_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_apu_init_mt_axi_s_awlen,
    input  logic                                    i_apu_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_apu_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_apu_init_mt_axi_s_awqos,
    output logic                                    o_apu_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_apu_init_mt_axi_s_awsize,
    input  logic                                    i_apu_init_mt_axi_s_awvalid,
    output logic[8:0]                               o_apu_init_mt_axi_s_bid,
    input  logic                                    i_apu_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_apu_init_mt_axi_s_bresp,
    output logic                                    o_apu_init_mt_axi_s_bvalid,
    input  apu_pkg::apu_axi_mt_data_t               i_apu_init_mt_axi_s_wdata,
    input  logic                                    i_apu_init_mt_axi_s_wlast,
    output logic                                    o_apu_init_mt_axi_s_wready,
    input  apu_pkg::apu_axi_mt_wstrb_t              i_apu_init_mt_axi_s_wstrb,
    input  logic                                    i_apu_init_mt_axi_s_wvalid,
    output logic                                    o_apu_pwr_idle_val,
    output logic                                    o_apu_pwr_idle_ack,
    input  logic                                    i_apu_pwr_idle_req,
    output chip_pkg::chip_axi_addr_t                o_apu_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_apu_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_apu_targ_lt_axi_m_arcache,
    output logic[7:0]                               o_apu_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_apu_targ_lt_axi_m_arlen,
    output logic                                    o_apu_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_apu_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_apu_targ_lt_axi_m_arqos,
    input  logic                                    i_apu_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_apu_targ_lt_axi_m_arsize,
    output logic                                    o_apu_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_apu_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_apu_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_apu_targ_lt_axi_m_awcache,
    output logic[7:0]                               o_apu_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_apu_targ_lt_axi_m_awlen,
    output logic                                    o_apu_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_apu_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_apu_targ_lt_axi_m_awqos,
    input  logic                                    i_apu_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_apu_targ_lt_axi_m_awsize,
    output logic                                    o_apu_targ_lt_axi_m_awvalid,
    input  logic[7:0]                               i_apu_targ_lt_axi_m_bid,
    output logic                                    o_apu_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_apu_targ_lt_axi_m_bresp,
    input  logic                                    i_apu_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_apu_targ_lt_axi_m_rdata,
    input  logic[7:0]                               i_apu_targ_lt_axi_m_rid,
    input  logic                                    i_apu_targ_lt_axi_m_rlast,
    output logic                                    o_apu_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_apu_targ_lt_axi_m_rresp,
    input  logic                                    i_apu_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_apu_targ_lt_axi_m_wdata,
    output logic                                    o_apu_targ_lt_axi_m_wlast,
    input  logic                                    i_apu_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_apu_targ_lt_axi_m_wstrb,
    output logic                                    o_apu_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_apu_targ_syscfg_apb_m_paddr,
    output logic                                    o_apu_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_apu_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_apu_targ_syscfg_apb_m_prdata,
    input  logic                                    i_apu_targ_syscfg_apb_m_pready,
    output logic                                    o_apu_targ_syscfg_apb_m_psel,
    input  logic                                    i_apu_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_apu_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_apu_targ_syscfg_apb_m_pwdata,
    output logic                                    o_apu_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_apu_x_clk,
    input  wire                                     i_apu_x_clken,
    input  wire                                     i_apu_x_rst_n,
    input  wire                                     i_dcd_aon_clk,
    input  wire                                     i_dcd_aon_rst_n,
    input  wire                                     i_dcd_codec_clk,
    input  wire                                     i_dcd_codec_clken,
    input  wire                                     i_dcd_codec_rst_n,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_0_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_0_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_0_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_0_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_0_init_mt_axi_s_arlen,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_0_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_0_init_mt_axi_s_arqos,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_0_init_mt_axi_s_arsize,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_arvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_data_t    o_dcd_dec_0_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_0_init_mt_axi_s_rid,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_rlast,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_0_init_mt_axi_s_rresp,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_0_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_0_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_0_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_0_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_0_init_mt_axi_s_awlen,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_0_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_0_init_mt_axi_s_awqos,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_0_init_mt_axi_s_awsize,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_0_init_mt_axi_s_bid,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_0_init_mt_axi_s_bresp,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_bvalid,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_data_t    i_dcd_dec_0_init_mt_axi_s_wdata,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_wlast,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_wready,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_strb_t    i_dcd_dec_0_init_mt_axi_s_wstrb,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_1_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_1_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_1_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_1_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_1_init_mt_axi_s_arlen,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_1_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_1_init_mt_axi_s_arqos,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_1_init_mt_axi_s_arsize,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_arvalid,
    output dcd_pkg::dcd_dec_1_init_mt_axi_data_t    o_dcd_dec_1_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_1_init_mt_axi_s_rid,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_rlast,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_1_init_mt_axi_s_rresp,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_1_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_1_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_1_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_1_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_1_init_mt_axi_s_awlen,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_1_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_1_init_mt_axi_s_awqos,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_1_init_mt_axi_s_awsize,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_1_init_mt_axi_s_bid,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_1_init_mt_axi_s_bresp,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_bvalid,
    input  dcd_pkg::dcd_dec_1_init_mt_axi_data_t    i_dcd_dec_1_init_mt_axi_s_wdata,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_wlast,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_wready,
    input  dcd_pkg::dcd_dec_1_init_mt_axi_strb_t    i_dcd_dec_1_init_mt_axi_s_wstrb,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_2_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_2_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_2_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_2_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_2_init_mt_axi_s_arlen,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_2_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_2_init_mt_axi_s_arqos,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_2_init_mt_axi_s_arsize,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_arvalid,
    output logic [127:0]                            o_dcd_dec_2_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_2_init_mt_axi_s_rid,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_rlast,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_2_init_mt_axi_s_rresp,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_2_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_2_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_2_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_2_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_2_init_mt_axi_s_awlen,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_2_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_2_init_mt_axi_s_awqos,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_2_init_mt_axi_s_awsize,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_2_init_mt_axi_s_bid,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_2_init_mt_axi_s_bresp,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_bvalid,
    input  logic [127:0]                            i_dcd_dec_2_init_mt_axi_s_wdata,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_wlast,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_wready,
    input  logic [15:0]                             i_dcd_dec_2_init_mt_axi_s_wstrb,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_wvalid,
    input  wire                                     i_dcd_mcu_clk,
    input  wire                                     i_dcd_mcu_clken,
    input  chip_pkg::chip_axi_addr_t                i_dcd_mcu_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_dcd_mcu_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_dcd_mcu_init_lt_axi_s_arcache,
    input  dcd_pkg::dcd_mcu_init_lt_axi_id_t        i_dcd_mcu_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_dcd_mcu_init_lt_axi_s_arlen,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_dcd_mcu_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_dcd_mcu_init_lt_axi_s_arqos,
    output logic                                    o_dcd_mcu_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_dcd_mcu_init_lt_axi_s_arsize,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_arvalid,
    output dcd_pkg::dcd_mcu_init_lt_axi_data_t      o_dcd_mcu_init_lt_axi_s_rdata,
    output dcd_pkg::dcd_mcu_init_lt_axi_id_t        o_dcd_mcu_init_lt_axi_s_rid,
    output logic                                    o_dcd_mcu_init_lt_axi_s_rlast,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_dcd_mcu_init_lt_axi_s_rresp,
    output logic                                    o_dcd_mcu_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_mcu_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_dcd_mcu_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_dcd_mcu_init_lt_axi_s_awcache,
    input  dcd_pkg::dcd_mcu_init_lt_axi_id_t        i_dcd_mcu_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_dcd_mcu_init_lt_axi_s_awlen,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_dcd_mcu_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_dcd_mcu_init_lt_axi_s_awqos,
    output logic                                    o_dcd_mcu_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_dcd_mcu_init_lt_axi_s_awsize,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_awvalid,
    output dcd_pkg::dcd_mcu_init_lt_axi_id_t        o_dcd_mcu_init_lt_axi_s_bid,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_dcd_mcu_init_lt_axi_s_bresp,
    output logic                                    o_dcd_mcu_init_lt_axi_s_bvalid,
    input  dcd_pkg::dcd_mcu_init_lt_axi_data_t      i_dcd_mcu_init_lt_axi_s_wdata,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_wlast,
    output logic                                    o_dcd_mcu_init_lt_axi_s_wready,
    input  dcd_pkg::dcd_mcu_init_lt_axi_strb_t      i_dcd_mcu_init_lt_axi_s_wstrb,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_wvalid,
    output logic                                    o_dcd_mcu_pwr_idle_val,
    output logic                                    o_dcd_mcu_pwr_idle_ack,
    input  logic                                    i_dcd_mcu_pwr_idle_req,
    input  wire                                     i_dcd_mcu_rst_n,
    output logic                                    o_dcd_pwr_idle_val,
    output logic                                    o_dcd_pwr_idle_ack,
    input  logic                                    i_dcd_pwr_idle_req,
    output dcd_pkg::dcd_targ_cfg_apb_addr_t         o_dcd_targ_cfg_apb_m_paddr,
    output logic                                    o_dcd_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_dcd_targ_cfg_apb_m_pprot,
    input  dcd_pkg::dcd_targ_cfg_apb_data_t         i_dcd_targ_cfg_apb_m_prdata,
    input  logic                                    i_dcd_targ_cfg_apb_m_pready,
    output logic                                    o_dcd_targ_cfg_apb_m_psel,
    input  logic                                    i_dcd_targ_cfg_apb_m_pslverr,
    output dcd_pkg::dcd_targ_cfg_apb_strb_t         o_dcd_targ_cfg_apb_m_pstrb,
    output dcd_pkg::dcd_targ_cfg_apb_data_t         o_dcd_targ_cfg_apb_m_pwdata,
    output logic                                    o_dcd_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_syscfg_addr_t             o_dcd_targ_syscfg_apb_m_paddr,
    output logic                                    o_dcd_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_dcd_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_dcd_targ_syscfg_apb_m_prdata,
    input  logic                                    i_dcd_targ_syscfg_apb_m_pready,
    output logic                                    o_dcd_targ_syscfg_apb_m_psel,
    input  logic                                    i_dcd_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_dcd_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_dcd_targ_syscfg_apb_m_pwdata,
    output logic                                    o_dcd_targ_syscfg_apb_m_pwrite,
    input  logic [686:0]                            i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld,
    output logic [108:0]                            o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld,
    input  logic [686:0]                            i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld,
    output logic [108:0]                            o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld,
    input  logic [146:0]                            i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld,
    output logic [686:0]                            o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld,
    input  logic [146:0]                            i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld,
    output logic [686:0]                            o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld,
    input  logic [182:0]                            i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld,
    output logic [182:0]                            o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld,
    input  logic [182:0]                            i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data,
    input  logic                                    i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head,
    output logic                                    o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy,
    input  logic                                    i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail,
    input  logic                                    i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld,
    output logic [182:0]                            o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data,
    output logic                                    o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head,
    input  logic                                    i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy,
    output logic                                    o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail,
    output logic                                    o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld,
    output logic [398:0]                            o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld,
    input  logic [398:0]                            i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld,
    output logic [398:0]                            o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld,
    input  logic [398:0]                            i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld,
    output logic [398:0]                            o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld,
    input  logic [398:0]                            i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld,
    output logic [398:0]                            o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld,
    input  logic [398:0]                            i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld,
    output logic [182:0]                            o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld,
    input  logic [182:0]                            i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld,
    output logic [686:0]                            o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld,
    input  logic [108:0]                            i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld,
    output logic [146:0]                            o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld,
    input  logic [686:0]                            i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld,
    output logic [182:0]                            o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld,
    input  logic [182:0]                            i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld,
    input  logic                                    i_l2_addr_mode_port_b0,
    input  logic                                    i_l2_addr_mode_port_b1,
    input  logic                                    i_l2_intr_mode_port_b0,
    input  logic                                    i_l2_intr_mode_port_b1,
    input  logic                                    i_lpddr_graph_addr_mode_port_b0,
    input  logic                                    i_lpddr_graph_addr_mode_port_b1,
    input  logic                                    i_lpddr_graph_intr_mode_port_b0,
    input  logic                                    i_lpddr_graph_intr_mode_port_b1,
    input  logic                                    i_lpddr_ppp_addr_mode_port_b0,
    input  logic                                    i_lpddr_ppp_addr_mode_port_b1,
    input  logic                                    i_lpddr_ppp_intr_mode_port_b0,
    input  logic                                    i_lpddr_ppp_intr_mode_port_b1,
    input  wire                                     i_noc_clk,
    input  wire                                     i_noc_rst_n,
    input  wire                                     i_pcie_aon_clk,
    input  wire                                     i_pcie_aon_rst_n,
    input  wire                                     i_pcie_init_mt_clk,
    input  wire                                     i_pcie_init_mt_clken,
    output logic                                    o_pcie_init_mt_pwr_idle_val,
    output logic                                    o_pcie_init_mt_pwr_idle_ack,
    input  logic                                    i_pcie_init_mt_pwr_idle_req,
    input  chip_pkg::chip_axi_addr_t                i_pcie_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pcie_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pcie_init_mt_axi_s_arcache,
    input  pcie_pkg::pcie_init_mt_axi_id_t          i_pcie_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pcie_init_mt_axi_s_arlen,
    input  logic                                    i_pcie_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pcie_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_pcie_init_mt_axi_s_arqos,
    output logic                                    o_pcie_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pcie_init_mt_axi_s_arsize,
    input  logic                                    i_pcie_init_mt_axi_s_arvalid,
    output pcie_pkg::pcie_init_mt_axi_data_t        o_pcie_init_mt_axi_s_rdata,
    output pcie_pkg::pcie_init_mt_axi_id_t          o_pcie_init_mt_axi_s_rid,
    output logic                                    o_pcie_init_mt_axi_s_rlast,
    input  logic                                    i_pcie_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pcie_init_mt_axi_s_rresp,
    output logic                                    o_pcie_init_mt_axi_s_rvalid,
    input  wire                                     i_pcie_init_mt_rst_n,
    input  chip_pkg::chip_axi_addr_t                i_pcie_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pcie_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pcie_init_mt_axi_s_awcache,
    input  pcie_pkg::pcie_init_mt_axi_id_t          i_pcie_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pcie_init_mt_axi_s_awlen,
    input  logic                                    i_pcie_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pcie_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_pcie_init_mt_axi_s_awqos,
    output logic                                    o_pcie_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pcie_init_mt_axi_s_awsize,
    input  logic                                    i_pcie_init_mt_axi_s_awvalid,
    output pcie_pkg::pcie_init_mt_axi_id_t          o_pcie_init_mt_axi_s_bid,
    input  logic                                    i_pcie_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pcie_init_mt_axi_s_bresp,
    output logic                                    o_pcie_init_mt_axi_s_bvalid,
    input  pcie_pkg::pcie_init_mt_axi_data_t        i_pcie_init_mt_axi_s_wdata,
    input  logic                                    i_pcie_init_mt_axi_s_wlast,
    output logic                                    o_pcie_init_mt_axi_s_wready,
    input  pcie_pkg::pcie_init_mt_axi_strb_t        i_pcie_init_mt_axi_s_wstrb,
    input  logic                                    i_pcie_init_mt_axi_s_wvalid,
    output pcie_pkg::pcie_targ_cfg_apb3_addr_t      o_pcie_targ_cfg_apb_m_paddr,
    output logic                                    o_pcie_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_pcie_targ_cfg_apb_m_pprot,
    input  pcie_pkg::pcie_targ_cfg_apb3_data_t      i_pcie_targ_cfg_apb_m_prdata,
    input  logic                                    i_pcie_targ_cfg_apb_m_pready,
    output logic                                    o_pcie_targ_cfg_apb_m_psel,
    input  logic                                    i_pcie_targ_cfg_apb_m_pslverr,
    output logic [3:0]                              o_pcie_targ_cfg_apb_m_pstrb,
    output pcie_pkg::pcie_targ_cfg_apb3_data_t      o_pcie_targ_cfg_apb_m_pwdata,
    output logic                                    o_pcie_targ_cfg_apb_m_pwrite,
    input  wire                                     i_pcie_targ_cfg_clk,
    input  wire                                     i_pcie_targ_cfg_clken,
    output chip_pkg::chip_axi_addr_t                o_pcie_targ_cfg_dbi_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_pcie_targ_cfg_dbi_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_pcie_targ_cfg_dbi_axi_m_arcache,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_id_t     o_pcie_targ_cfg_dbi_axi_m_arid,
    output axi_pkg::axi_len_t                       o_pcie_targ_cfg_dbi_axi_m_arlen,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_pcie_targ_cfg_dbi_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_pcie_targ_cfg_dbi_axi_m_arqos,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_arready,
    output axi_pkg::axi_size_t                      o_pcie_targ_cfg_dbi_axi_m_arsize,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_pcie_targ_cfg_dbi_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_pcie_targ_cfg_dbi_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_pcie_targ_cfg_dbi_axi_m_awcache,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_id_t     o_pcie_targ_cfg_dbi_axi_m_awid,
    output axi_pkg::axi_len_t                       o_pcie_targ_cfg_dbi_axi_m_awlen,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_pcie_targ_cfg_dbi_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_pcie_targ_cfg_dbi_axi_m_awqos,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_awready,
    output axi_pkg::axi_size_t                      o_pcie_targ_cfg_dbi_axi_m_awsize,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_awvalid,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_id_t     i_pcie_targ_cfg_dbi_axi_m_bid,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_pcie_targ_cfg_dbi_axi_m_bresp,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_bvalid,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_data_t   i_pcie_targ_cfg_dbi_axi_m_rdata,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_id_t     i_pcie_targ_cfg_dbi_axi_m_rid,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_rlast,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_pcie_targ_cfg_dbi_axi_m_rresp,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_rvalid,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_data_t   o_pcie_targ_cfg_dbi_axi_m_wdata,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_wlast,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_wready,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_strb_t   o_pcie_targ_cfg_dbi_axi_m_wstrb,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_wvalid,
    input  wire                                     i_pcie_targ_cfg_dbi_clk,
    input  wire                                     i_pcie_targ_cfg_dbi_clken,
    output logic                                    o_pcie_targ_cfg_dbi_pwr_idle_val,
    output logic                                    o_pcie_targ_cfg_dbi_pwr_idle_ack,
    input  logic                                    i_pcie_targ_cfg_dbi_pwr_idle_req,
    input  wire                                     i_pcie_targ_cfg_dbi_rst_n,
    output logic                                    o_pcie_targ_cfg_pwr_idle_val,
    output logic                                    o_pcie_targ_cfg_pwr_idle_ack,
    input  logic                                    i_pcie_targ_cfg_pwr_idle_req,
    input  wire                                     i_pcie_targ_cfg_rst_n,
    input  wire                                     i_pcie_targ_mt_clk,
    input  wire                                     i_pcie_targ_mt_clken,
    output logic                                    o_pcie_targ_mt_pwr_idle_val,
    output logic                                    o_pcie_targ_mt_pwr_idle_ack,
    input  logic                                    i_pcie_targ_mt_pwr_idle_req,
    output chip_pkg::chip_axi_addr_t                o_pcie_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_pcie_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_pcie_targ_mt_axi_m_arcache,
    output pcie_pkg::pcie_targ_mt_axi_id_t          o_pcie_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_pcie_targ_mt_axi_m_arlen,
    output logic                                    o_pcie_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_pcie_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_pcie_targ_mt_axi_m_arqos,
    input  logic                                    i_pcie_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_pcie_targ_mt_axi_m_arsize,
    output logic                                    o_pcie_targ_mt_axi_m_arvalid,
    input  pcie_pkg::pcie_targ_mt_axi_data_t        i_pcie_targ_mt_axi_m_rdata,
    input  pcie_pkg::pcie_targ_mt_axi_id_t          i_pcie_targ_mt_axi_m_rid,
    input  logic                                    i_pcie_targ_mt_axi_m_rlast,
    output logic                                    o_pcie_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_pcie_targ_mt_axi_m_rresp,
    input  logic                                    i_pcie_targ_mt_axi_m_rvalid,
    input  wire                                     i_pcie_targ_mt_rst_n,
    output chip_pkg::chip_axi_addr_t                o_pcie_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_pcie_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_pcie_targ_mt_axi_m_awcache,
    output pcie_pkg::pcie_targ_mt_axi_id_t          o_pcie_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_pcie_targ_mt_axi_m_awlen,
    output logic                                    o_pcie_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_pcie_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_pcie_targ_mt_axi_m_awqos,
    input  logic                                    i_pcie_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_pcie_targ_mt_axi_m_awsize,
    output logic                                    o_pcie_targ_mt_axi_m_awvalid,
    input  pcie_pkg::pcie_targ_mt_axi_id_t          i_pcie_targ_mt_axi_m_bid,
    output logic                                    o_pcie_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_pcie_targ_mt_axi_m_bresp,
    input  logic                                    i_pcie_targ_mt_axi_m_bvalid,
    output pcie_pkg::pcie_targ_mt_axi_data_t        o_pcie_targ_mt_axi_m_wdata,
    output logic                                    o_pcie_targ_mt_axi_m_wlast,
    input  logic                                    i_pcie_targ_mt_axi_m_wready,
    output pcie_pkg::pcie_targ_mt_axi_strb_t        o_pcie_targ_mt_axi_m_wstrb,
    output logic                                    o_pcie_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_pcie_targ_syscfg_apb_m_paddr,
    output logic                                    o_pcie_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_pcie_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_pcie_targ_syscfg_apb_m_prdata,
    input  logic                                    i_pcie_targ_syscfg_apb_m_pready,
    output logic                                    o_pcie_targ_syscfg_apb_m_psel,
    input  logic                                    i_pcie_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_pcie_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_pcie_targ_syscfg_apb_m_pwdata,
    output logic                                    o_pcie_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_pve_0_aon_clk,
    input  wire                                     i_pve_0_aon_rst_n,
    input  wire                                     i_pve_0_clk,
    input  wire                                     i_pve_0_clken,
    input  chip_pkg::chip_axi_addr_t                i_pve_0_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pve_0_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pve_0_init_ht_axi_s_arcache,
    input  pve_pkg::pve_ht_axi_m_id_t               i_pve_0_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pve_0_init_ht_axi_s_arlen,
    input  logic                                    i_pve_0_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pve_0_init_ht_axi_s_arprot,
    output logic                                    o_pve_0_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pve_0_init_ht_axi_s_arsize,
    input  logic                                    i_pve_0_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t             o_pve_0_init_ht_axi_s_rdata,
    output pve_pkg::pve_ht_axi_m_id_t               o_pve_0_init_ht_axi_s_rid,
    output logic                                    o_pve_0_init_ht_axi_s_rlast,
    input  logic                                    i_pve_0_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pve_0_init_ht_axi_s_rresp,
    output logic                                    o_pve_0_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_0_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pve_0_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pve_0_init_ht_axi_s_awcache,
    input  pve_pkg::pve_ht_axi_m_id_t               i_pve_0_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pve_0_init_ht_axi_s_awlen,
    input  logic                                    i_pve_0_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pve_0_init_ht_axi_s_awprot,
    output logic                                    o_pve_0_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pve_0_init_ht_axi_s_awsize,
    input  logic                                    i_pve_0_init_ht_axi_s_awvalid,
    output pve_pkg::pve_ht_axi_m_id_t               o_pve_0_init_ht_axi_s_bid,
    input  logic                                    i_pve_0_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pve_0_init_ht_axi_s_bresp,
    output logic                                    o_pve_0_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t             i_pve_0_init_ht_axi_s_wdata,
    input  logic                                    i_pve_0_init_ht_axi_s_wlast,
    output logic                                    o_pve_0_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t            i_pve_0_init_ht_axi_s_wstrb,
    input  logic                                    i_pve_0_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_0_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pve_0_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pve_0_init_lt_axi_s_arcache,
    input  pve_pkg::pve_lt_axi_m_id_t               i_pve_0_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pve_0_init_lt_axi_s_arlen,
    input  logic                                    i_pve_0_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pve_0_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_pve_0_init_lt_axi_s_arqos,
    output logic                                    o_pve_0_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pve_0_init_lt_axi_s_arsize,
    input  logic                                    i_pve_0_init_lt_axi_s_arvalid,
    output chip_pkg::chip_axi_lt_data_t             o_pve_0_init_lt_axi_s_rdata,
    output pve_pkg::pve_lt_axi_m_id_t               o_pve_0_init_lt_axi_s_rid,
    output logic                                    o_pve_0_init_lt_axi_s_rlast,
    input  logic                                    i_pve_0_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pve_0_init_lt_axi_s_rresp,
    output logic                                    o_pve_0_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_0_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pve_0_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pve_0_init_lt_axi_s_awcache,
    input  pve_pkg::pve_lt_axi_m_id_t               i_pve_0_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pve_0_init_lt_axi_s_awlen,
    input  logic                                    i_pve_0_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pve_0_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_pve_0_init_lt_axi_s_awqos,
    output logic                                    o_pve_0_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pve_0_init_lt_axi_s_awsize,
    input  logic                                    i_pve_0_init_lt_axi_s_awvalid,
    output pve_pkg::pve_lt_axi_m_id_t               o_pve_0_init_lt_axi_s_bid,
    input  logic                                    i_pve_0_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pve_0_init_lt_axi_s_bresp,
    output logic                                    o_pve_0_init_lt_axi_s_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_pve_0_init_lt_axi_s_wdata,
    input  logic                                    i_pve_0_init_lt_axi_s_wlast,
    output logic                                    o_pve_0_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t            i_pve_0_init_lt_axi_s_wstrb,
    input  logic                                    i_pve_0_init_lt_axi_s_wvalid,
    output logic                                    o_pve_0_pwr_idle_val,
    output logic                                    o_pve_0_pwr_idle_ack,
    input  logic                                    i_pve_0_pwr_idle_req,
    input  wire                                     i_pve_0_rst_n,
    output chip_pkg::chip_axi_addr_t                o_pve_0_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_pve_0_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_pve_0_targ_lt_axi_m_arcache,
    output pve_pkg::pve_lt_axi_s_id_t               o_pve_0_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_pve_0_targ_lt_axi_m_arlen,
    output logic                                    o_pve_0_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_pve_0_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_pve_0_targ_lt_axi_m_arqos,
    input  logic                                    i_pve_0_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_pve_0_targ_lt_axi_m_arsize,
    output logic                                    o_pve_0_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_pve_0_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_pve_0_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_pve_0_targ_lt_axi_m_awcache,
    output pve_pkg::pve_lt_axi_s_id_t               o_pve_0_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_pve_0_targ_lt_axi_m_awlen,
    output logic                                    o_pve_0_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_pve_0_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_pve_0_targ_lt_axi_m_awqos,
    input  logic                                    i_pve_0_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_pve_0_targ_lt_axi_m_awsize,
    output logic                                    o_pve_0_targ_lt_axi_m_awvalid,
    input  pve_pkg::pve_lt_axi_s_id_t               i_pve_0_targ_lt_axi_m_bid,
    output logic                                    o_pve_0_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_pve_0_targ_lt_axi_m_bresp,
    input  logic                                    i_pve_0_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_pve_0_targ_lt_axi_m_rdata,
    input  pve_pkg::pve_lt_axi_s_id_t               i_pve_0_targ_lt_axi_m_rid,
    input  logic                                    i_pve_0_targ_lt_axi_m_rlast,
    output logic                                    o_pve_0_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_pve_0_targ_lt_axi_m_rresp,
    input  logic                                    i_pve_0_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_pve_0_targ_lt_axi_m_wdata,
    output logic                                    o_pve_0_targ_lt_axi_m_wlast,
    input  logic                                    i_pve_0_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_pve_0_targ_lt_axi_m_wstrb,
    output logic                                    o_pve_0_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_pve_0_targ_syscfg_apb_m_paddr,
    output logic                                    o_pve_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_pve_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_pve_0_targ_syscfg_apb_m_prdata,
    input  logic                                    i_pve_0_targ_syscfg_apb_m_pready,
    output logic                                    o_pve_0_targ_syscfg_apb_m_psel,
    input  logic                                    i_pve_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_pve_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_pve_0_targ_syscfg_apb_m_pwdata,
    output logic                                    o_pve_0_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_pve_1_aon_clk,
    input  wire                                     i_pve_1_aon_rst_n,
    input  wire                                     i_pve_1_clk,
    input  wire                                     i_pve_1_clken,
    input  chip_pkg::chip_axi_addr_t                i_pve_1_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pve_1_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pve_1_init_ht_axi_s_arcache,
    input  pve_pkg::pve_ht_axi_m_id_t               i_pve_1_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pve_1_init_ht_axi_s_arlen,
    input  logic                                    i_pve_1_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pve_1_init_ht_axi_s_arprot,
    output logic                                    o_pve_1_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pve_1_init_ht_axi_s_arsize,
    input  logic                                    i_pve_1_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t             o_pve_1_init_ht_axi_s_rdata,
    output pve_pkg::pve_ht_axi_m_id_t               o_pve_1_init_ht_axi_s_rid,
    output logic                                    o_pve_1_init_ht_axi_s_rlast,
    input  logic                                    i_pve_1_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pve_1_init_ht_axi_s_rresp,
    output logic                                    o_pve_1_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_1_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pve_1_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pve_1_init_ht_axi_s_awcache,
    input  pve_pkg::pve_ht_axi_m_id_t               i_pve_1_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pve_1_init_ht_axi_s_awlen,
    input  logic                                    i_pve_1_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pve_1_init_ht_axi_s_awprot,
    output logic                                    o_pve_1_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pve_1_init_ht_axi_s_awsize,
    input  logic                                    i_pve_1_init_ht_axi_s_awvalid,
    output pve_pkg::pve_ht_axi_m_id_t               o_pve_1_init_ht_axi_s_bid,
    input  logic                                    i_pve_1_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pve_1_init_ht_axi_s_bresp,
    output logic                                    o_pve_1_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t             i_pve_1_init_ht_axi_s_wdata,
    input  logic                                    i_pve_1_init_ht_axi_s_wlast,
    output logic                                    o_pve_1_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t            i_pve_1_init_ht_axi_s_wstrb,
    input  logic                                    i_pve_1_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_1_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pve_1_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pve_1_init_lt_axi_s_arcache,
    input  pve_pkg::pve_lt_axi_m_id_t               i_pve_1_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pve_1_init_lt_axi_s_arlen,
    input  logic                                    i_pve_1_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pve_1_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_pve_1_init_lt_axi_s_arqos,
    output logic                                    o_pve_1_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pve_1_init_lt_axi_s_arsize,
    input  logic                                    i_pve_1_init_lt_axi_s_arvalid,
    output chip_pkg::chip_axi_lt_data_t             o_pve_1_init_lt_axi_s_rdata,
    output pve_pkg::pve_lt_axi_m_id_t               o_pve_1_init_lt_axi_s_rid,
    output logic                                    o_pve_1_init_lt_axi_s_rlast,
    input  logic                                    i_pve_1_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pve_1_init_lt_axi_s_rresp,
    output logic                                    o_pve_1_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_1_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pve_1_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pve_1_init_lt_axi_s_awcache,
    input  pve_pkg::pve_lt_axi_m_id_t               i_pve_1_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pve_1_init_lt_axi_s_awlen,
    input  logic                                    i_pve_1_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pve_1_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_pve_1_init_lt_axi_s_awqos,
    output logic                                    o_pve_1_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pve_1_init_lt_axi_s_awsize,
    input  logic                                    i_pve_1_init_lt_axi_s_awvalid,
    output pve_pkg::pve_lt_axi_m_id_t               o_pve_1_init_lt_axi_s_bid,
    input  logic                                    i_pve_1_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pve_1_init_lt_axi_s_bresp,
    output logic                                    o_pve_1_init_lt_axi_s_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_pve_1_init_lt_axi_s_wdata,
    input  logic                                    i_pve_1_init_lt_axi_s_wlast,
    output logic                                    o_pve_1_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t            i_pve_1_init_lt_axi_s_wstrb,
    input  logic                                    i_pve_1_init_lt_axi_s_wvalid,
    output logic                                    o_pve_1_pwr_idle_val,
    output logic                                    o_pve_1_pwr_idle_ack,
    input  logic                                    i_pve_1_pwr_idle_req,
    input  wire                                     i_pve_1_rst_n,
    output chip_pkg::chip_axi_addr_t                o_pve_1_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_pve_1_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_pve_1_targ_lt_axi_m_arcache,
    output pve_pkg::pve_lt_axi_s_id_t               o_pve_1_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_pve_1_targ_lt_axi_m_arlen,
    output logic                                    o_pve_1_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_pve_1_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_pve_1_targ_lt_axi_m_arqos,
    input  logic                                    i_pve_1_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_pve_1_targ_lt_axi_m_arsize,
    output logic                                    o_pve_1_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_pve_1_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_pve_1_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_pve_1_targ_lt_axi_m_awcache,
    output pve_pkg::pve_lt_axi_s_id_t               o_pve_1_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_pve_1_targ_lt_axi_m_awlen,
    output logic                                    o_pve_1_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_pve_1_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_pve_1_targ_lt_axi_m_awqos,
    input  logic                                    i_pve_1_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_pve_1_targ_lt_axi_m_awsize,
    output logic                                    o_pve_1_targ_lt_axi_m_awvalid,
    input  pve_pkg::pve_lt_axi_s_id_t               i_pve_1_targ_lt_axi_m_bid,
    output logic                                    o_pve_1_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_pve_1_targ_lt_axi_m_bresp,
    input  logic                                    i_pve_1_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_pve_1_targ_lt_axi_m_rdata,
    input  pve_pkg::pve_lt_axi_s_id_t               i_pve_1_targ_lt_axi_m_rid,
    input  logic                                    i_pve_1_targ_lt_axi_m_rlast,
    output logic                                    o_pve_1_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_pve_1_targ_lt_axi_m_rresp,
    input  logic                                    i_pve_1_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_pve_1_targ_lt_axi_m_wdata,
    output logic                                    o_pve_1_targ_lt_axi_m_wlast,
    input  logic                                    i_pve_1_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_pve_1_targ_lt_axi_m_wstrb,
    output logic                                    o_pve_1_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_pve_1_targ_syscfg_apb_m_paddr,
    output logic                                    o_pve_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_pve_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_pve_1_targ_syscfg_apb_m_prdata,
    input  logic                                    i_pve_1_targ_syscfg_apb_m_pready,
    output logic                                    o_pve_1_targ_syscfg_apb_m_psel,
    input  logic                                    i_pve_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_pve_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_pve_1_targ_syscfg_apb_m_pwdata,
    output logic                                    o_pve_1_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_soc_mgmt_aon_clk,
    input  wire                                     i_soc_mgmt_aon_rst_n,
    input  wire                                     i_soc_mgmt_clk,
    input  wire                                     i_soc_mgmt_clken,
    input  chip_pkg::chip_axi_addr_t                i_soc_mgmt_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_soc_mgmt_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_soc_mgmt_init_lt_axi_s_arcache,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t     i_soc_mgmt_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_soc_mgmt_init_lt_axi_s_arlen,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_soc_mgmt_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_soc_mgmt_init_lt_axi_s_arqos,
    output logic                                    o_soc_mgmt_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_soc_mgmt_init_lt_axi_s_arsize,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                i_soc_mgmt_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_soc_mgmt_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_soc_mgmt_init_lt_axi_s_awcache,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t     i_soc_mgmt_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_soc_mgmt_init_lt_axi_s_awlen,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_soc_mgmt_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_soc_mgmt_init_lt_axi_s_awqos,
    output logic                                    o_soc_mgmt_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_soc_mgmt_init_lt_axi_s_awsize,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_awvalid,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t     o_soc_mgmt_init_lt_axi_s_bid,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_soc_mgmt_init_lt_axi_s_bresp,
    output logic                                    o_soc_mgmt_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t             o_soc_mgmt_init_lt_axi_s_rdata,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t     o_soc_mgmt_init_lt_axi_s_rid,
    output logic                                    o_soc_mgmt_init_lt_axi_s_rlast,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_soc_mgmt_init_lt_axi_s_rresp,
    output logic                                    o_soc_mgmt_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_soc_mgmt_init_lt_axi_s_wdata,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_wlast,
    output logic                                    o_soc_mgmt_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t            i_soc_mgmt_init_lt_axi_s_wstrb,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_wvalid,
    output logic                                    o_soc_mgmt_pwr_idle_val,
    output logic                                    o_soc_mgmt_pwr_idle_ack,
    input  logic                                    i_soc_mgmt_pwr_idle_req,
    input  wire                                     i_soc_mgmt_rst_n,
    output chip_pkg::chip_axi_addr_t                o_soc_mgmt_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_soc_mgmt_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_soc_mgmt_targ_lt_axi_m_arcache,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t     o_soc_mgmt_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_soc_mgmt_targ_lt_axi_m_arlen,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_soc_mgmt_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_soc_mgmt_targ_lt_axi_m_arqos,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_soc_mgmt_targ_lt_axi_m_arsize,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_soc_mgmt_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_soc_mgmt_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_soc_mgmt_targ_lt_axi_m_awcache,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t     o_soc_mgmt_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_soc_mgmt_targ_lt_axi_m_awlen,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_soc_mgmt_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_soc_mgmt_targ_lt_axi_m_awqos,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_soc_mgmt_targ_lt_axi_m_awsize,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_awvalid,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t     i_soc_mgmt_targ_lt_axi_m_bid,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_soc_mgmt_targ_lt_axi_m_bresp,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_soc_mgmt_targ_lt_axi_m_rdata,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t     i_soc_mgmt_targ_lt_axi_m_rid,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_rlast,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_soc_mgmt_targ_lt_axi_m_rresp,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_soc_mgmt_targ_lt_axi_m_wdata,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_wlast,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_soc_mgmt_targ_lt_axi_m_wstrb,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_soc_mgmt_syscfg_addr_t    o_soc_mgmt_targ_syscfg_apb_m_paddr,
    output logic                                    o_soc_mgmt_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_soc_mgmt_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_soc_mgmt_targ_syscfg_apb_m_prdata,
    input  logic                                    i_soc_mgmt_targ_syscfg_apb_m_pready,
    output logic                                    o_soc_mgmt_targ_syscfg_apb_m_psel,
    input  logic                                    i_soc_mgmt_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_soc_mgmt_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_soc_mgmt_targ_syscfg_apb_m_pwdata,
    output logic                                    o_soc_mgmt_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_sys_spm_aon_clk,
    input  wire                                     i_sys_spm_aon_rst_n,
    input  wire                                     i_sys_spm_clk,
    input  wire                                     i_sys_spm_clken,
    output logic                                    o_sys_spm_pwr_idle_val,
    output logic                                    o_sys_spm_pwr_idle_ack,
    input  logic                                    i_sys_spm_pwr_idle_req,
    input  wire                                     i_sys_spm_rst_n,
    output chip_pkg::chip_axi_addr_t                o_sys_spm_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_sys_spm_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_sys_spm_targ_lt_axi_m_arcache,
    output sys_spm_pkg::sys_spm_targ_lt_axi_id_t    o_sys_spm_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_sys_spm_targ_lt_axi_m_arlen,
    output logic                                    o_sys_spm_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_sys_spm_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_sys_spm_targ_lt_axi_m_arqos,
    input  logic                                    i_sys_spm_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_sys_spm_targ_lt_axi_m_arsize,
    output logic                                    o_sys_spm_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_sys_spm_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_sys_spm_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_sys_spm_targ_lt_axi_m_awcache,
    output sys_spm_pkg::sys_spm_targ_lt_axi_id_t    o_sys_spm_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_sys_spm_targ_lt_axi_m_awlen,
    output logic                                    o_sys_spm_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_sys_spm_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_sys_spm_targ_lt_axi_m_awqos,
    input  logic                                    i_sys_spm_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_sys_spm_targ_lt_axi_m_awsize,
    output logic                                    o_sys_spm_targ_lt_axi_m_awvalid,
    input  sys_spm_pkg::sys_spm_targ_lt_axi_id_t    i_sys_spm_targ_lt_axi_m_bid,
    output logic                                    o_sys_spm_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_sys_spm_targ_lt_axi_m_bresp,
    input  logic                                    i_sys_spm_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_sys_spm_targ_lt_axi_m_rdata,
    input  sys_spm_pkg::sys_spm_targ_lt_axi_id_t    i_sys_spm_targ_lt_axi_m_rid,
    input  logic                                    i_sys_spm_targ_lt_axi_m_rlast,
    output logic                                    o_sys_spm_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_sys_spm_targ_lt_axi_m_rresp,
    input  logic                                    i_sys_spm_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_sys_spm_targ_lt_axi_m_wdata,
    output logic                                    o_sys_spm_targ_lt_axi_m_wlast,
    input  logic                                    i_sys_spm_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_sys_spm_targ_lt_axi_m_wstrb,
    output logic                                    o_sys_spm_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_sys_spm_targ_syscfg_apb_m_paddr,
    output logic                                    o_sys_spm_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_sys_spm_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_sys_spm_targ_syscfg_apb_m_prdata,
    input  logic                                    i_sys_spm_targ_syscfg_apb_m_pready,
    output logic                                    o_sys_spm_targ_syscfg_apb_m_psel,
    input  logic                                    i_sys_spm_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_sys_spm_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_sys_spm_targ_syscfg_apb_m_pwdata,
    output logic                                    o_sys_spm_targ_syscfg_apb_m_pwrite,
    // DFT Interface
    input  wire           tck,
    input  wire           trst,
    input  logic          tms,
    input  logic          tdi,
    output logic          tdo_en,
    output logic          tdo,
    input  wire           test_clk,
    input  logic          test_mode,
    input  logic          edt_update,
    input  logic          scan_en,
    input  logic [30-1:0] scan_in,
    output logic [30-1:0] scan_out,
    input  wire            bisr_clk,
    input  wire            bisr_reset,
    input  logic           bisr_shift_en,
    input  logic           bisr_si,
    output logic           bisr_so
);

logic [2:0] apu_targ_tok_ocpl_m_mcmd_ext;
assign o_apu_targ_tok_ocpl_m_mcmd = apu_targ_tok_ocpl_m_mcmd_ext[0];


    // -- Automatically-generated Reset Synchronizers -- //
    wire sys_spm_aon_rst_n_synced;
    wire soc_mgmt_aon_rst_n_synced;
    wire pve_1_aon_rst_n_synced;
    wire pve_0_aon_rst_n_synced;
    wire pcie_aon_rst_n_synced;
    wire dcd_aon_rst_n_synced;
    wire apu_aon_rst_n_synced;

    // SYS SPM AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_sys_spm_aon_rst_n_sync (
        .i_clk          (i_sys_spm_aon_clk),
        .i_rst_n        (i_sys_spm_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (sys_spm_aon_rst_n_synced)
    );

    // SOC MGMT AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_soc_mgmt_aon_rst_n_sync (
        .i_clk          (i_soc_mgmt_aon_clk),
        .i_rst_n        (i_soc_mgmt_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (soc_mgmt_aon_rst_n_synced)
    );

    // PVE 1 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_pve_1_aon_rst_n_sync (
        .i_clk          (i_pve_1_aon_clk),
        .i_rst_n        (i_pve_1_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (pve_1_aon_rst_n_synced)
    );

    // PVE 0 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_pve_0_aon_rst_n_sync (
        .i_clk          (i_pve_0_aon_clk),
        .i_rst_n        (i_pve_0_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (pve_0_aon_rst_n_synced)
    );

    // PCIE AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_pcie_aon_rst_n_sync (
        .i_clk          (i_pcie_aon_clk),
        .i_rst_n        (i_pcie_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (pcie_aon_rst_n_synced)
    );

    // DCD AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_dcd_aon_rst_n_sync (
        .i_clk          (i_dcd_aon_clk),
        .i_rst_n        (i_dcd_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (dcd_aon_rst_n_synced)
    );

    // APU AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_apu_aon_rst_n_sync (
        .i_clk          (i_apu_aon_clk),
        .i_rst_n        (i_apu_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (apu_aon_rst_n_synced)
    );
    // -- Automatically-generated Memory Interface -- //
    localparam int unsigned MEM_INTERFACES = 30;

    axe_tcl_sram_pkg::impl_inp_t mem_impl_in;
    axe_tcl_sram_pkg::impl_oup_t mem_impl_out;
    axe_tcl_sram_pkg::impl_inp_t[MEM_INTERFACES-1:0] impl_to_mem;
    axe_tcl_sram_pkg::impl_oup_t[MEM_INTERFACES-1:0] impl_from_mem;

    logic mem_pde;
    logic mem_prn;
    logic mem_ret;

    // TODO(psarras; bronze; drive mem_pde by CSRs)
    assign mem_pde = '0;
    // TODO(psarras; bronze; connect mem_prn to CSRs)
    // assign CSR = mem_prn;
    // Wiring: 1st interface in the chain
    assign mem_impl_in = axe_tcl_sram_pkg::impl_inp_t'{
        ret: mem_ret,
        pde: mem_pde,
        se: scan_en,
        default: '0
    };
    // Wiring: Last interface in the chain
    assign mem_prn = mem_impl_out.prn;
    // Wiring: Intermediate interfaces
    axe_tcl_sram_cfg #(
        .NUM_SRAMS(MEM_INTERFACES)
    ) u_sram_cfg_impl (
        .i_s(mem_impl_in),
        .o_s(mem_impl_out),
        .o_m(impl_to_mem),
        .i_m(impl_from_mem)
    );

    noc_soc u_noc_soc (
    .i_apu_aon_clk(i_apu_aon_clk),
    .i_apu_aon_rst_n(apu_aon_rst_n_synced),
    .i_apu_init_lt_axi_s_araddr(i_apu_init_lt_axi_s_araddr),
    .i_apu_init_lt_axi_s_arburst(i_apu_init_lt_axi_s_arburst),
    .i_apu_init_lt_axi_s_arcache(i_apu_init_lt_axi_s_arcache),
    .i_apu_init_lt_axi_s_arid(i_apu_init_lt_axi_s_arid),
    .i_apu_init_lt_axi_s_arlen(i_apu_init_lt_axi_s_arlen),
    .i_apu_init_lt_axi_s_arlock(i_apu_init_lt_axi_s_arlock),
    .i_apu_init_lt_axi_s_arprot(i_apu_init_lt_axi_s_arprot),
    .i_apu_init_lt_axi_s_arqos(i_apu_init_lt_axi_s_arqos),
    .o_apu_init_lt_axi_s_arready(o_apu_init_lt_axi_s_arready),
    .i_apu_init_lt_axi_s_arsize(i_apu_init_lt_axi_s_arsize),
    .i_apu_init_lt_axi_s_arvalid(i_apu_init_lt_axi_s_arvalid),
    .i_apu_init_lt_axi_s_awaddr(i_apu_init_lt_axi_s_awaddr),
    .i_apu_init_lt_axi_s_awburst(i_apu_init_lt_axi_s_awburst),
    .i_apu_init_lt_axi_s_awcache(i_apu_init_lt_axi_s_awcache),
    .i_apu_init_lt_axi_s_awid(i_apu_init_lt_axi_s_awid),
    .i_apu_init_lt_axi_s_awlen(i_apu_init_lt_axi_s_awlen),
    .i_apu_init_lt_axi_s_awlock(i_apu_init_lt_axi_s_awlock),
    .i_apu_init_lt_axi_s_awprot(i_apu_init_lt_axi_s_awprot),
    .i_apu_init_lt_axi_s_awqos(i_apu_init_lt_axi_s_awqos),
    .o_apu_init_lt_axi_s_awready(o_apu_init_lt_axi_s_awready),
    .i_apu_init_lt_axi_s_awsize(i_apu_init_lt_axi_s_awsize),
    .i_apu_init_lt_axi_s_awvalid(i_apu_init_lt_axi_s_awvalid),
    .o_apu_init_lt_axi_s_bid(o_apu_init_lt_axi_s_bid),
    .i_apu_init_lt_axi_s_bready(i_apu_init_lt_axi_s_bready),
    .o_apu_init_lt_axi_s_bresp(o_apu_init_lt_axi_s_bresp),
    .o_apu_init_lt_axi_s_bvalid(o_apu_init_lt_axi_s_bvalid),
    .o_apu_init_lt_axi_s_rdata(o_apu_init_lt_axi_s_rdata),
    .o_apu_init_lt_axi_s_rid(o_apu_init_lt_axi_s_rid),
    .o_apu_init_lt_axi_s_rlast(o_apu_init_lt_axi_s_rlast),
    .i_apu_init_lt_axi_s_rready(i_apu_init_lt_axi_s_rready),
    .o_apu_init_lt_axi_s_rresp(o_apu_init_lt_axi_s_rresp),
    .o_apu_init_lt_axi_s_rvalid(o_apu_init_lt_axi_s_rvalid),
    .i_apu_init_lt_axi_s_wdata(i_apu_init_lt_axi_s_wdata),
    .i_apu_init_lt_axi_s_wlast(i_apu_init_lt_axi_s_wlast),
    .o_apu_init_lt_axi_s_wready(o_apu_init_lt_axi_s_wready),
    .i_apu_init_lt_axi_s_wstrb(i_apu_init_lt_axi_s_wstrb),
    .i_apu_init_lt_axi_s_wvalid(i_apu_init_lt_axi_s_wvalid),
    .i_apu_init_mt_axi_s_araddr(i_apu_init_mt_axi_s_araddr),
    .i_apu_init_mt_axi_s_arburst(i_apu_init_mt_axi_s_arburst),
    .i_apu_init_mt_axi_s_arcache(i_apu_init_mt_axi_s_arcache),
    .i_apu_init_mt_axi_s_arid(i_apu_init_mt_axi_s_arid),
    .i_apu_init_mt_axi_s_arlen(i_apu_init_mt_axi_s_arlen),
    .i_apu_init_mt_axi_s_arlock(i_apu_init_mt_axi_s_arlock),
    .i_apu_init_mt_axi_s_arprot(i_apu_init_mt_axi_s_arprot),
    .i_apu_init_mt_axi_s_arqos(i_apu_init_mt_axi_s_arqos),
    .o_apu_init_mt_axi_s_arready(o_apu_init_mt_axi_s_arready),
    .i_apu_init_mt_axi_s_arsize(i_apu_init_mt_axi_s_arsize),
    .i_apu_init_mt_axi_s_arvalid(i_apu_init_mt_axi_s_arvalid),
    .o_apu_init_mt_axi_s_rdata(o_apu_init_mt_axi_s_rdata),
    .o_apu_init_mt_axi_s_rid(o_apu_init_mt_axi_s_rid),
    .o_apu_init_mt_axi_s_rlast(o_apu_init_mt_axi_s_rlast),
    .i_apu_init_mt_axi_s_rready(i_apu_init_mt_axi_s_rready),
    .o_apu_init_mt_axi_s_rresp(o_apu_init_mt_axi_s_rresp),
    .o_apu_init_mt_axi_s_rvalid(o_apu_init_mt_axi_s_rvalid),
    .i_apu_init_mt_axi_s_awaddr(i_apu_init_mt_axi_s_awaddr),
    .i_apu_init_mt_axi_s_awburst(i_apu_init_mt_axi_s_awburst),
    .i_apu_init_mt_axi_s_awcache(i_apu_init_mt_axi_s_awcache),
    .i_apu_init_mt_axi_s_awid(i_apu_init_mt_axi_s_awid),
    .i_apu_init_mt_axi_s_awlen(i_apu_init_mt_axi_s_awlen),
    .i_apu_init_mt_axi_s_awlock(i_apu_init_mt_axi_s_awlock),
    .i_apu_init_mt_axi_s_awprot(i_apu_init_mt_axi_s_awprot),
    .i_apu_init_mt_axi_s_awqos(i_apu_init_mt_axi_s_awqos),
    .o_apu_init_mt_axi_s_awready(o_apu_init_mt_axi_s_awready),
    .i_apu_init_mt_axi_s_awsize(i_apu_init_mt_axi_s_awsize),
    .i_apu_init_mt_axi_s_awvalid(i_apu_init_mt_axi_s_awvalid),
    .o_apu_init_mt_axi_s_bid(o_apu_init_mt_axi_s_bid),
    .i_apu_init_mt_axi_s_bready(i_apu_init_mt_axi_s_bready),
    .o_apu_init_mt_axi_s_bresp(o_apu_init_mt_axi_s_bresp),
    .o_apu_init_mt_axi_s_bvalid(o_apu_init_mt_axi_s_bvalid),
    .i_apu_init_mt_axi_s_wdata(i_apu_init_mt_axi_s_wdata),
    .i_apu_init_mt_axi_s_wlast(i_apu_init_mt_axi_s_wlast),
    .o_apu_init_mt_axi_s_wready(o_apu_init_mt_axi_s_wready),
    .i_apu_init_mt_axi_s_wstrb(i_apu_init_mt_axi_s_wstrb),
    .i_apu_init_mt_axi_s_wvalid(i_apu_init_mt_axi_s_wvalid),
    .o_apu_pwr_idle_val(o_apu_pwr_idle_val),
    .o_apu_pwr_idle_ack(o_apu_pwr_idle_ack),
    .i_apu_pwr_idle_req(i_apu_pwr_idle_req),
    .o_apu_targ_lt_axi_m_araddr(o_apu_targ_lt_axi_m_araddr),
    .o_apu_targ_lt_axi_m_arburst(o_apu_targ_lt_axi_m_arburst),
    .o_apu_targ_lt_axi_m_arcache(o_apu_targ_lt_axi_m_arcache),
    .o_apu_targ_lt_axi_m_arid(o_apu_targ_lt_axi_m_arid),
    .o_apu_targ_lt_axi_m_arlen(o_apu_targ_lt_axi_m_arlen),
    .o_apu_targ_lt_axi_m_arlock(o_apu_targ_lt_axi_m_arlock),
    .o_apu_targ_lt_axi_m_arprot(o_apu_targ_lt_axi_m_arprot),
    .o_apu_targ_lt_axi_m_arqos(o_apu_targ_lt_axi_m_arqos),
    .i_apu_targ_lt_axi_m_arready(i_apu_targ_lt_axi_m_arready),
    .o_apu_targ_lt_axi_m_arsize(o_apu_targ_lt_axi_m_arsize),
    .o_apu_targ_lt_axi_m_arvalid(o_apu_targ_lt_axi_m_arvalid),
    .o_apu_targ_lt_axi_m_awaddr(o_apu_targ_lt_axi_m_awaddr),
    .o_apu_targ_lt_axi_m_awburst(o_apu_targ_lt_axi_m_awburst),
    .o_apu_targ_lt_axi_m_awcache(o_apu_targ_lt_axi_m_awcache),
    .o_apu_targ_lt_axi_m_awid(o_apu_targ_lt_axi_m_awid),
    .o_apu_targ_lt_axi_m_awlen(o_apu_targ_lt_axi_m_awlen),
    .o_apu_targ_lt_axi_m_awlock(o_apu_targ_lt_axi_m_awlock),
    .o_apu_targ_lt_axi_m_awprot(o_apu_targ_lt_axi_m_awprot),
    .o_apu_targ_lt_axi_m_awqos(o_apu_targ_lt_axi_m_awqos),
    .i_apu_targ_lt_axi_m_awready(i_apu_targ_lt_axi_m_awready),
    .o_apu_targ_lt_axi_m_awsize(o_apu_targ_lt_axi_m_awsize),
    .o_apu_targ_lt_axi_m_awvalid(o_apu_targ_lt_axi_m_awvalid),
    .i_apu_targ_lt_axi_m_bid(i_apu_targ_lt_axi_m_bid),
    .o_apu_targ_lt_axi_m_bready(o_apu_targ_lt_axi_m_bready),
    .i_apu_targ_lt_axi_m_bresp(i_apu_targ_lt_axi_m_bresp),
    .i_apu_targ_lt_axi_m_bvalid(i_apu_targ_lt_axi_m_bvalid),
    .i_apu_targ_lt_axi_m_rdata(i_apu_targ_lt_axi_m_rdata),
    .i_apu_targ_lt_axi_m_rid(i_apu_targ_lt_axi_m_rid),
    .i_apu_targ_lt_axi_m_rlast(i_apu_targ_lt_axi_m_rlast),
    .o_apu_targ_lt_axi_m_rready(o_apu_targ_lt_axi_m_rready),
    .i_apu_targ_lt_axi_m_rresp(i_apu_targ_lt_axi_m_rresp),
    .i_apu_targ_lt_axi_m_rvalid(i_apu_targ_lt_axi_m_rvalid),
    .o_apu_targ_lt_axi_m_wdata(o_apu_targ_lt_axi_m_wdata),
    .o_apu_targ_lt_axi_m_wlast(o_apu_targ_lt_axi_m_wlast),
    .i_apu_targ_lt_axi_m_wready(i_apu_targ_lt_axi_m_wready),
    .o_apu_targ_lt_axi_m_wstrb(o_apu_targ_lt_axi_m_wstrb),
    .o_apu_targ_lt_axi_m_wvalid(o_apu_targ_lt_axi_m_wvalid),
    .o_apu_targ_syscfg_apb_m_paddr(o_apu_targ_syscfg_apb_m_paddr),
    .o_apu_targ_syscfg_apb_m_penable(o_apu_targ_syscfg_apb_m_penable),
    .o_apu_targ_syscfg_apb_m_pprot(o_apu_targ_syscfg_apb_m_pprot),
    .i_apu_targ_syscfg_apb_m_prdata(i_apu_targ_syscfg_apb_m_prdata),
    .i_apu_targ_syscfg_apb_m_pready(i_apu_targ_syscfg_apb_m_pready),
    .o_apu_targ_syscfg_apb_m_psel(o_apu_targ_syscfg_apb_m_psel),
    .i_apu_targ_syscfg_apb_m_pslverr(i_apu_targ_syscfg_apb_m_pslverr),
    .o_apu_targ_syscfg_apb_m_pstrb(o_apu_targ_syscfg_apb_m_pstrb),
    .o_apu_targ_syscfg_apb_m_pwdata(o_apu_targ_syscfg_apb_m_pwdata),
    .o_apu_targ_syscfg_apb_m_pwrite(o_apu_targ_syscfg_apb_m_pwrite),
    .i_apu_x_clk(i_apu_x_clk),
    .i_apu_x_clken(i_apu_x_clken),
    .i_apu_x_rst_n(i_apu_x_rst_n),
    .i_dcd_aon_clk(i_dcd_aon_clk),
    .i_dcd_aon_rst_n(dcd_aon_rst_n_synced),
    .i_dcd_codec_clk(i_dcd_codec_clk),
    .i_dcd_codec_clken(i_dcd_codec_clken),
    .i_dcd_codec_rst_n(i_dcd_codec_rst_n),
    .i_dcd_dec_0_init_mt_axi_s_araddr(i_dcd_dec_0_init_mt_axi_s_araddr),
    .i_dcd_dec_0_init_mt_axi_s_arburst(i_dcd_dec_0_init_mt_axi_s_arburst),
    .i_dcd_dec_0_init_mt_axi_s_arcache(i_dcd_dec_0_init_mt_axi_s_arcache),
    .i_dcd_dec_0_init_mt_axi_s_arid(i_dcd_dec_0_init_mt_axi_s_arid),
    .i_dcd_dec_0_init_mt_axi_s_arlen(i_dcd_dec_0_init_mt_axi_s_arlen),
    .i_dcd_dec_0_init_mt_axi_s_arlock(i_dcd_dec_0_init_mt_axi_s_arlock),
    .i_dcd_dec_0_init_mt_axi_s_arprot(i_dcd_dec_0_init_mt_axi_s_arprot),
    .i_dcd_dec_0_init_mt_axi_s_arqos(i_dcd_dec_0_init_mt_axi_s_arqos),
    .o_dcd_dec_0_init_mt_axi_s_arready(o_dcd_dec_0_init_mt_axi_s_arready),
    .i_dcd_dec_0_init_mt_axi_s_arsize(i_dcd_dec_0_init_mt_axi_s_arsize),
    .i_dcd_dec_0_init_mt_axi_s_arvalid(i_dcd_dec_0_init_mt_axi_s_arvalid),
    .o_dcd_dec_0_init_mt_axi_s_rdata(o_dcd_dec_0_init_mt_axi_s_rdata),
    .o_dcd_dec_0_init_mt_axi_s_rid(o_dcd_dec_0_init_mt_axi_s_rid),
    .o_dcd_dec_0_init_mt_axi_s_rlast(o_dcd_dec_0_init_mt_axi_s_rlast),
    .i_dcd_dec_0_init_mt_axi_s_rready(i_dcd_dec_0_init_mt_axi_s_rready),
    .o_dcd_dec_0_init_mt_axi_s_rresp(o_dcd_dec_0_init_mt_axi_s_rresp),
    .o_dcd_dec_0_init_mt_axi_s_rvalid(o_dcd_dec_0_init_mt_axi_s_rvalid),
    .i_dcd_dec_0_init_mt_axi_s_awaddr(i_dcd_dec_0_init_mt_axi_s_awaddr),
    .i_dcd_dec_0_init_mt_axi_s_awburst(i_dcd_dec_0_init_mt_axi_s_awburst),
    .i_dcd_dec_0_init_mt_axi_s_awcache(i_dcd_dec_0_init_mt_axi_s_awcache),
    .i_dcd_dec_0_init_mt_axi_s_awid(i_dcd_dec_0_init_mt_axi_s_awid),
    .i_dcd_dec_0_init_mt_axi_s_awlen(i_dcd_dec_0_init_mt_axi_s_awlen),
    .i_dcd_dec_0_init_mt_axi_s_awlock(i_dcd_dec_0_init_mt_axi_s_awlock),
    .i_dcd_dec_0_init_mt_axi_s_awprot(i_dcd_dec_0_init_mt_axi_s_awprot),
    .i_dcd_dec_0_init_mt_axi_s_awqos(i_dcd_dec_0_init_mt_axi_s_awqos),
    .o_dcd_dec_0_init_mt_axi_s_awready(o_dcd_dec_0_init_mt_axi_s_awready),
    .i_dcd_dec_0_init_mt_axi_s_awsize(i_dcd_dec_0_init_mt_axi_s_awsize),
    .i_dcd_dec_0_init_mt_axi_s_awvalid(i_dcd_dec_0_init_mt_axi_s_awvalid),
    .o_dcd_dec_0_init_mt_axi_s_bid(o_dcd_dec_0_init_mt_axi_s_bid),
    .i_dcd_dec_0_init_mt_axi_s_bready(i_dcd_dec_0_init_mt_axi_s_bready),
    .o_dcd_dec_0_init_mt_axi_s_bresp(o_dcd_dec_0_init_mt_axi_s_bresp),
    .o_dcd_dec_0_init_mt_axi_s_bvalid(o_dcd_dec_0_init_mt_axi_s_bvalid),
    .i_dcd_dec_0_init_mt_axi_s_wdata(i_dcd_dec_0_init_mt_axi_s_wdata),
    .i_dcd_dec_0_init_mt_axi_s_wlast(i_dcd_dec_0_init_mt_axi_s_wlast),
    .o_dcd_dec_0_init_mt_axi_s_wready(o_dcd_dec_0_init_mt_axi_s_wready),
    .i_dcd_dec_0_init_mt_axi_s_wstrb(i_dcd_dec_0_init_mt_axi_s_wstrb),
    .i_dcd_dec_0_init_mt_axi_s_wvalid(i_dcd_dec_0_init_mt_axi_s_wvalid),
    .i_dcd_dec_1_init_mt_axi_s_araddr(i_dcd_dec_1_init_mt_axi_s_araddr),
    .i_dcd_dec_1_init_mt_axi_s_arburst(i_dcd_dec_1_init_mt_axi_s_arburst),
    .i_dcd_dec_1_init_mt_axi_s_arcache(i_dcd_dec_1_init_mt_axi_s_arcache),
    .i_dcd_dec_1_init_mt_axi_s_arid(i_dcd_dec_1_init_mt_axi_s_arid),
    .i_dcd_dec_1_init_mt_axi_s_arlen(i_dcd_dec_1_init_mt_axi_s_arlen),
    .i_dcd_dec_1_init_mt_axi_s_arlock(i_dcd_dec_1_init_mt_axi_s_arlock),
    .i_dcd_dec_1_init_mt_axi_s_arprot(i_dcd_dec_1_init_mt_axi_s_arprot),
    .i_dcd_dec_1_init_mt_axi_s_arqos(i_dcd_dec_1_init_mt_axi_s_arqos),
    .o_dcd_dec_1_init_mt_axi_s_arready(o_dcd_dec_1_init_mt_axi_s_arready),
    .i_dcd_dec_1_init_mt_axi_s_arsize(i_dcd_dec_1_init_mt_axi_s_arsize),
    .i_dcd_dec_1_init_mt_axi_s_arvalid(i_dcd_dec_1_init_mt_axi_s_arvalid),
    .o_dcd_dec_1_init_mt_axi_s_rdata(o_dcd_dec_1_init_mt_axi_s_rdata),
    .o_dcd_dec_1_init_mt_axi_s_rid(o_dcd_dec_1_init_mt_axi_s_rid),
    .o_dcd_dec_1_init_mt_axi_s_rlast(o_dcd_dec_1_init_mt_axi_s_rlast),
    .i_dcd_dec_1_init_mt_axi_s_rready(i_dcd_dec_1_init_mt_axi_s_rready),
    .o_dcd_dec_1_init_mt_axi_s_rresp(o_dcd_dec_1_init_mt_axi_s_rresp),
    .o_dcd_dec_1_init_mt_axi_s_rvalid(o_dcd_dec_1_init_mt_axi_s_rvalid),
    .i_dcd_dec_1_init_mt_axi_s_awaddr(i_dcd_dec_1_init_mt_axi_s_awaddr),
    .i_dcd_dec_1_init_mt_axi_s_awburst(i_dcd_dec_1_init_mt_axi_s_awburst),
    .i_dcd_dec_1_init_mt_axi_s_awcache(i_dcd_dec_1_init_mt_axi_s_awcache),
    .i_dcd_dec_1_init_mt_axi_s_awid(i_dcd_dec_1_init_mt_axi_s_awid),
    .i_dcd_dec_1_init_mt_axi_s_awlen(i_dcd_dec_1_init_mt_axi_s_awlen),
    .i_dcd_dec_1_init_mt_axi_s_awlock(i_dcd_dec_1_init_mt_axi_s_awlock),
    .i_dcd_dec_1_init_mt_axi_s_awprot(i_dcd_dec_1_init_mt_axi_s_awprot),
    .i_dcd_dec_1_init_mt_axi_s_awqos(i_dcd_dec_1_init_mt_axi_s_awqos),
    .o_dcd_dec_1_init_mt_axi_s_awready(o_dcd_dec_1_init_mt_axi_s_awready),
    .i_dcd_dec_1_init_mt_axi_s_awsize(i_dcd_dec_1_init_mt_axi_s_awsize),
    .i_dcd_dec_1_init_mt_axi_s_awvalid(i_dcd_dec_1_init_mt_axi_s_awvalid),
    .o_dcd_dec_1_init_mt_axi_s_bid(o_dcd_dec_1_init_mt_axi_s_bid),
    .i_dcd_dec_1_init_mt_axi_s_bready(i_dcd_dec_1_init_mt_axi_s_bready),
    .o_dcd_dec_1_init_mt_axi_s_bresp(o_dcd_dec_1_init_mt_axi_s_bresp),
    .o_dcd_dec_1_init_mt_axi_s_bvalid(o_dcd_dec_1_init_mt_axi_s_bvalid),
    .i_dcd_dec_1_init_mt_axi_s_wdata(i_dcd_dec_1_init_mt_axi_s_wdata),
    .i_dcd_dec_1_init_mt_axi_s_wlast(i_dcd_dec_1_init_mt_axi_s_wlast),
    .o_dcd_dec_1_init_mt_axi_s_wready(o_dcd_dec_1_init_mt_axi_s_wready),
    .i_dcd_dec_1_init_mt_axi_s_wstrb(i_dcd_dec_1_init_mt_axi_s_wstrb),
    .i_dcd_dec_1_init_mt_axi_s_wvalid(i_dcd_dec_1_init_mt_axi_s_wvalid),
    .i_dcd_dec_2_init_mt_axi_s_araddr(i_dcd_dec_2_init_mt_axi_s_araddr),
    .i_dcd_dec_2_init_mt_axi_s_arburst(i_dcd_dec_2_init_mt_axi_s_arburst),
    .i_dcd_dec_2_init_mt_axi_s_arcache(i_dcd_dec_2_init_mt_axi_s_arcache),
    .i_dcd_dec_2_init_mt_axi_s_arid(i_dcd_dec_2_init_mt_axi_s_arid),
    .i_dcd_dec_2_init_mt_axi_s_arlen(i_dcd_dec_2_init_mt_axi_s_arlen),
    .i_dcd_dec_2_init_mt_axi_s_arlock(i_dcd_dec_2_init_mt_axi_s_arlock),
    .i_dcd_dec_2_init_mt_axi_s_arprot(i_dcd_dec_2_init_mt_axi_s_arprot),
    .i_dcd_dec_2_init_mt_axi_s_arqos(i_dcd_dec_2_init_mt_axi_s_arqos),
    .o_dcd_dec_2_init_mt_axi_s_arready(o_dcd_dec_2_init_mt_axi_s_arready),
    .i_dcd_dec_2_init_mt_axi_s_arsize(i_dcd_dec_2_init_mt_axi_s_arsize),
    .i_dcd_dec_2_init_mt_axi_s_arvalid(i_dcd_dec_2_init_mt_axi_s_arvalid),
    .o_dcd_dec_2_init_mt_axi_s_rdata(o_dcd_dec_2_init_mt_axi_s_rdata),
    .o_dcd_dec_2_init_mt_axi_s_rid(o_dcd_dec_2_init_mt_axi_s_rid),
    .o_dcd_dec_2_init_mt_axi_s_rlast(o_dcd_dec_2_init_mt_axi_s_rlast),
    .i_dcd_dec_2_init_mt_axi_s_rready(i_dcd_dec_2_init_mt_axi_s_rready),
    .o_dcd_dec_2_init_mt_axi_s_rresp(o_dcd_dec_2_init_mt_axi_s_rresp),
    .o_dcd_dec_2_init_mt_axi_s_rvalid(o_dcd_dec_2_init_mt_axi_s_rvalid),
    .i_dcd_dec_2_init_mt_axi_s_awaddr(i_dcd_dec_2_init_mt_axi_s_awaddr),
    .i_dcd_dec_2_init_mt_axi_s_awburst(i_dcd_dec_2_init_mt_axi_s_awburst),
    .i_dcd_dec_2_init_mt_axi_s_awcache(i_dcd_dec_2_init_mt_axi_s_awcache),
    .i_dcd_dec_2_init_mt_axi_s_awid(i_dcd_dec_2_init_mt_axi_s_awid),
    .i_dcd_dec_2_init_mt_axi_s_awlen(i_dcd_dec_2_init_mt_axi_s_awlen),
    .i_dcd_dec_2_init_mt_axi_s_awlock(i_dcd_dec_2_init_mt_axi_s_awlock),
    .i_dcd_dec_2_init_mt_axi_s_awprot(i_dcd_dec_2_init_mt_axi_s_awprot),
    .i_dcd_dec_2_init_mt_axi_s_awqos(i_dcd_dec_2_init_mt_axi_s_awqos),
    .o_dcd_dec_2_init_mt_axi_s_awready(o_dcd_dec_2_init_mt_axi_s_awready),
    .i_dcd_dec_2_init_mt_axi_s_awsize(i_dcd_dec_2_init_mt_axi_s_awsize),
    .i_dcd_dec_2_init_mt_axi_s_awvalid(i_dcd_dec_2_init_mt_axi_s_awvalid),
    .o_dcd_dec_2_init_mt_axi_s_bid(o_dcd_dec_2_init_mt_axi_s_bid),
    .i_dcd_dec_2_init_mt_axi_s_bready(i_dcd_dec_2_init_mt_axi_s_bready),
    .o_dcd_dec_2_init_mt_axi_s_bresp(o_dcd_dec_2_init_mt_axi_s_bresp),
    .o_dcd_dec_2_init_mt_axi_s_bvalid(o_dcd_dec_2_init_mt_axi_s_bvalid),
    .i_dcd_dec_2_init_mt_axi_s_wdata(i_dcd_dec_2_init_mt_axi_s_wdata),
    .i_dcd_dec_2_init_mt_axi_s_wlast(i_dcd_dec_2_init_mt_axi_s_wlast),
    .o_dcd_dec_2_init_mt_axi_s_wready(o_dcd_dec_2_init_mt_axi_s_wready),
    .i_dcd_dec_2_init_mt_axi_s_wstrb(i_dcd_dec_2_init_mt_axi_s_wstrb),
    .i_dcd_dec_2_init_mt_axi_s_wvalid(i_dcd_dec_2_init_mt_axi_s_wvalid),
    .i_dcd_mcu_clk(i_dcd_mcu_clk),
    .i_dcd_mcu_clken(i_dcd_mcu_clken),
    .i_dcd_mcu_init_lt_axi_s_araddr(i_dcd_mcu_init_lt_axi_s_araddr),
    .i_dcd_mcu_init_lt_axi_s_arburst(i_dcd_mcu_init_lt_axi_s_arburst),
    .i_dcd_mcu_init_lt_axi_s_arcache(i_dcd_mcu_init_lt_axi_s_arcache),
    .i_dcd_mcu_init_lt_axi_s_arid(i_dcd_mcu_init_lt_axi_s_arid),
    .i_dcd_mcu_init_lt_axi_s_arlen(i_dcd_mcu_init_lt_axi_s_arlen),
    .i_dcd_mcu_init_lt_axi_s_arlock(i_dcd_mcu_init_lt_axi_s_arlock),
    .i_dcd_mcu_init_lt_axi_s_arprot(i_dcd_mcu_init_lt_axi_s_arprot),
    .i_dcd_mcu_init_lt_axi_s_arqos(i_dcd_mcu_init_lt_axi_s_arqos),
    .o_dcd_mcu_init_lt_axi_s_arready(o_dcd_mcu_init_lt_axi_s_arready),
    .i_dcd_mcu_init_lt_axi_s_arsize(i_dcd_mcu_init_lt_axi_s_arsize),
    .i_dcd_mcu_init_lt_axi_s_arvalid(i_dcd_mcu_init_lt_axi_s_arvalid),
    .o_dcd_mcu_init_lt_axi_s_rdata(o_dcd_mcu_init_lt_axi_s_rdata),
    .o_dcd_mcu_init_lt_axi_s_rid(o_dcd_mcu_init_lt_axi_s_rid),
    .o_dcd_mcu_init_lt_axi_s_rlast(o_dcd_mcu_init_lt_axi_s_rlast),
    .i_dcd_mcu_init_lt_axi_s_rready(i_dcd_mcu_init_lt_axi_s_rready),
    .o_dcd_mcu_init_lt_axi_s_rresp(o_dcd_mcu_init_lt_axi_s_rresp),
    .o_dcd_mcu_init_lt_axi_s_rvalid(o_dcd_mcu_init_lt_axi_s_rvalid),
    .i_dcd_mcu_init_lt_axi_s_awaddr(i_dcd_mcu_init_lt_axi_s_awaddr),
    .i_dcd_mcu_init_lt_axi_s_awburst(i_dcd_mcu_init_lt_axi_s_awburst),
    .i_dcd_mcu_init_lt_axi_s_awcache(i_dcd_mcu_init_lt_axi_s_awcache),
    .i_dcd_mcu_init_lt_axi_s_awid(i_dcd_mcu_init_lt_axi_s_awid),
    .i_dcd_mcu_init_lt_axi_s_awlen(i_dcd_mcu_init_lt_axi_s_awlen),
    .i_dcd_mcu_init_lt_axi_s_awlock(i_dcd_mcu_init_lt_axi_s_awlock),
    .i_dcd_mcu_init_lt_axi_s_awprot(i_dcd_mcu_init_lt_axi_s_awprot),
    .i_dcd_mcu_init_lt_axi_s_awqos(i_dcd_mcu_init_lt_axi_s_awqos),
    .o_dcd_mcu_init_lt_axi_s_awready(o_dcd_mcu_init_lt_axi_s_awready),
    .i_dcd_mcu_init_lt_axi_s_awsize(i_dcd_mcu_init_lt_axi_s_awsize),
    .i_dcd_mcu_init_lt_axi_s_awvalid(i_dcd_mcu_init_lt_axi_s_awvalid),
    .o_dcd_mcu_init_lt_axi_s_bid(o_dcd_mcu_init_lt_axi_s_bid),
    .i_dcd_mcu_init_lt_axi_s_bready(i_dcd_mcu_init_lt_axi_s_bready),
    .o_dcd_mcu_init_lt_axi_s_bresp(o_dcd_mcu_init_lt_axi_s_bresp),
    .o_dcd_mcu_init_lt_axi_s_bvalid(o_dcd_mcu_init_lt_axi_s_bvalid),
    .i_dcd_mcu_init_lt_axi_s_wdata(i_dcd_mcu_init_lt_axi_s_wdata),
    .i_dcd_mcu_init_lt_axi_s_wlast(i_dcd_mcu_init_lt_axi_s_wlast),
    .o_dcd_mcu_init_lt_axi_s_wready(o_dcd_mcu_init_lt_axi_s_wready),
    .i_dcd_mcu_init_lt_axi_s_wstrb(i_dcd_mcu_init_lt_axi_s_wstrb),
    .i_dcd_mcu_init_lt_axi_s_wvalid(i_dcd_mcu_init_lt_axi_s_wvalid),
    .o_dcd_mcu_pwr_idle_val(o_dcd_mcu_pwr_idle_val),
    .o_dcd_mcu_pwr_idle_ack(o_dcd_mcu_pwr_idle_ack),
    .i_dcd_mcu_pwr_idle_req(i_dcd_mcu_pwr_idle_req),
    .i_dcd_mcu_rst_n(i_dcd_mcu_rst_n),
    .o_dcd_pwr_idle_val(o_dcd_pwr_idle_val),
    .o_dcd_pwr_idle_ack(o_dcd_pwr_idle_ack),
    .i_dcd_pwr_idle_req(i_dcd_pwr_idle_req),
    .o_dcd_targ_cfg_apb_m_paddr(o_dcd_targ_cfg_apb_m_paddr),
    .o_dcd_targ_cfg_apb_m_penable(o_dcd_targ_cfg_apb_m_penable),
    .o_dcd_targ_cfg_apb_m_pprot(o_dcd_targ_cfg_apb_m_pprot),
    .i_dcd_targ_cfg_apb_m_prdata(i_dcd_targ_cfg_apb_m_prdata),
    .i_dcd_targ_cfg_apb_m_pready(i_dcd_targ_cfg_apb_m_pready),
    .o_dcd_targ_cfg_apb_m_psel(o_dcd_targ_cfg_apb_m_psel),
    .i_dcd_targ_cfg_apb_m_pslverr(i_dcd_targ_cfg_apb_m_pslverr),
    .o_dcd_targ_cfg_apb_m_pstrb(o_dcd_targ_cfg_apb_m_pstrb),
    .o_dcd_targ_cfg_apb_m_pwdata(o_dcd_targ_cfg_apb_m_pwdata),
    .o_dcd_targ_cfg_apb_m_pwrite(o_dcd_targ_cfg_apb_m_pwrite),
    .o_dcd_targ_syscfg_apb_m_paddr(o_dcd_targ_syscfg_apb_m_paddr),
    .o_dcd_targ_syscfg_apb_m_penable(o_dcd_targ_syscfg_apb_m_penable),
    .o_dcd_targ_syscfg_apb_m_pprot(o_dcd_targ_syscfg_apb_m_pprot),
    .i_dcd_targ_syscfg_apb_m_prdata(i_dcd_targ_syscfg_apb_m_prdata),
    .i_dcd_targ_syscfg_apb_m_pready(i_dcd_targ_syscfg_apb_m_pready),
    .o_dcd_targ_syscfg_apb_m_psel(o_dcd_targ_syscfg_apb_m_psel),
    .i_dcd_targ_syscfg_apb_m_pslverr(i_dcd_targ_syscfg_apb_m_pslverr),
    .o_dcd_targ_syscfg_apb_m_pstrb(o_dcd_targ_syscfg_apb_m_pstrb),
    .o_dcd_targ_syscfg_apb_m_pwdata(o_dcd_targ_syscfg_apb_m_pwdata),
    .o_dcd_targ_syscfg_apb_m_pwrite(o_dcd_targ_syscfg_apb_m_pwrite),
    .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data),
    .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head),
    .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy),
    .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail),
    .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld),
    .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data),
    .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head),
    .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data),
    .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head),
    .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy),
    .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail),
    .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld),
    .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data),
    .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head),
    .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data),
    .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head),
    .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy),
    .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail),
    .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld),
    .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data),
    .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head),
    .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data),
    .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head),
    .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy),
    .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail),
    .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld),
    .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data),
    .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head),
    .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data),
    .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head),
    .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy),
    .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail),
    .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld),
    .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data),
    .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head),
    .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy),
    .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail),
    .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld),
    .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data),
    .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head),
    .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy),
    .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail),
    .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld),
    .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data),
    .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head),
    .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy),
    .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail),
    .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head),
    .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head),
    .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head),
    .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head),
    .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld),
    .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data),
    .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head),
    .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy),
    .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail),
    .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld),
    .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data),
    .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head),
    .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy),
    .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail),
    .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld),
    .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data),
    .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head),
    .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy),
    .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail),
    .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld),
    .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data),
    .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head),
    .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data),
    .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head),
    .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy),
    .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail),
    .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld),
    .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data),
    .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head),
    .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data),
    .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head),
    .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy),
    .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail),
    .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld),
    .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data),
    .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head),
    .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy),
    .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail),
    .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld),
    .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .lnk_buff_dec_128_to_256_ddr_e0_req_mainpde(impl_to_mem[0].pde),
    .lnk_buff_dec_128_to_256_ddr_e0_req_mainprn(impl_from_mem[0].prn),
    .lnk_buff_dec_128_to_256_ddr_e0_req_mainret(impl_to_mem[0].ret),
    .lnk_buff_dec_128_to_256_ddr_e0_req_mainse(impl_to_mem[0].se),
    .lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainpde(impl_to_mem[1].pde),
    .lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainprn(impl_from_mem[1].prn),
    .lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainret(impl_to_mem[1].ret),
    .lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainse(impl_to_mem[1].se),
    .lnk_buff_dec_128_to_256_ddr_e1_req_mainpde(impl_to_mem[2].pde),
    .lnk_buff_dec_128_to_256_ddr_e1_req_mainprn(impl_from_mem[2].prn),
    .lnk_buff_dec_128_to_256_ddr_e1_req_mainret(impl_to_mem[2].ret),
    .lnk_buff_dec_128_to_256_ddr_e1_req_mainse(impl_to_mem[2].se),
    .lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainpde(impl_to_mem[3].pde),
    .lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainprn(impl_from_mem[3].prn),
    .lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainret(impl_to_mem[3].ret),
    .lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainse(impl_to_mem[3].se),
    .lnk_buff_dec_128_to_256_ddr_e2_req_mainpde(impl_to_mem[4].pde),
    .lnk_buff_dec_128_to_256_ddr_e2_req_mainprn(impl_from_mem[4].prn),
    .lnk_buff_dec_128_to_256_ddr_e2_req_mainret(impl_to_mem[4].ret),
    .lnk_buff_dec_128_to_256_ddr_e2_req_mainse(impl_to_mem[4].se),
    .lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainpde(impl_to_mem[5].pde),
    .lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainprn(impl_from_mem[5].prn),
    .lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainret(impl_to_mem[5].ret),
    .lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainse(impl_to_mem[5].se),
    .lnk_buff_dec_128_to_256_ddr_e3_req_mainpde(impl_to_mem[6].pde),
    .lnk_buff_dec_128_to_256_ddr_e3_req_mainprn(impl_from_mem[6].prn),
    .lnk_buff_dec_128_to_256_ddr_e3_req_mainret(impl_to_mem[6].ret),
    .lnk_buff_dec_128_to_256_ddr_e3_req_mainse(impl_to_mem[6].se),
    .lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainpde(impl_to_mem[7].pde),
    .lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainprn(impl_from_mem[7].prn),
    .lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainret(impl_to_mem[7].ret),
    .lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainse(impl_to_mem[7].se),
    .lnk_buff_soc_128_to_256_lt_req_mainpde(impl_to_mem[8].pde),
    .lnk_buff_soc_128_to_256_lt_req_mainprn(impl_from_mem[8].prn),
    .lnk_buff_soc_128_to_256_lt_req_mainret(impl_to_mem[8].ret),
    .lnk_buff_soc_128_to_256_lt_req_mainse(impl_to_mem[8].se),
    .lnk_buff_soc_128_to_256_lt_req_resp_mainpde(impl_to_mem[9].pde),
    .lnk_buff_soc_128_to_256_lt_req_resp_mainprn(impl_from_mem[9].prn),
    .lnk_buff_soc_128_to_256_lt_req_resp_mainret(impl_to_mem[9].ret),
    .lnk_buff_soc_128_to_256_lt_req_resp_mainse(impl_to_mem[9].se),
    .lnk_buff_soc_128_to_256_rd_req_resp_mainpde(impl_to_mem[10].pde),
    .lnk_buff_soc_128_to_256_rd_req_resp_mainprn(impl_from_mem[10].prn),
    .lnk_buff_soc_128_to_256_rd_req_resp_mainret(impl_to_mem[10].ret),
    .lnk_buff_soc_128_to_256_rd_req_resp_mainse(impl_to_mem[10].se),
    .lnk_buff_soc_128_to_256_wr_req_mainpde(impl_to_mem[11].pde),
    .lnk_buff_soc_128_to_256_wr_req_mainprn(impl_from_mem[11].prn),
    .lnk_buff_soc_128_to_256_wr_req_mainret(impl_to_mem[11].ret),
    .lnk_buff_soc_128_to_256_wr_req_mainse(impl_to_mem[11].se),
    .lnk_buff_soc_128_to_64_req_mainpde(impl_to_mem[12].pde),
    .lnk_buff_soc_128_to_64_req_mainprn(impl_from_mem[12].prn),
    .lnk_buff_soc_128_to_64_req_mainret(impl_to_mem[12].ret),
    .lnk_buff_soc_128_to_64_req_mainse(impl_to_mem[12].se),
    .lnk_buff_soc_128_to_64_req_resp_mainpde(impl_to_mem[13].pde),
    .lnk_buff_soc_128_to_64_req_resp_mainprn(impl_from_mem[13].prn),
    .lnk_buff_soc_128_to_64_req_resp_mainret(impl_to_mem[13].ret),
    .lnk_buff_soc_128_to_64_req_resp_mainse(impl_to_mem[13].se),
    .lnk_buff_soc_256_to_128_rd_req_resp_mainpde(impl_to_mem[14].pde),
    .lnk_buff_soc_256_to_128_rd_req_resp_mainprn(impl_from_mem[14].prn),
    .lnk_buff_soc_256_to_128_rd_req_resp_mainret(impl_to_mem[14].ret),
    .lnk_buff_soc_256_to_128_rd_req_resp_mainse(impl_to_mem[14].se),
    .lnk_buff_soc_256_to_128_wr_req_mainpde(impl_to_mem[15].pde),
    .lnk_buff_soc_256_to_128_wr_req_mainprn(impl_from_mem[15].prn),
    .lnk_buff_soc_256_to_128_wr_req_mainret(impl_to_mem[15].ret),
    .lnk_buff_soc_256_to_128_wr_req_mainse(impl_to_mem[15].se),
    .lnk_buff_soc_256_to_512_rd_req_resp_mainpde(impl_to_mem[16].pde),
    .lnk_buff_soc_256_to_512_rd_req_resp_mainprn(impl_from_mem[16].prn),
    .lnk_buff_soc_256_to_512_rd_req_resp_mainret(impl_to_mem[16].ret),
    .lnk_buff_soc_256_to_512_rd_req_resp_mainse(impl_to_mem[16].se),
    .lnk_buff_soc_256_to_512_wr_req_mainpde(impl_to_mem[17].pde),
    .lnk_buff_soc_256_to_512_wr_req_mainprn(impl_from_mem[17].prn),
    .lnk_buff_soc_256_to_512_wr_req_mainret(impl_to_mem[17].ret),
    .lnk_buff_soc_256_to_512_wr_req_mainse(impl_to_mem[17].se),
    .lnk_buff_soc_512_to_256_ddr_e0_req_mainpde(impl_to_mem[18].pde),
    .lnk_buff_soc_512_to_256_ddr_e0_req_mainprn(impl_from_mem[18].prn),
    .lnk_buff_soc_512_to_256_ddr_e0_req_mainret(impl_to_mem[18].ret),
    .lnk_buff_soc_512_to_256_ddr_e0_req_mainse(impl_to_mem[18].se),
    .lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainpde(impl_to_mem[19].pde),
    .lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainprn(impl_from_mem[19].prn),
    .lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainret(impl_to_mem[19].ret),
    .lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainse(impl_to_mem[19].se),
    .lnk_buff_soc_512_to_256_ddr_e1_req_mainpde(impl_to_mem[20].pde),
    .lnk_buff_soc_512_to_256_ddr_e1_req_mainprn(impl_from_mem[20].prn),
    .lnk_buff_soc_512_to_256_ddr_e1_req_mainret(impl_to_mem[20].ret),
    .lnk_buff_soc_512_to_256_ddr_e1_req_mainse(impl_to_mem[20].se),
    .lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainpde(impl_to_mem[21].pde),
    .lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainprn(impl_from_mem[21].prn),
    .lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainret(impl_to_mem[21].ret),
    .lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainse(impl_to_mem[21].se),
    .lnk_buff_soc_512_to_256_ddr_e2_req_mainpde(impl_to_mem[22].pde),
    .lnk_buff_soc_512_to_256_ddr_e2_req_mainprn(impl_from_mem[22].prn),
    .lnk_buff_soc_512_to_256_ddr_e2_req_mainret(impl_to_mem[22].ret),
    .lnk_buff_soc_512_to_256_ddr_e2_req_mainse(impl_to_mem[22].se),
    .lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainpde(impl_to_mem[23].pde),
    .lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainprn(impl_from_mem[23].prn),
    .lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainret(impl_to_mem[23].ret),
    .lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainse(impl_to_mem[23].se),
    .lnk_buff_soc_512_to_256_ddr_e3_req_mainpde(impl_to_mem[24].pde),
    .lnk_buff_soc_512_to_256_ddr_e3_req_mainprn(impl_from_mem[24].prn),
    .lnk_buff_soc_512_to_256_ddr_e3_req_mainret(impl_to_mem[24].ret),
    .lnk_buff_soc_512_to_256_ddr_e3_req_mainse(impl_to_mem[24].se),
    .lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainpde(impl_to_mem[25].pde),
    .lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainprn(impl_from_mem[25].prn),
    .lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainret(impl_to_mem[25].ret),
    .lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainse(impl_to_mem[25].se),
    .lnk_buff_soc_512_to_256_rd_req_resp_mainpde(impl_to_mem[26].pde),
    .lnk_buff_soc_512_to_256_rd_req_resp_mainprn(impl_from_mem[26].prn),
    .lnk_buff_soc_512_to_256_rd_req_resp_mainret(impl_to_mem[26].ret),
    .lnk_buff_soc_512_to_256_rd_req_resp_mainse(impl_to_mem[26].se),
    .lnk_buff_soc_512_to_256_wr_req_mainpde(impl_to_mem[27].pde),
    .lnk_buff_soc_512_to_256_wr_req_mainprn(impl_from_mem[27].prn),
    .lnk_buff_soc_512_to_256_wr_req_mainret(impl_to_mem[27].ret),
    .lnk_buff_soc_512_to_256_wr_req_mainse(impl_to_mem[27].se),
    .lnk_buff_soc_64_to_128_lt_req_mainpde(impl_to_mem[28].pde),
    .lnk_buff_soc_64_to_128_lt_req_mainprn(impl_from_mem[28].prn),
    .lnk_buff_soc_64_to_128_lt_req_mainret(impl_to_mem[28].ret),
    .lnk_buff_soc_64_to_128_lt_req_mainse(impl_to_mem[28].se),
    .lnk_buff_soc_64_to_128_lt_req_resp_mainpde(impl_to_mem[29].pde),
    .lnk_buff_soc_64_to_128_lt_req_resp_mainprn(impl_from_mem[29].prn),
    .lnk_buff_soc_64_to_128_lt_req_resp_mainret(impl_to_mem[29].ret),
    .lnk_buff_soc_64_to_128_lt_req_resp_mainse(impl_to_mem[29].se),
    .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .i_noc_clk(i_noc_clk),
    .i_noc_rst_n(i_noc_rst_n),
    .i_pcie_aon_clk(i_pcie_aon_clk),
    .i_pcie_aon_rst_n(pcie_aon_rst_n_synced),
    .i_pcie_init_mt_clk(i_pcie_init_mt_clk),
    .i_pcie_init_mt_clken(i_pcie_init_mt_clken),
    .o_pcie_init_mt_pwr_idle_val(o_pcie_init_mt_pwr_idle_val),
    .o_pcie_init_mt_pwr_idle_ack(o_pcie_init_mt_pwr_idle_ack),
    .i_pcie_init_mt_pwr_idle_req(i_pcie_init_mt_pwr_idle_req),
    .i_pcie_init_mt_axi_s_araddr(i_pcie_init_mt_axi_s_araddr),
    .i_pcie_init_mt_axi_s_arburst(i_pcie_init_mt_axi_s_arburst),
    .i_pcie_init_mt_axi_s_arcache(i_pcie_init_mt_axi_s_arcache),
    .i_pcie_init_mt_axi_s_arid(i_pcie_init_mt_axi_s_arid),
    .i_pcie_init_mt_axi_s_arlen(i_pcie_init_mt_axi_s_arlen),
    .i_pcie_init_mt_axi_s_arlock(i_pcie_init_mt_axi_s_arlock),
    .i_pcie_init_mt_axi_s_arprot(i_pcie_init_mt_axi_s_arprot),
    .i_pcie_init_mt_axi_s_arqos(i_pcie_init_mt_axi_s_arqos),
    .o_pcie_init_mt_axi_s_arready(o_pcie_init_mt_axi_s_arready),
    .i_pcie_init_mt_axi_s_arsize(i_pcie_init_mt_axi_s_arsize),
    .i_pcie_init_mt_axi_s_arvalid(i_pcie_init_mt_axi_s_arvalid),
    .o_pcie_init_mt_axi_s_rdata(o_pcie_init_mt_axi_s_rdata),
    .o_pcie_init_mt_axi_s_rid(o_pcie_init_mt_axi_s_rid),
    .o_pcie_init_mt_axi_s_rlast(o_pcie_init_mt_axi_s_rlast),
    .i_pcie_init_mt_axi_s_rready(i_pcie_init_mt_axi_s_rready),
    .o_pcie_init_mt_axi_s_rresp(o_pcie_init_mt_axi_s_rresp),
    .o_pcie_init_mt_axi_s_rvalid(o_pcie_init_mt_axi_s_rvalid),
    .i_pcie_init_mt_rst_n(i_pcie_init_mt_rst_n),
    .i_pcie_init_mt_axi_s_awaddr(i_pcie_init_mt_axi_s_awaddr),
    .i_pcie_init_mt_axi_s_awburst(i_pcie_init_mt_axi_s_awburst),
    .i_pcie_init_mt_axi_s_awcache(i_pcie_init_mt_axi_s_awcache),
    .i_pcie_init_mt_axi_s_awid(i_pcie_init_mt_axi_s_awid),
    .i_pcie_init_mt_axi_s_awlen(i_pcie_init_mt_axi_s_awlen),
    .i_pcie_init_mt_axi_s_awlock(i_pcie_init_mt_axi_s_awlock),
    .i_pcie_init_mt_axi_s_awprot(i_pcie_init_mt_axi_s_awprot),
    .i_pcie_init_mt_axi_s_awqos(i_pcie_init_mt_axi_s_awqos),
    .o_pcie_init_mt_axi_s_awready(o_pcie_init_mt_axi_s_awready),
    .i_pcie_init_mt_axi_s_awsize(i_pcie_init_mt_axi_s_awsize),
    .i_pcie_init_mt_axi_s_awvalid(i_pcie_init_mt_axi_s_awvalid),
    .o_pcie_init_mt_axi_s_bid(o_pcie_init_mt_axi_s_bid),
    .i_pcie_init_mt_axi_s_bready(i_pcie_init_mt_axi_s_bready),
    .o_pcie_init_mt_axi_s_bresp(o_pcie_init_mt_axi_s_bresp),
    .o_pcie_init_mt_axi_s_bvalid(o_pcie_init_mt_axi_s_bvalid),
    .i_pcie_init_mt_axi_s_wdata(i_pcie_init_mt_axi_s_wdata),
    .i_pcie_init_mt_axi_s_wlast(i_pcie_init_mt_axi_s_wlast),
    .o_pcie_init_mt_axi_s_wready(o_pcie_init_mt_axi_s_wready),
    .i_pcie_init_mt_axi_s_wstrb(i_pcie_init_mt_axi_s_wstrb),
    .i_pcie_init_mt_axi_s_wvalid(i_pcie_init_mt_axi_s_wvalid),
    .o_pcie_targ_cfg_apb_m_paddr(o_pcie_targ_cfg_apb_m_paddr),
    .o_pcie_targ_cfg_apb_m_penable(o_pcie_targ_cfg_apb_m_penable),
    .o_pcie_targ_cfg_apb_m_pprot(o_pcie_targ_cfg_apb_m_pprot),
    .i_pcie_targ_cfg_apb_m_prdata(i_pcie_targ_cfg_apb_m_prdata),
    .i_pcie_targ_cfg_apb_m_pready(i_pcie_targ_cfg_apb_m_pready),
    .o_pcie_targ_cfg_apb_m_psel(o_pcie_targ_cfg_apb_m_psel),
    .i_pcie_targ_cfg_apb_m_pslverr(i_pcie_targ_cfg_apb_m_pslverr),
    .o_pcie_targ_cfg_apb_m_pstrb(o_pcie_targ_cfg_apb_m_pstrb),
    .o_pcie_targ_cfg_apb_m_pwdata(o_pcie_targ_cfg_apb_m_pwdata),
    .o_pcie_targ_cfg_apb_m_pwrite(o_pcie_targ_cfg_apb_m_pwrite),
    .i_pcie_targ_cfg_clk(i_pcie_targ_cfg_clk),
    .i_pcie_targ_cfg_clken(i_pcie_targ_cfg_clken),
    .o_pcie_targ_cfg_dbi_axi_m_araddr(o_pcie_targ_cfg_dbi_axi_m_araddr),
    .o_pcie_targ_cfg_dbi_axi_m_arburst(o_pcie_targ_cfg_dbi_axi_m_arburst),
    .o_pcie_targ_cfg_dbi_axi_m_arcache(o_pcie_targ_cfg_dbi_axi_m_arcache),
    .o_pcie_targ_cfg_dbi_axi_m_arid(o_pcie_targ_cfg_dbi_axi_m_arid),
    .o_pcie_targ_cfg_dbi_axi_m_arlen(o_pcie_targ_cfg_dbi_axi_m_arlen),
    .o_pcie_targ_cfg_dbi_axi_m_arlock(o_pcie_targ_cfg_dbi_axi_m_arlock),
    .o_pcie_targ_cfg_dbi_axi_m_arprot(o_pcie_targ_cfg_dbi_axi_m_arprot),
    .o_pcie_targ_cfg_dbi_axi_m_arqos(o_pcie_targ_cfg_dbi_axi_m_arqos),
    .i_pcie_targ_cfg_dbi_axi_m_arready(i_pcie_targ_cfg_dbi_axi_m_arready),
    .o_pcie_targ_cfg_dbi_axi_m_arsize(o_pcie_targ_cfg_dbi_axi_m_arsize),
    .o_pcie_targ_cfg_dbi_axi_m_arvalid(o_pcie_targ_cfg_dbi_axi_m_arvalid),
    .o_pcie_targ_cfg_dbi_axi_m_awaddr(o_pcie_targ_cfg_dbi_axi_m_awaddr),
    .o_pcie_targ_cfg_dbi_axi_m_awburst(o_pcie_targ_cfg_dbi_axi_m_awburst),
    .o_pcie_targ_cfg_dbi_axi_m_awcache(o_pcie_targ_cfg_dbi_axi_m_awcache),
    .o_pcie_targ_cfg_dbi_axi_m_awid(o_pcie_targ_cfg_dbi_axi_m_awid),
    .o_pcie_targ_cfg_dbi_axi_m_awlen(o_pcie_targ_cfg_dbi_axi_m_awlen),
    .o_pcie_targ_cfg_dbi_axi_m_awlock(o_pcie_targ_cfg_dbi_axi_m_awlock),
    .o_pcie_targ_cfg_dbi_axi_m_awprot(o_pcie_targ_cfg_dbi_axi_m_awprot),
    .o_pcie_targ_cfg_dbi_axi_m_awqos(o_pcie_targ_cfg_dbi_axi_m_awqos),
    .i_pcie_targ_cfg_dbi_axi_m_awready(i_pcie_targ_cfg_dbi_axi_m_awready),
    .o_pcie_targ_cfg_dbi_axi_m_awsize(o_pcie_targ_cfg_dbi_axi_m_awsize),
    .o_pcie_targ_cfg_dbi_axi_m_awvalid(o_pcie_targ_cfg_dbi_axi_m_awvalid),
    .i_pcie_targ_cfg_dbi_axi_m_bid(i_pcie_targ_cfg_dbi_axi_m_bid),
    .o_pcie_targ_cfg_dbi_axi_m_bready(o_pcie_targ_cfg_dbi_axi_m_bready),
    .i_pcie_targ_cfg_dbi_axi_m_bresp(i_pcie_targ_cfg_dbi_axi_m_bresp),
    .i_pcie_targ_cfg_dbi_axi_m_bvalid(i_pcie_targ_cfg_dbi_axi_m_bvalid),
    .i_pcie_targ_cfg_dbi_axi_m_rdata(i_pcie_targ_cfg_dbi_axi_m_rdata),
    .i_pcie_targ_cfg_dbi_axi_m_rid(i_pcie_targ_cfg_dbi_axi_m_rid),
    .i_pcie_targ_cfg_dbi_axi_m_rlast(i_pcie_targ_cfg_dbi_axi_m_rlast),
    .o_pcie_targ_cfg_dbi_axi_m_rready(o_pcie_targ_cfg_dbi_axi_m_rready),
    .i_pcie_targ_cfg_dbi_axi_m_rresp(i_pcie_targ_cfg_dbi_axi_m_rresp),
    .i_pcie_targ_cfg_dbi_axi_m_rvalid(i_pcie_targ_cfg_dbi_axi_m_rvalid),
    .o_pcie_targ_cfg_dbi_axi_m_wdata(o_pcie_targ_cfg_dbi_axi_m_wdata),
    .o_pcie_targ_cfg_dbi_axi_m_wlast(o_pcie_targ_cfg_dbi_axi_m_wlast),
    .i_pcie_targ_cfg_dbi_axi_m_wready(i_pcie_targ_cfg_dbi_axi_m_wready),
    .o_pcie_targ_cfg_dbi_axi_m_wstrb(o_pcie_targ_cfg_dbi_axi_m_wstrb),
    .o_pcie_targ_cfg_dbi_axi_m_wvalid(o_pcie_targ_cfg_dbi_axi_m_wvalid),
    .i_pcie_targ_cfg_dbi_clk(i_pcie_targ_cfg_dbi_clk),
    .i_pcie_targ_cfg_dbi_clken(i_pcie_targ_cfg_dbi_clken),
    .o_pcie_targ_cfg_dbi_pwr_idle_val(o_pcie_targ_cfg_dbi_pwr_idle_val),
    .o_pcie_targ_cfg_dbi_pwr_idle_ack(o_pcie_targ_cfg_dbi_pwr_idle_ack),
    .i_pcie_targ_cfg_dbi_pwr_idle_req(i_pcie_targ_cfg_dbi_pwr_idle_req),
    .i_pcie_targ_cfg_dbi_rst_n(i_pcie_targ_cfg_dbi_rst_n),
    .o_pcie_targ_cfg_pwr_idle_val(o_pcie_targ_cfg_pwr_idle_val),
    .o_pcie_targ_cfg_pwr_idle_ack(o_pcie_targ_cfg_pwr_idle_ack),
    .i_pcie_targ_cfg_pwr_idle_req(i_pcie_targ_cfg_pwr_idle_req),
    .i_pcie_targ_cfg_rst_n(i_pcie_targ_cfg_rst_n),
    .i_pcie_targ_mt_clk(i_pcie_targ_mt_clk),
    .i_pcie_targ_mt_clken(i_pcie_targ_mt_clken),
    .o_pcie_targ_mt_pwr_idle_val(o_pcie_targ_mt_pwr_idle_val),
    .o_pcie_targ_mt_pwr_idle_ack(o_pcie_targ_mt_pwr_idle_ack),
    .i_pcie_targ_mt_pwr_idle_req(i_pcie_targ_mt_pwr_idle_req),
    .o_pcie_targ_mt_axi_m_araddr(o_pcie_targ_mt_axi_m_araddr),
    .o_pcie_targ_mt_axi_m_arburst(o_pcie_targ_mt_axi_m_arburst),
    .o_pcie_targ_mt_axi_m_arcache(o_pcie_targ_mt_axi_m_arcache),
    .o_pcie_targ_mt_axi_m_arid(o_pcie_targ_mt_axi_m_arid),
    .o_pcie_targ_mt_axi_m_arlen(o_pcie_targ_mt_axi_m_arlen),
    .o_pcie_targ_mt_axi_m_arlock(o_pcie_targ_mt_axi_m_arlock),
    .o_pcie_targ_mt_axi_m_arprot(o_pcie_targ_mt_axi_m_arprot),
    .o_pcie_targ_mt_axi_m_arqos(o_pcie_targ_mt_axi_m_arqos),
    .i_pcie_targ_mt_axi_m_arready(i_pcie_targ_mt_axi_m_arready),
    .o_pcie_targ_mt_axi_m_arsize(o_pcie_targ_mt_axi_m_arsize),
    .o_pcie_targ_mt_axi_m_arvalid(o_pcie_targ_mt_axi_m_arvalid),
    .i_pcie_targ_mt_axi_m_rdata(i_pcie_targ_mt_axi_m_rdata),
    .i_pcie_targ_mt_axi_m_rid(i_pcie_targ_mt_axi_m_rid),
    .i_pcie_targ_mt_axi_m_rlast(i_pcie_targ_mt_axi_m_rlast),
    .o_pcie_targ_mt_axi_m_rready(o_pcie_targ_mt_axi_m_rready),
    .i_pcie_targ_mt_axi_m_rresp(i_pcie_targ_mt_axi_m_rresp),
    .i_pcie_targ_mt_axi_m_rvalid(i_pcie_targ_mt_axi_m_rvalid),
    .i_pcie_targ_mt_rst_n(i_pcie_targ_mt_rst_n),
    .o_pcie_targ_mt_axi_m_awaddr(o_pcie_targ_mt_axi_m_awaddr),
    .o_pcie_targ_mt_axi_m_awburst(o_pcie_targ_mt_axi_m_awburst),
    .o_pcie_targ_mt_axi_m_awcache(o_pcie_targ_mt_axi_m_awcache),
    .o_pcie_targ_mt_axi_m_awid(o_pcie_targ_mt_axi_m_awid),
    .o_pcie_targ_mt_axi_m_awlen(o_pcie_targ_mt_axi_m_awlen),
    .o_pcie_targ_mt_axi_m_awlock(o_pcie_targ_mt_axi_m_awlock),
    .o_pcie_targ_mt_axi_m_awprot(o_pcie_targ_mt_axi_m_awprot),
    .o_pcie_targ_mt_axi_m_awqos(o_pcie_targ_mt_axi_m_awqos),
    .i_pcie_targ_mt_axi_m_awready(i_pcie_targ_mt_axi_m_awready),
    .o_pcie_targ_mt_axi_m_awsize(o_pcie_targ_mt_axi_m_awsize),
    .o_pcie_targ_mt_axi_m_awvalid(o_pcie_targ_mt_axi_m_awvalid),
    .i_pcie_targ_mt_axi_m_bid(i_pcie_targ_mt_axi_m_bid),
    .o_pcie_targ_mt_axi_m_bready(o_pcie_targ_mt_axi_m_bready),
    .i_pcie_targ_mt_axi_m_bresp(i_pcie_targ_mt_axi_m_bresp),
    .i_pcie_targ_mt_axi_m_bvalid(i_pcie_targ_mt_axi_m_bvalid),
    .o_pcie_targ_mt_axi_m_wdata(o_pcie_targ_mt_axi_m_wdata),
    .o_pcie_targ_mt_axi_m_wlast(o_pcie_targ_mt_axi_m_wlast),
    .i_pcie_targ_mt_axi_m_wready(i_pcie_targ_mt_axi_m_wready),
    .o_pcie_targ_mt_axi_m_wstrb(o_pcie_targ_mt_axi_m_wstrb),
    .o_pcie_targ_mt_axi_m_wvalid(o_pcie_targ_mt_axi_m_wvalid),
    .o_pcie_targ_syscfg_apb_m_paddr(o_pcie_targ_syscfg_apb_m_paddr),
    .o_pcie_targ_syscfg_apb_m_penable(o_pcie_targ_syscfg_apb_m_penable),
    .o_pcie_targ_syscfg_apb_m_pprot(o_pcie_targ_syscfg_apb_m_pprot),
    .i_pcie_targ_syscfg_apb_m_prdata(i_pcie_targ_syscfg_apb_m_prdata),
    .i_pcie_targ_syscfg_apb_m_pready(i_pcie_targ_syscfg_apb_m_pready),
    .o_pcie_targ_syscfg_apb_m_psel(o_pcie_targ_syscfg_apb_m_psel),
    .i_pcie_targ_syscfg_apb_m_pslverr(i_pcie_targ_syscfg_apb_m_pslverr),
    .o_pcie_targ_syscfg_apb_m_pstrb(o_pcie_targ_syscfg_apb_m_pstrb),
    .o_pcie_targ_syscfg_apb_m_pwdata(o_pcie_targ_syscfg_apb_m_pwdata),
    .o_pcie_targ_syscfg_apb_m_pwrite(o_pcie_targ_syscfg_apb_m_pwrite),
    .i_pve_0_aon_clk(i_pve_0_aon_clk),
    .i_pve_0_aon_rst_n(pve_0_aon_rst_n_synced),
    .i_pve_0_clk(i_pve_0_clk),
    .i_pve_0_clken(i_pve_0_clken),
    .i_pve_0_init_ht_axi_s_araddr(i_pve_0_init_ht_axi_s_araddr),
    .i_pve_0_init_ht_axi_s_arburst(i_pve_0_init_ht_axi_s_arburst),
    .i_pve_0_init_ht_axi_s_arcache(i_pve_0_init_ht_axi_s_arcache),
    .i_pve_0_init_ht_axi_s_arid(i_pve_0_init_ht_axi_s_arid),
    .i_pve_0_init_ht_axi_s_arlen(i_pve_0_init_ht_axi_s_arlen),
    .i_pve_0_init_ht_axi_s_arlock(i_pve_0_init_ht_axi_s_arlock),
    .i_pve_0_init_ht_axi_s_arprot(i_pve_0_init_ht_axi_s_arprot),
    .o_pve_0_init_ht_axi_s_arready(o_pve_0_init_ht_axi_s_arready),
    .i_pve_0_init_ht_axi_s_arsize(i_pve_0_init_ht_axi_s_arsize),
    .i_pve_0_init_ht_axi_s_arvalid(i_pve_0_init_ht_axi_s_arvalid),
    .o_pve_0_init_ht_axi_s_rdata(o_pve_0_init_ht_axi_s_rdata),
    .o_pve_0_init_ht_axi_s_rid(o_pve_0_init_ht_axi_s_rid),
    .o_pve_0_init_ht_axi_s_rlast(o_pve_0_init_ht_axi_s_rlast),
    .i_pve_0_init_ht_axi_s_rready(i_pve_0_init_ht_axi_s_rready),
    .o_pve_0_init_ht_axi_s_rresp(o_pve_0_init_ht_axi_s_rresp),
    .o_pve_0_init_ht_axi_s_rvalid(o_pve_0_init_ht_axi_s_rvalid),
    .i_pve_0_init_ht_axi_s_awaddr(i_pve_0_init_ht_axi_s_awaddr),
    .i_pve_0_init_ht_axi_s_awburst(i_pve_0_init_ht_axi_s_awburst),
    .i_pve_0_init_ht_axi_s_awcache(i_pve_0_init_ht_axi_s_awcache),
    .i_pve_0_init_ht_axi_s_awid(i_pve_0_init_ht_axi_s_awid),
    .i_pve_0_init_ht_axi_s_awlen(i_pve_0_init_ht_axi_s_awlen),
    .i_pve_0_init_ht_axi_s_awlock(i_pve_0_init_ht_axi_s_awlock),
    .i_pve_0_init_ht_axi_s_awprot(i_pve_0_init_ht_axi_s_awprot),
    .o_pve_0_init_ht_axi_s_awready(o_pve_0_init_ht_axi_s_awready),
    .i_pve_0_init_ht_axi_s_awsize(i_pve_0_init_ht_axi_s_awsize),
    .i_pve_0_init_ht_axi_s_awvalid(i_pve_0_init_ht_axi_s_awvalid),
    .o_pve_0_init_ht_axi_s_bid(o_pve_0_init_ht_axi_s_bid),
    .i_pve_0_init_ht_axi_s_bready(i_pve_0_init_ht_axi_s_bready),
    .o_pve_0_init_ht_axi_s_bresp(o_pve_0_init_ht_axi_s_bresp),
    .o_pve_0_init_ht_axi_s_bvalid(o_pve_0_init_ht_axi_s_bvalid),
    .i_pve_0_init_ht_axi_s_wdata(i_pve_0_init_ht_axi_s_wdata),
    .i_pve_0_init_ht_axi_s_wlast(i_pve_0_init_ht_axi_s_wlast),
    .o_pve_0_init_ht_axi_s_wready(o_pve_0_init_ht_axi_s_wready),
    .i_pve_0_init_ht_axi_s_wstrb(i_pve_0_init_ht_axi_s_wstrb),
    .i_pve_0_init_ht_axi_s_wvalid(i_pve_0_init_ht_axi_s_wvalid),
    .i_pve_0_init_lt_axi_s_araddr(i_pve_0_init_lt_axi_s_araddr),
    .i_pve_0_init_lt_axi_s_arburst(i_pve_0_init_lt_axi_s_arburst),
    .i_pve_0_init_lt_axi_s_arcache(i_pve_0_init_lt_axi_s_arcache),
    .i_pve_0_init_lt_axi_s_arid(i_pve_0_init_lt_axi_s_arid),
    .i_pve_0_init_lt_axi_s_arlen(i_pve_0_init_lt_axi_s_arlen),
    .i_pve_0_init_lt_axi_s_arlock(i_pve_0_init_lt_axi_s_arlock),
    .i_pve_0_init_lt_axi_s_arprot(i_pve_0_init_lt_axi_s_arprot),
    .i_pve_0_init_lt_axi_s_arqos(i_pve_0_init_lt_axi_s_arqos),
    .o_pve_0_init_lt_axi_s_arready(o_pve_0_init_lt_axi_s_arready),
    .i_pve_0_init_lt_axi_s_arsize(i_pve_0_init_lt_axi_s_arsize),
    .i_pve_0_init_lt_axi_s_arvalid(i_pve_0_init_lt_axi_s_arvalid),
    .o_pve_0_init_lt_axi_s_rdata(o_pve_0_init_lt_axi_s_rdata),
    .o_pve_0_init_lt_axi_s_rid(o_pve_0_init_lt_axi_s_rid),
    .o_pve_0_init_lt_axi_s_rlast(o_pve_0_init_lt_axi_s_rlast),
    .i_pve_0_init_lt_axi_s_rready(i_pve_0_init_lt_axi_s_rready),
    .o_pve_0_init_lt_axi_s_rresp(o_pve_0_init_lt_axi_s_rresp),
    .o_pve_0_init_lt_axi_s_rvalid(o_pve_0_init_lt_axi_s_rvalid),
    .i_pve_0_init_lt_axi_s_awaddr(i_pve_0_init_lt_axi_s_awaddr),
    .i_pve_0_init_lt_axi_s_awburst(i_pve_0_init_lt_axi_s_awburst),
    .i_pve_0_init_lt_axi_s_awcache(i_pve_0_init_lt_axi_s_awcache),
    .i_pve_0_init_lt_axi_s_awid(i_pve_0_init_lt_axi_s_awid),
    .i_pve_0_init_lt_axi_s_awlen(i_pve_0_init_lt_axi_s_awlen),
    .i_pve_0_init_lt_axi_s_awlock(i_pve_0_init_lt_axi_s_awlock),
    .i_pve_0_init_lt_axi_s_awprot(i_pve_0_init_lt_axi_s_awprot),
    .i_pve_0_init_lt_axi_s_awqos(i_pve_0_init_lt_axi_s_awqos),
    .o_pve_0_init_lt_axi_s_awready(o_pve_0_init_lt_axi_s_awready),
    .i_pve_0_init_lt_axi_s_awsize(i_pve_0_init_lt_axi_s_awsize),
    .i_pve_0_init_lt_axi_s_awvalid(i_pve_0_init_lt_axi_s_awvalid),
    .o_pve_0_init_lt_axi_s_bid(o_pve_0_init_lt_axi_s_bid),
    .i_pve_0_init_lt_axi_s_bready(i_pve_0_init_lt_axi_s_bready),
    .o_pve_0_init_lt_axi_s_bresp(o_pve_0_init_lt_axi_s_bresp),
    .o_pve_0_init_lt_axi_s_bvalid(o_pve_0_init_lt_axi_s_bvalid),
    .i_pve_0_init_lt_axi_s_wdata(i_pve_0_init_lt_axi_s_wdata),
    .i_pve_0_init_lt_axi_s_wlast(i_pve_0_init_lt_axi_s_wlast),
    .o_pve_0_init_lt_axi_s_wready(o_pve_0_init_lt_axi_s_wready),
    .i_pve_0_init_lt_axi_s_wstrb(i_pve_0_init_lt_axi_s_wstrb),
    .i_pve_0_init_lt_axi_s_wvalid(i_pve_0_init_lt_axi_s_wvalid),
    .o_pve_0_pwr_idle_val(o_pve_0_pwr_idle_val),
    .o_pve_0_pwr_idle_ack(o_pve_0_pwr_idle_ack),
    .i_pve_0_pwr_idle_req(i_pve_0_pwr_idle_req),
    .i_pve_0_rst_n(i_pve_0_rst_n),
    .o_pve_0_targ_lt_axi_m_araddr(o_pve_0_targ_lt_axi_m_araddr),
    .o_pve_0_targ_lt_axi_m_arburst(o_pve_0_targ_lt_axi_m_arburst),
    .o_pve_0_targ_lt_axi_m_arcache(o_pve_0_targ_lt_axi_m_arcache),
    .o_pve_0_targ_lt_axi_m_arid(o_pve_0_targ_lt_axi_m_arid),
    .o_pve_0_targ_lt_axi_m_arlen(o_pve_0_targ_lt_axi_m_arlen),
    .o_pve_0_targ_lt_axi_m_arlock(o_pve_0_targ_lt_axi_m_arlock),
    .o_pve_0_targ_lt_axi_m_arprot(o_pve_0_targ_lt_axi_m_arprot),
    .o_pve_0_targ_lt_axi_m_arqos(o_pve_0_targ_lt_axi_m_arqos),
    .i_pve_0_targ_lt_axi_m_arready(i_pve_0_targ_lt_axi_m_arready),
    .o_pve_0_targ_lt_axi_m_arsize(o_pve_0_targ_lt_axi_m_arsize),
    .o_pve_0_targ_lt_axi_m_arvalid(o_pve_0_targ_lt_axi_m_arvalid),
    .o_pve_0_targ_lt_axi_m_awaddr(o_pve_0_targ_lt_axi_m_awaddr),
    .o_pve_0_targ_lt_axi_m_awburst(o_pve_0_targ_lt_axi_m_awburst),
    .o_pve_0_targ_lt_axi_m_awcache(o_pve_0_targ_lt_axi_m_awcache),
    .o_pve_0_targ_lt_axi_m_awid(o_pve_0_targ_lt_axi_m_awid),
    .o_pve_0_targ_lt_axi_m_awlen(o_pve_0_targ_lt_axi_m_awlen),
    .o_pve_0_targ_lt_axi_m_awlock(o_pve_0_targ_lt_axi_m_awlock),
    .o_pve_0_targ_lt_axi_m_awprot(o_pve_0_targ_lt_axi_m_awprot),
    .o_pve_0_targ_lt_axi_m_awqos(o_pve_0_targ_lt_axi_m_awqos),
    .i_pve_0_targ_lt_axi_m_awready(i_pve_0_targ_lt_axi_m_awready),
    .o_pve_0_targ_lt_axi_m_awsize(o_pve_0_targ_lt_axi_m_awsize),
    .o_pve_0_targ_lt_axi_m_awvalid(o_pve_0_targ_lt_axi_m_awvalid),
    .i_pve_0_targ_lt_axi_m_bid(i_pve_0_targ_lt_axi_m_bid),
    .o_pve_0_targ_lt_axi_m_bready(o_pve_0_targ_lt_axi_m_bready),
    .i_pve_0_targ_lt_axi_m_bresp(i_pve_0_targ_lt_axi_m_bresp),
    .i_pve_0_targ_lt_axi_m_bvalid(i_pve_0_targ_lt_axi_m_bvalid),
    .i_pve_0_targ_lt_axi_m_rdata(i_pve_0_targ_lt_axi_m_rdata),
    .i_pve_0_targ_lt_axi_m_rid(i_pve_0_targ_lt_axi_m_rid),
    .i_pve_0_targ_lt_axi_m_rlast(i_pve_0_targ_lt_axi_m_rlast),
    .o_pve_0_targ_lt_axi_m_rready(o_pve_0_targ_lt_axi_m_rready),
    .i_pve_0_targ_lt_axi_m_rresp(i_pve_0_targ_lt_axi_m_rresp),
    .i_pve_0_targ_lt_axi_m_rvalid(i_pve_0_targ_lt_axi_m_rvalid),
    .o_pve_0_targ_lt_axi_m_wdata(o_pve_0_targ_lt_axi_m_wdata),
    .o_pve_0_targ_lt_axi_m_wlast(o_pve_0_targ_lt_axi_m_wlast),
    .i_pve_0_targ_lt_axi_m_wready(i_pve_0_targ_lt_axi_m_wready),
    .o_pve_0_targ_lt_axi_m_wstrb(o_pve_0_targ_lt_axi_m_wstrb),
    .o_pve_0_targ_lt_axi_m_wvalid(o_pve_0_targ_lt_axi_m_wvalid),
    .o_pve_0_targ_syscfg_apb_m_paddr(o_pve_0_targ_syscfg_apb_m_paddr),
    .o_pve_0_targ_syscfg_apb_m_penable(o_pve_0_targ_syscfg_apb_m_penable),
    .o_pve_0_targ_syscfg_apb_m_pprot(o_pve_0_targ_syscfg_apb_m_pprot),
    .i_pve_0_targ_syscfg_apb_m_prdata(i_pve_0_targ_syscfg_apb_m_prdata),
    .i_pve_0_targ_syscfg_apb_m_pready(i_pve_0_targ_syscfg_apb_m_pready),
    .o_pve_0_targ_syscfg_apb_m_psel(o_pve_0_targ_syscfg_apb_m_psel),
    .i_pve_0_targ_syscfg_apb_m_pslverr(i_pve_0_targ_syscfg_apb_m_pslverr),
    .o_pve_0_targ_syscfg_apb_m_pstrb(o_pve_0_targ_syscfg_apb_m_pstrb),
    .o_pve_0_targ_syscfg_apb_m_pwdata(o_pve_0_targ_syscfg_apb_m_pwdata),
    .o_pve_0_targ_syscfg_apb_m_pwrite(o_pve_0_targ_syscfg_apb_m_pwrite),
    .i_pve_1_aon_clk(i_pve_1_aon_clk),
    .i_pve_1_aon_rst_n(pve_1_aon_rst_n_synced),
    .i_pve_1_clk(i_pve_1_clk),
    .i_pve_1_clken(i_pve_1_clken),
    .i_pve_1_init_ht_axi_s_araddr(i_pve_1_init_ht_axi_s_araddr),
    .i_pve_1_init_ht_axi_s_arburst(i_pve_1_init_ht_axi_s_arburst),
    .i_pve_1_init_ht_axi_s_arcache(i_pve_1_init_ht_axi_s_arcache),
    .i_pve_1_init_ht_axi_s_arid(i_pve_1_init_ht_axi_s_arid),
    .i_pve_1_init_ht_axi_s_arlen(i_pve_1_init_ht_axi_s_arlen),
    .i_pve_1_init_ht_axi_s_arlock(i_pve_1_init_ht_axi_s_arlock),
    .i_pve_1_init_ht_axi_s_arprot(i_pve_1_init_ht_axi_s_arprot),
    .o_pve_1_init_ht_axi_s_arready(o_pve_1_init_ht_axi_s_arready),
    .i_pve_1_init_ht_axi_s_arsize(i_pve_1_init_ht_axi_s_arsize),
    .i_pve_1_init_ht_axi_s_arvalid(i_pve_1_init_ht_axi_s_arvalid),
    .o_pve_1_init_ht_axi_s_rdata(o_pve_1_init_ht_axi_s_rdata),
    .o_pve_1_init_ht_axi_s_rid(o_pve_1_init_ht_axi_s_rid),
    .o_pve_1_init_ht_axi_s_rlast(o_pve_1_init_ht_axi_s_rlast),
    .i_pve_1_init_ht_axi_s_rready(i_pve_1_init_ht_axi_s_rready),
    .o_pve_1_init_ht_axi_s_rresp(o_pve_1_init_ht_axi_s_rresp),
    .o_pve_1_init_ht_axi_s_rvalid(o_pve_1_init_ht_axi_s_rvalid),
    .i_pve_1_init_ht_axi_s_awaddr(i_pve_1_init_ht_axi_s_awaddr),
    .i_pve_1_init_ht_axi_s_awburst(i_pve_1_init_ht_axi_s_awburst),
    .i_pve_1_init_ht_axi_s_awcache(i_pve_1_init_ht_axi_s_awcache),
    .i_pve_1_init_ht_axi_s_awid(i_pve_1_init_ht_axi_s_awid),
    .i_pve_1_init_ht_axi_s_awlen(i_pve_1_init_ht_axi_s_awlen),
    .i_pve_1_init_ht_axi_s_awlock(i_pve_1_init_ht_axi_s_awlock),
    .i_pve_1_init_ht_axi_s_awprot(i_pve_1_init_ht_axi_s_awprot),
    .o_pve_1_init_ht_axi_s_awready(o_pve_1_init_ht_axi_s_awready),
    .i_pve_1_init_ht_axi_s_awsize(i_pve_1_init_ht_axi_s_awsize),
    .i_pve_1_init_ht_axi_s_awvalid(i_pve_1_init_ht_axi_s_awvalid),
    .o_pve_1_init_ht_axi_s_bid(o_pve_1_init_ht_axi_s_bid),
    .i_pve_1_init_ht_axi_s_bready(i_pve_1_init_ht_axi_s_bready),
    .o_pve_1_init_ht_axi_s_bresp(o_pve_1_init_ht_axi_s_bresp),
    .o_pve_1_init_ht_axi_s_bvalid(o_pve_1_init_ht_axi_s_bvalid),
    .i_pve_1_init_ht_axi_s_wdata(i_pve_1_init_ht_axi_s_wdata),
    .i_pve_1_init_ht_axi_s_wlast(i_pve_1_init_ht_axi_s_wlast),
    .o_pve_1_init_ht_axi_s_wready(o_pve_1_init_ht_axi_s_wready),
    .i_pve_1_init_ht_axi_s_wstrb(i_pve_1_init_ht_axi_s_wstrb),
    .i_pve_1_init_ht_axi_s_wvalid(i_pve_1_init_ht_axi_s_wvalid),
    .i_pve_1_init_lt_axi_s_araddr(i_pve_1_init_lt_axi_s_araddr),
    .i_pve_1_init_lt_axi_s_arburst(i_pve_1_init_lt_axi_s_arburst),
    .i_pve_1_init_lt_axi_s_arcache(i_pve_1_init_lt_axi_s_arcache),
    .i_pve_1_init_lt_axi_s_arid(i_pve_1_init_lt_axi_s_arid),
    .i_pve_1_init_lt_axi_s_arlen(i_pve_1_init_lt_axi_s_arlen),
    .i_pve_1_init_lt_axi_s_arlock(i_pve_1_init_lt_axi_s_arlock),
    .i_pve_1_init_lt_axi_s_arprot(i_pve_1_init_lt_axi_s_arprot),
    .i_pve_1_init_lt_axi_s_arqos(i_pve_1_init_lt_axi_s_arqos),
    .o_pve_1_init_lt_axi_s_arready(o_pve_1_init_lt_axi_s_arready),
    .i_pve_1_init_lt_axi_s_arsize(i_pve_1_init_lt_axi_s_arsize),
    .i_pve_1_init_lt_axi_s_arvalid(i_pve_1_init_lt_axi_s_arvalid),
    .o_pve_1_init_lt_axi_s_rdata(o_pve_1_init_lt_axi_s_rdata),
    .o_pve_1_init_lt_axi_s_rid(o_pve_1_init_lt_axi_s_rid),
    .o_pve_1_init_lt_axi_s_rlast(o_pve_1_init_lt_axi_s_rlast),
    .i_pve_1_init_lt_axi_s_rready(i_pve_1_init_lt_axi_s_rready),
    .o_pve_1_init_lt_axi_s_rresp(o_pve_1_init_lt_axi_s_rresp),
    .o_pve_1_init_lt_axi_s_rvalid(o_pve_1_init_lt_axi_s_rvalid),
    .i_pve_1_init_lt_axi_s_awaddr(i_pve_1_init_lt_axi_s_awaddr),
    .i_pve_1_init_lt_axi_s_awburst(i_pve_1_init_lt_axi_s_awburst),
    .i_pve_1_init_lt_axi_s_awcache(i_pve_1_init_lt_axi_s_awcache),
    .i_pve_1_init_lt_axi_s_awid(i_pve_1_init_lt_axi_s_awid),
    .i_pve_1_init_lt_axi_s_awlen(i_pve_1_init_lt_axi_s_awlen),
    .i_pve_1_init_lt_axi_s_awlock(i_pve_1_init_lt_axi_s_awlock),
    .i_pve_1_init_lt_axi_s_awprot(i_pve_1_init_lt_axi_s_awprot),
    .i_pve_1_init_lt_axi_s_awqos(i_pve_1_init_lt_axi_s_awqos),
    .o_pve_1_init_lt_axi_s_awready(o_pve_1_init_lt_axi_s_awready),
    .i_pve_1_init_lt_axi_s_awsize(i_pve_1_init_lt_axi_s_awsize),
    .i_pve_1_init_lt_axi_s_awvalid(i_pve_1_init_lt_axi_s_awvalid),
    .o_pve_1_init_lt_axi_s_bid(o_pve_1_init_lt_axi_s_bid),
    .i_pve_1_init_lt_axi_s_bready(i_pve_1_init_lt_axi_s_bready),
    .o_pve_1_init_lt_axi_s_bresp(o_pve_1_init_lt_axi_s_bresp),
    .o_pve_1_init_lt_axi_s_bvalid(o_pve_1_init_lt_axi_s_bvalid),
    .i_pve_1_init_lt_axi_s_wdata(i_pve_1_init_lt_axi_s_wdata),
    .i_pve_1_init_lt_axi_s_wlast(i_pve_1_init_lt_axi_s_wlast),
    .o_pve_1_init_lt_axi_s_wready(o_pve_1_init_lt_axi_s_wready),
    .i_pve_1_init_lt_axi_s_wstrb(i_pve_1_init_lt_axi_s_wstrb),
    .i_pve_1_init_lt_axi_s_wvalid(i_pve_1_init_lt_axi_s_wvalid),
    .o_pve_1_pwr_idle_val(o_pve_1_pwr_idle_val),
    .o_pve_1_pwr_idle_ack(o_pve_1_pwr_idle_ack),
    .i_pve_1_pwr_idle_req(i_pve_1_pwr_idle_req),
    .i_pve_1_rst_n(i_pve_1_rst_n),
    .o_pve_1_targ_lt_axi_m_araddr(o_pve_1_targ_lt_axi_m_araddr),
    .o_pve_1_targ_lt_axi_m_arburst(o_pve_1_targ_lt_axi_m_arburst),
    .o_pve_1_targ_lt_axi_m_arcache(o_pve_1_targ_lt_axi_m_arcache),
    .o_pve_1_targ_lt_axi_m_arid(o_pve_1_targ_lt_axi_m_arid),
    .o_pve_1_targ_lt_axi_m_arlen(o_pve_1_targ_lt_axi_m_arlen),
    .o_pve_1_targ_lt_axi_m_arlock(o_pve_1_targ_lt_axi_m_arlock),
    .o_pve_1_targ_lt_axi_m_arprot(o_pve_1_targ_lt_axi_m_arprot),
    .o_pve_1_targ_lt_axi_m_arqos(o_pve_1_targ_lt_axi_m_arqos),
    .i_pve_1_targ_lt_axi_m_arready(i_pve_1_targ_lt_axi_m_arready),
    .o_pve_1_targ_lt_axi_m_arsize(o_pve_1_targ_lt_axi_m_arsize),
    .o_pve_1_targ_lt_axi_m_arvalid(o_pve_1_targ_lt_axi_m_arvalid),
    .o_pve_1_targ_lt_axi_m_awaddr(o_pve_1_targ_lt_axi_m_awaddr),
    .o_pve_1_targ_lt_axi_m_awburst(o_pve_1_targ_lt_axi_m_awburst),
    .o_pve_1_targ_lt_axi_m_awcache(o_pve_1_targ_lt_axi_m_awcache),
    .o_pve_1_targ_lt_axi_m_awid(o_pve_1_targ_lt_axi_m_awid),
    .o_pve_1_targ_lt_axi_m_awlen(o_pve_1_targ_lt_axi_m_awlen),
    .o_pve_1_targ_lt_axi_m_awlock(o_pve_1_targ_lt_axi_m_awlock),
    .o_pve_1_targ_lt_axi_m_awprot(o_pve_1_targ_lt_axi_m_awprot),
    .o_pve_1_targ_lt_axi_m_awqos(o_pve_1_targ_lt_axi_m_awqos),
    .i_pve_1_targ_lt_axi_m_awready(i_pve_1_targ_lt_axi_m_awready),
    .o_pve_1_targ_lt_axi_m_awsize(o_pve_1_targ_lt_axi_m_awsize),
    .o_pve_1_targ_lt_axi_m_awvalid(o_pve_1_targ_lt_axi_m_awvalid),
    .i_pve_1_targ_lt_axi_m_bid(i_pve_1_targ_lt_axi_m_bid),
    .o_pve_1_targ_lt_axi_m_bready(o_pve_1_targ_lt_axi_m_bready),
    .i_pve_1_targ_lt_axi_m_bresp(i_pve_1_targ_lt_axi_m_bresp),
    .i_pve_1_targ_lt_axi_m_bvalid(i_pve_1_targ_lt_axi_m_bvalid),
    .i_pve_1_targ_lt_axi_m_rdata(i_pve_1_targ_lt_axi_m_rdata),
    .i_pve_1_targ_lt_axi_m_rid(i_pve_1_targ_lt_axi_m_rid),
    .i_pve_1_targ_lt_axi_m_rlast(i_pve_1_targ_lt_axi_m_rlast),
    .o_pve_1_targ_lt_axi_m_rready(o_pve_1_targ_lt_axi_m_rready),
    .i_pve_1_targ_lt_axi_m_rresp(i_pve_1_targ_lt_axi_m_rresp),
    .i_pve_1_targ_lt_axi_m_rvalid(i_pve_1_targ_lt_axi_m_rvalid),
    .o_pve_1_targ_lt_axi_m_wdata(o_pve_1_targ_lt_axi_m_wdata),
    .o_pve_1_targ_lt_axi_m_wlast(o_pve_1_targ_lt_axi_m_wlast),
    .i_pve_1_targ_lt_axi_m_wready(i_pve_1_targ_lt_axi_m_wready),
    .o_pve_1_targ_lt_axi_m_wstrb(o_pve_1_targ_lt_axi_m_wstrb),
    .o_pve_1_targ_lt_axi_m_wvalid(o_pve_1_targ_lt_axi_m_wvalid),
    .o_pve_1_targ_syscfg_apb_m_paddr(o_pve_1_targ_syscfg_apb_m_paddr),
    .o_pve_1_targ_syscfg_apb_m_penable(o_pve_1_targ_syscfg_apb_m_penable),
    .o_pve_1_targ_syscfg_apb_m_pprot(o_pve_1_targ_syscfg_apb_m_pprot),
    .i_pve_1_targ_syscfg_apb_m_prdata(i_pve_1_targ_syscfg_apb_m_prdata),
    .i_pve_1_targ_syscfg_apb_m_pready(i_pve_1_targ_syscfg_apb_m_pready),
    .o_pve_1_targ_syscfg_apb_m_psel(o_pve_1_targ_syscfg_apb_m_psel),
    .i_pve_1_targ_syscfg_apb_m_pslverr(i_pve_1_targ_syscfg_apb_m_pslverr),
    .o_pve_1_targ_syscfg_apb_m_pstrb(o_pve_1_targ_syscfg_apb_m_pstrb),
    .o_pve_1_targ_syscfg_apb_m_pwdata(o_pve_1_targ_syscfg_apb_m_pwdata),
    .o_pve_1_targ_syscfg_apb_m_pwrite(o_pve_1_targ_syscfg_apb_m_pwrite),
    .scan_en(scan_en),
    .i_soc_mgmt_aon_clk(i_soc_mgmt_aon_clk),
    .i_soc_mgmt_aon_rst_n(soc_mgmt_aon_rst_n_synced),
    .i_soc_mgmt_clk(i_soc_mgmt_clk),
    .i_soc_mgmt_clken(i_soc_mgmt_clken),
    .i_soc_mgmt_init_lt_axi_s_araddr(i_soc_mgmt_init_lt_axi_s_araddr),
    .i_soc_mgmt_init_lt_axi_s_arburst(i_soc_mgmt_init_lt_axi_s_arburst),
    .i_soc_mgmt_init_lt_axi_s_arcache(i_soc_mgmt_init_lt_axi_s_arcache),
    .i_soc_mgmt_init_lt_axi_s_arid(i_soc_mgmt_init_lt_axi_s_arid),
    .i_soc_mgmt_init_lt_axi_s_arlen(i_soc_mgmt_init_lt_axi_s_arlen),
    .i_soc_mgmt_init_lt_axi_s_arlock(i_soc_mgmt_init_lt_axi_s_arlock),
    .i_soc_mgmt_init_lt_axi_s_arprot(i_soc_mgmt_init_lt_axi_s_arprot),
    .i_soc_mgmt_init_lt_axi_s_arqos(i_soc_mgmt_init_lt_axi_s_arqos),
    .o_soc_mgmt_init_lt_axi_s_arready(o_soc_mgmt_init_lt_axi_s_arready),
    .i_soc_mgmt_init_lt_axi_s_arsize(i_soc_mgmt_init_lt_axi_s_arsize),
    .i_soc_mgmt_init_lt_axi_s_arvalid(i_soc_mgmt_init_lt_axi_s_arvalid),
    .i_soc_mgmt_init_lt_axi_s_awaddr(i_soc_mgmt_init_lt_axi_s_awaddr),
    .i_soc_mgmt_init_lt_axi_s_awburst(i_soc_mgmt_init_lt_axi_s_awburst),
    .i_soc_mgmt_init_lt_axi_s_awcache(i_soc_mgmt_init_lt_axi_s_awcache),
    .i_soc_mgmt_init_lt_axi_s_awid(i_soc_mgmt_init_lt_axi_s_awid),
    .i_soc_mgmt_init_lt_axi_s_awlen(i_soc_mgmt_init_lt_axi_s_awlen),
    .i_soc_mgmt_init_lt_axi_s_awlock(i_soc_mgmt_init_lt_axi_s_awlock),
    .i_soc_mgmt_init_lt_axi_s_awprot(i_soc_mgmt_init_lt_axi_s_awprot),
    .i_soc_mgmt_init_lt_axi_s_awqos(i_soc_mgmt_init_lt_axi_s_awqos),
    .o_soc_mgmt_init_lt_axi_s_awready(o_soc_mgmt_init_lt_axi_s_awready),
    .i_soc_mgmt_init_lt_axi_s_awsize(i_soc_mgmt_init_lt_axi_s_awsize),
    .i_soc_mgmt_init_lt_axi_s_awvalid(i_soc_mgmt_init_lt_axi_s_awvalid),
    .o_soc_mgmt_init_lt_axi_s_bid(o_soc_mgmt_init_lt_axi_s_bid),
    .i_soc_mgmt_init_lt_axi_s_bready(i_soc_mgmt_init_lt_axi_s_bready),
    .o_soc_mgmt_init_lt_axi_s_bresp(o_soc_mgmt_init_lt_axi_s_bresp),
    .o_soc_mgmt_init_lt_axi_s_bvalid(o_soc_mgmt_init_lt_axi_s_bvalid),
    .o_soc_mgmt_init_lt_axi_s_rdata(o_soc_mgmt_init_lt_axi_s_rdata),
    .o_soc_mgmt_init_lt_axi_s_rid(o_soc_mgmt_init_lt_axi_s_rid),
    .o_soc_mgmt_init_lt_axi_s_rlast(o_soc_mgmt_init_lt_axi_s_rlast),
    .i_soc_mgmt_init_lt_axi_s_rready(i_soc_mgmt_init_lt_axi_s_rready),
    .o_soc_mgmt_init_lt_axi_s_rresp(o_soc_mgmt_init_lt_axi_s_rresp),
    .o_soc_mgmt_init_lt_axi_s_rvalid(o_soc_mgmt_init_lt_axi_s_rvalid),
    .i_soc_mgmt_init_lt_axi_s_wdata(i_soc_mgmt_init_lt_axi_s_wdata),
    .i_soc_mgmt_init_lt_axi_s_wlast(i_soc_mgmt_init_lt_axi_s_wlast),
    .o_soc_mgmt_init_lt_axi_s_wready(o_soc_mgmt_init_lt_axi_s_wready),
    .i_soc_mgmt_init_lt_axi_s_wstrb(i_soc_mgmt_init_lt_axi_s_wstrb),
    .i_soc_mgmt_init_lt_axi_s_wvalid(i_soc_mgmt_init_lt_axi_s_wvalid),
    .o_soc_mgmt_pwr_idle_val(o_soc_mgmt_pwr_idle_val),
    .o_soc_mgmt_pwr_idle_ack(o_soc_mgmt_pwr_idle_ack),
    .i_soc_mgmt_pwr_idle_req(i_soc_mgmt_pwr_idle_req),
    .i_soc_mgmt_rst_n(i_soc_mgmt_rst_n),
    .o_soc_mgmt_targ_lt_axi_m_araddr(o_soc_mgmt_targ_lt_axi_m_araddr),
    .o_soc_mgmt_targ_lt_axi_m_arburst(o_soc_mgmt_targ_lt_axi_m_arburst),
    .o_soc_mgmt_targ_lt_axi_m_arcache(o_soc_mgmt_targ_lt_axi_m_arcache),
    .o_soc_mgmt_targ_lt_axi_m_arid(o_soc_mgmt_targ_lt_axi_m_arid),
    .o_soc_mgmt_targ_lt_axi_m_arlen(o_soc_mgmt_targ_lt_axi_m_arlen),
    .o_soc_mgmt_targ_lt_axi_m_arlock(o_soc_mgmt_targ_lt_axi_m_arlock),
    .o_soc_mgmt_targ_lt_axi_m_arprot(o_soc_mgmt_targ_lt_axi_m_arprot),
    .o_soc_mgmt_targ_lt_axi_m_arqos(o_soc_mgmt_targ_lt_axi_m_arqos),
    .i_soc_mgmt_targ_lt_axi_m_arready(i_soc_mgmt_targ_lt_axi_m_arready),
    .o_soc_mgmt_targ_lt_axi_m_arsize(o_soc_mgmt_targ_lt_axi_m_arsize),
    .o_soc_mgmt_targ_lt_axi_m_arvalid(o_soc_mgmt_targ_lt_axi_m_arvalid),
    .o_soc_mgmt_targ_lt_axi_m_awaddr(o_soc_mgmt_targ_lt_axi_m_awaddr),
    .o_soc_mgmt_targ_lt_axi_m_awburst(o_soc_mgmt_targ_lt_axi_m_awburst),
    .o_soc_mgmt_targ_lt_axi_m_awcache(o_soc_mgmt_targ_lt_axi_m_awcache),
    .o_soc_mgmt_targ_lt_axi_m_awid(o_soc_mgmt_targ_lt_axi_m_awid),
    .o_soc_mgmt_targ_lt_axi_m_awlen(o_soc_mgmt_targ_lt_axi_m_awlen),
    .o_soc_mgmt_targ_lt_axi_m_awlock(o_soc_mgmt_targ_lt_axi_m_awlock),
    .o_soc_mgmt_targ_lt_axi_m_awprot(o_soc_mgmt_targ_lt_axi_m_awprot),
    .o_soc_mgmt_targ_lt_axi_m_awqos(o_soc_mgmt_targ_lt_axi_m_awqos),
    .i_soc_mgmt_targ_lt_axi_m_awready(i_soc_mgmt_targ_lt_axi_m_awready),
    .o_soc_mgmt_targ_lt_axi_m_awsize(o_soc_mgmt_targ_lt_axi_m_awsize),
    .o_soc_mgmt_targ_lt_axi_m_awvalid(o_soc_mgmt_targ_lt_axi_m_awvalid),
    .i_soc_mgmt_targ_lt_axi_m_bid(i_soc_mgmt_targ_lt_axi_m_bid),
    .o_soc_mgmt_targ_lt_axi_m_bready(o_soc_mgmt_targ_lt_axi_m_bready),
    .i_soc_mgmt_targ_lt_axi_m_bresp(i_soc_mgmt_targ_lt_axi_m_bresp),
    .i_soc_mgmt_targ_lt_axi_m_bvalid(i_soc_mgmt_targ_lt_axi_m_bvalid),
    .i_soc_mgmt_targ_lt_axi_m_rdata(i_soc_mgmt_targ_lt_axi_m_rdata),
    .i_soc_mgmt_targ_lt_axi_m_rid(i_soc_mgmt_targ_lt_axi_m_rid),
    .i_soc_mgmt_targ_lt_axi_m_rlast(i_soc_mgmt_targ_lt_axi_m_rlast),
    .o_soc_mgmt_targ_lt_axi_m_rready(o_soc_mgmt_targ_lt_axi_m_rready),
    .i_soc_mgmt_targ_lt_axi_m_rresp(i_soc_mgmt_targ_lt_axi_m_rresp),
    .i_soc_mgmt_targ_lt_axi_m_rvalid(i_soc_mgmt_targ_lt_axi_m_rvalid),
    .o_soc_mgmt_targ_lt_axi_m_wdata(o_soc_mgmt_targ_lt_axi_m_wdata),
    .o_soc_mgmt_targ_lt_axi_m_wlast(o_soc_mgmt_targ_lt_axi_m_wlast),
    .i_soc_mgmt_targ_lt_axi_m_wready(i_soc_mgmt_targ_lt_axi_m_wready),
    .o_soc_mgmt_targ_lt_axi_m_wstrb(o_soc_mgmt_targ_lt_axi_m_wstrb),
    .o_soc_mgmt_targ_lt_axi_m_wvalid(o_soc_mgmt_targ_lt_axi_m_wvalid),
    .o_soc_mgmt_targ_syscfg_apb_m_paddr(o_soc_mgmt_targ_syscfg_apb_m_paddr),
    .o_soc_mgmt_targ_syscfg_apb_m_penable(o_soc_mgmt_targ_syscfg_apb_m_penable),
    .o_soc_mgmt_targ_syscfg_apb_m_pprot(o_soc_mgmt_targ_syscfg_apb_m_pprot),
    .i_soc_mgmt_targ_syscfg_apb_m_prdata(i_soc_mgmt_targ_syscfg_apb_m_prdata),
    .i_soc_mgmt_targ_syscfg_apb_m_pready(i_soc_mgmt_targ_syscfg_apb_m_pready),
    .o_soc_mgmt_targ_syscfg_apb_m_psel(o_soc_mgmt_targ_syscfg_apb_m_psel),
    .i_soc_mgmt_targ_syscfg_apb_m_pslverr(i_soc_mgmt_targ_syscfg_apb_m_pslverr),
    .o_soc_mgmt_targ_syscfg_apb_m_pstrb(o_soc_mgmt_targ_syscfg_apb_m_pstrb),
    .o_soc_mgmt_targ_syscfg_apb_m_pwdata(o_soc_mgmt_targ_syscfg_apb_m_pwdata),
    .o_soc_mgmt_targ_syscfg_apb_m_pwrite(o_soc_mgmt_targ_syscfg_apb_m_pwrite),
    .i_sys_spm_aon_clk(i_sys_spm_aon_clk),
    .i_sys_spm_aon_rst_n(sys_spm_aon_rst_n_synced),
    .i_sys_spm_clk(i_sys_spm_clk),
    .i_sys_spm_clken(i_sys_spm_clken),
    .o_sys_spm_pwr_idle_val(o_sys_spm_pwr_idle_val),
    .o_sys_spm_pwr_idle_ack(o_sys_spm_pwr_idle_ack),
    .i_sys_spm_pwr_idle_req(i_sys_spm_pwr_idle_req),
    .i_sys_spm_rst_n(i_sys_spm_rst_n),
    .o_sys_spm_targ_lt_axi_m_araddr(o_sys_spm_targ_lt_axi_m_araddr),
    .o_sys_spm_targ_lt_axi_m_arburst(o_sys_spm_targ_lt_axi_m_arburst),
    .o_sys_spm_targ_lt_axi_m_arcache(o_sys_spm_targ_lt_axi_m_arcache),
    .o_sys_spm_targ_lt_axi_m_arid(o_sys_spm_targ_lt_axi_m_arid),
    .o_sys_spm_targ_lt_axi_m_arlen(o_sys_spm_targ_lt_axi_m_arlen),
    .o_sys_spm_targ_lt_axi_m_arlock(o_sys_spm_targ_lt_axi_m_arlock),
    .o_sys_spm_targ_lt_axi_m_arprot(o_sys_spm_targ_lt_axi_m_arprot),
    .o_sys_spm_targ_lt_axi_m_arqos(o_sys_spm_targ_lt_axi_m_arqos),
    .i_sys_spm_targ_lt_axi_m_arready(i_sys_spm_targ_lt_axi_m_arready),
    .o_sys_spm_targ_lt_axi_m_arsize(o_sys_spm_targ_lt_axi_m_arsize),
    .o_sys_spm_targ_lt_axi_m_arvalid(o_sys_spm_targ_lt_axi_m_arvalid),
    .o_sys_spm_targ_lt_axi_m_awaddr(o_sys_spm_targ_lt_axi_m_awaddr),
    .o_sys_spm_targ_lt_axi_m_awburst(o_sys_spm_targ_lt_axi_m_awburst),
    .o_sys_spm_targ_lt_axi_m_awcache(o_sys_spm_targ_lt_axi_m_awcache),
    .o_sys_spm_targ_lt_axi_m_awid(o_sys_spm_targ_lt_axi_m_awid),
    .o_sys_spm_targ_lt_axi_m_awlen(o_sys_spm_targ_lt_axi_m_awlen),
    .o_sys_spm_targ_lt_axi_m_awlock(o_sys_spm_targ_lt_axi_m_awlock),
    .o_sys_spm_targ_lt_axi_m_awprot(o_sys_spm_targ_lt_axi_m_awprot),
    .o_sys_spm_targ_lt_axi_m_awqos(o_sys_spm_targ_lt_axi_m_awqos),
    .i_sys_spm_targ_lt_axi_m_awready(i_sys_spm_targ_lt_axi_m_awready),
    .o_sys_spm_targ_lt_axi_m_awsize(o_sys_spm_targ_lt_axi_m_awsize),
    .o_sys_spm_targ_lt_axi_m_awvalid(o_sys_spm_targ_lt_axi_m_awvalid),
    .i_sys_spm_targ_lt_axi_m_bid(i_sys_spm_targ_lt_axi_m_bid),
    .o_sys_spm_targ_lt_axi_m_bready(o_sys_spm_targ_lt_axi_m_bready),
    .i_sys_spm_targ_lt_axi_m_bresp(i_sys_spm_targ_lt_axi_m_bresp),
    .i_sys_spm_targ_lt_axi_m_bvalid(i_sys_spm_targ_lt_axi_m_bvalid),
    .i_sys_spm_targ_lt_axi_m_rdata(i_sys_spm_targ_lt_axi_m_rdata),
    .i_sys_spm_targ_lt_axi_m_rid(i_sys_spm_targ_lt_axi_m_rid),
    .i_sys_spm_targ_lt_axi_m_rlast(i_sys_spm_targ_lt_axi_m_rlast),
    .o_sys_spm_targ_lt_axi_m_rready(o_sys_spm_targ_lt_axi_m_rready),
    .i_sys_spm_targ_lt_axi_m_rresp(i_sys_spm_targ_lt_axi_m_rresp),
    .i_sys_spm_targ_lt_axi_m_rvalid(i_sys_spm_targ_lt_axi_m_rvalid),
    .o_sys_spm_targ_lt_axi_m_wdata(o_sys_spm_targ_lt_axi_m_wdata),
    .o_sys_spm_targ_lt_axi_m_wlast(o_sys_spm_targ_lt_axi_m_wlast),
    .i_sys_spm_targ_lt_axi_m_wready(i_sys_spm_targ_lt_axi_m_wready),
    .o_sys_spm_targ_lt_axi_m_wstrb(o_sys_spm_targ_lt_axi_m_wstrb),
    .o_sys_spm_targ_lt_axi_m_wvalid(o_sys_spm_targ_lt_axi_m_wvalid),
    .o_sys_spm_targ_syscfg_apb_m_paddr(o_sys_spm_targ_syscfg_apb_m_paddr),
    .o_sys_spm_targ_syscfg_apb_m_penable(o_sys_spm_targ_syscfg_apb_m_penable),
    .o_sys_spm_targ_syscfg_apb_m_pprot(o_sys_spm_targ_syscfg_apb_m_pprot),
    .i_sys_spm_targ_syscfg_apb_m_prdata(i_sys_spm_targ_syscfg_apb_m_prdata),
    .i_sys_spm_targ_syscfg_apb_m_pready(i_sys_spm_targ_syscfg_apb_m_pready),
    .o_sys_spm_targ_syscfg_apb_m_psel(o_sys_spm_targ_syscfg_apb_m_psel),
    .i_sys_spm_targ_syscfg_apb_m_pslverr(i_sys_spm_targ_syscfg_apb_m_pslverr),
    .o_sys_spm_targ_syscfg_apb_m_pstrb(o_sys_spm_targ_syscfg_apb_m_pstrb),
    .o_sys_spm_targ_syscfg_apb_m_pwdata(o_sys_spm_targ_syscfg_apb_m_pwdata),
    .o_sys_spm_targ_syscfg_apb_m_pwrite(o_sys_spm_targ_syscfg_apb_m_pwrite)
);

noc_tok_soc u_noc_tok_soc (
  .i_apu_init_tok_ocpl_s_maddr(i_apu_init_tok_ocpl_s_maddr),
  .i_apu_init_tok_ocpl_s_mcmd({{ 2'b0, i_apu_init_tok_ocpl_s_mcmd }}),
  .i_apu_init_tok_ocpl_s_mdata(i_apu_init_tok_ocpl_s_mdata),
  .o_apu_init_tok_ocpl_s_scmdaccept(o_apu_init_tok_ocpl_s_scmdaccept),
  .o_apu_pwr_tok_idle_val(o_apu_pwr_tok_idle_val),
  .o_apu_pwr_tok_idle_ack(o_apu_pwr_tok_idle_ack),
  .i_apu_pwr_tok_idle_req(i_apu_pwr_tok_idle_req),
  .o_apu_targ_tok_ocpl_m_maddr(o_apu_targ_tok_ocpl_m_maddr),
  .o_apu_targ_tok_ocpl_m_mcmd(apu_targ_tok_ocpl_m_mcmd_ext),
  .o_apu_targ_tok_ocpl_m_mdata(o_apu_targ_tok_ocpl_m_mdata),
  .i_apu_targ_tok_ocpl_m_scmdaccept(i_apu_targ_tok_ocpl_m_scmdaccept),
  .i_apu_x_clk(i_apu_x_clk),
  .i_apu_x_clken(i_apu_x_clken),
  .i_apu_x_rst_n(i_apu_x_rst_n),
  .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data),
  .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head),
  .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy),
  .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail),
  .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld),
  .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data),
  .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head),
  .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy),
  .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail),
  .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld),
  .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data),
  .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head),
  .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy),
  .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail),
  .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld),
  .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data),
  .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head),
  .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy),
  .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail),
  .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld),
  .i_noc_clk(i_noc_clk),
  .i_noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en)
);
endmodule
