const phy_init_data_t snps_phy_init_details[string][] = '{
"A" : '{
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd196642},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd200738},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd16496},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd20592},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd45168},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd49264},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd1065072},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd1069168},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd1093744},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd1097840},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd2113648},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd2117744},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd2142320},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd2146416},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd3162224},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd3166320},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd3190896},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd3194992},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd5},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd4101},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd8197},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd12293},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd16389},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd20485},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd28677},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd32773},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd36869},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd40965},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd45061},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd49157},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd656136},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd655362},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd917574},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd917575},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd917576},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd917577},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd921670},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd921671},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd921672},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd921673},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd921674},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd917579},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd921675},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd925766},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd925767},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd925768},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd925769},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd929862},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd929863},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd929864},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd929865},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd929866},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd925771},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd929867},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd933958},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd933959},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd933960},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd933961},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd938054},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd938055},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd938056},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd938057},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd938058},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd933963},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd938059},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd942150},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd942151},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd942152},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd942153},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd946246},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd946247},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd946248},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd946249},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd946250},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd942155},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd946251},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd196640},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd200736},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd5},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd4101},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd8197},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd12293},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd16389},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd20485},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd28677},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd32773},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd36869},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd40965},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd45061},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd49157},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd656136},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd655362},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917574},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917575},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917576},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917577},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921670},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921671},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921672},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921673},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921674},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd917579},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd921675},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925766},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925767},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925768},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925769},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929862},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929863},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929864},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929865},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929866},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd925771},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd929867},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd933958},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd933959},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd933960},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd933961},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd938054},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd938055},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd938056},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd938057},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd938058},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd933963},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd938059},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942150},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942151},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942152},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942153},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946246},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946247},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946248},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946249},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946250},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd942155},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd946251},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd131237},
'{step_type : REG_WRITE,	value : 32'd2047,	reg_addr : 32'd65687},
'{step_type : REG_WRITE,	value : 32'd2047,	reg_addr : 32'd69783},
'{step_type : REG_WRITE,	value : 32'd2047,	reg_addr : 32'd73879},
'{step_type : REG_WRITE,	value : 32'd2047,	reg_addr : 32'd77975},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd65599},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65599},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd69695},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69695},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd73791},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73791},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd77887},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd77887},
'{step_type : REG_WRITE,	value : 32'd9,	reg_addr : 32'd721667},
'{step_type : REG_WRITE,	value : 32'd38,	reg_addr : 32'd656130},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd721665},
'{step_type : REG_WRITE,	value : 32'd29,	reg_addr : 32'd721679},
'{step_type : REG_WRITE,	value : 32'd6272,	reg_addr : 32'd196782},
'{step_type : REG_WRITE,	value : 32'd6272,	reg_addr : 32'd196781},
'{step_type : REG_WRITE,	value : 32'd6272,	reg_addr : 32'd196780},
'{step_type : REG_WRITE,	value : 32'd6272,	reg_addr : 32'd200878},
'{step_type : REG_WRITE,	value : 32'd6272,	reg_addr : 32'd200877},
'{step_type : REG_WRITE,	value : 32'd6272,	reg_addr : 32'd200876},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd786566},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459035},
'{step_type : REG_WRITE,	value : 32'd2099,	reg_addr : 32'd65699},
'{step_type : REG_WRITE,	value : 32'd2099,	reg_addr : 32'd69795},
'{step_type : REG_WRITE,	value : 32'd2099,	reg_addr : 32'd73891},
'{step_type : REG_WRITE,	value : 32'd2099,	reg_addr : 32'd77987},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd786672},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd786673},
'{step_type : REG_WRITE,	value : 32'd7,	reg_addr : 32'd786674},
'{step_type : REG_WRITE,	value : 32'd52,	reg_addr : 32'd786675},
'{step_type : REG_WRITE,	value : 32'd45,	reg_addr : 32'd591667},
'{step_type : REG_WRITE,	value : 32'd5,	reg_addr : 32'd786676},
'{step_type : REG_WRITE,	value : 32'd61440,	reg_addr : 32'd786679},
'{step_type : REG_WRITE,	value : 32'd2560,	reg_addr : 32'd591671},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd591647},
'{step_type : REG_WRITE,	value : 32'd15,	reg_addr : 32'd591913},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd131079},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917626},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd921722},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925818},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd929914},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd934010},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd938106},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942202},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd946298},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd1566},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd5662},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd9758},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd13854},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd17950},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd22046},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd30238},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd34334},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd38430},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd42526},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd46622},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd50718},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69151},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73247},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd77343},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd81439},
'{step_type : REG_WRITE,	value : 32'd61030,	reg_addr : 32'd198663},
'{step_type : REG_WRITE,	value : 32'd61030,	reg_addr : 32'd202759},
'{step_type : REG_WRITE,	value : 32'd61030,	reg_addr : 32'd67591},
'{step_type : REG_WRITE,	value : 32'd61030,	reg_addr : 32'd71687},
'{step_type : REG_WRITE,	value : 32'd61030,	reg_addr : 32'd75783},
'{step_type : REG_WRITE,	value : 32'd61030,	reg_addr : 32'd79879},
'{step_type : REG_WRITE,	value : 32'd16383,	reg_addr : 32'd196768},
'{step_type : REG_WRITE,	value : 32'd16383,	reg_addr : 32'd200864},
'{step_type : REG_WRITE,	value : 32'd8191,	reg_addr : 32'd65673},
'{step_type : REG_WRITE,	value : 32'd2047,	reg_addr : 32'd65674},
'{step_type : REG_WRITE,	value : 32'd8191,	reg_addr : 32'd69769},
'{step_type : REG_WRITE,	value : 32'd2047,	reg_addr : 32'd69770},
'{step_type : REG_WRITE,	value : 32'd8191,	reg_addr : 32'd73865},
'{step_type : REG_WRITE,	value : 32'd2047,	reg_addr : 32'd73866},
'{step_type : REG_WRITE,	value : 32'd8191,	reg_addr : 32'd77961},
'{step_type : REG_WRITE,	value : 32'd2047,	reg_addr : 32'd77962},
'{step_type : REG_WRITE,	value : 32'd15,	reg_addr : 32'd131078},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd131084},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd917517},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd921613},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd925709},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd929805},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd933901},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd937997},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd942093},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd946189},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd196647},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd63},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd4159},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd8255},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd12351},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd16447},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd20543},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd200743},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd28735},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd32831},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd36927},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd41023},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd45119},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd49215},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd131211},
'{step_type : REG_WRITE,	value : 32'd49314,	reg_addr : 32'd591873},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591874},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd591878},
'{step_type : REG_WRITE,	value : 32'd16641,	reg_addr : 32'd656383},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd656139},
'{step_type : REG_WRITE,	value : 32'd11930,	reg_addr : 32'd393224},
'{step_type : REG_WRITE,	value : 32'd100,	reg_addr : 32'd592096},
'{step_type : REG_WRITE,	value : 32'd300,	reg_addr : 32'd592097},
'{step_type : REG_WRITE,	value : 32'd2000,	reg_addr : 32'd592098},
'{step_type : REG_WRITE,	value : 32'd88,	reg_addr : 32'd592099},
'{step_type : REG_WRITE,	value : 32'd20,	reg_addr : 32'd592100},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd592101},
'{step_type : REG_WRITE,	value : 32'd67,	reg_addr : 32'd592102},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd592103},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd592106},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd592107},
'{step_type : REG_WRITE,	value : 32'd10,	reg_addr : 32'd592108},
'{step_type : REG_WRITE,	value : 32'd78,	reg_addr : 32'd592109},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd131074},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd393280},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd131072},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65787},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69883},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73979},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd78075},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917515},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921611},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925707},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929803},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd933899},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd937995},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942091},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946187},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd65572},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd69668},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd73764},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd77860},
'{step_type : REG_WRITE,	value : 32'd44,	reg_addr : 32'd65573},
'{step_type : REG_WRITE,	value : 32'd44,	reg_addr : 32'd69669},
'{step_type : REG_WRITE,	value : 32'd44,	reg_addr : 32'd73765},
'{step_type : REG_WRITE,	value : 32'd44,	reg_addr : 32'd77861},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65540},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65539},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69636},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69635},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73732},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73731},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd77828},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd77827},
'{step_type : REG_WRITE,	value : 32'd800,	reg_addr : 32'd720900},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd656140},
'{step_type : REG_WRITE,	value : 32'd5,	reg_addr : 32'd65598},
'{step_type : REG_WRITE,	value : 32'd5,	reg_addr : 32'd69694},
'{step_type : REG_WRITE,	value : 32'd5,	reg_addr : 32'd73790},
'{step_type : REG_WRITE,	value : 32'd5,	reg_addr : 32'd77886},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd131075},
'{step_type : REG_WRITE,	value : 32'd4369,	reg_addr : 32'd131083},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65800},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69896},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73992},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd78088},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd458757},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd458767},
'{step_type : REG_WRITE,	value : 32'd4864,	reg_addr : 32'd65550},
'{step_type : REG_WRITE,	value : 32'd4864,	reg_addr : 32'd69646},
'{step_type : REG_WRITE,	value : 32'd4864,	reg_addr : 32'd73742},
'{step_type : REG_WRITE,	value : 32'd4864,	reg_addr : 32'd77838},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd131097},
'{step_type : REG_WRITE,	value : 32'd51,	reg_addr : 32'd917548},
'{step_type : REG_WRITE,	value : 32'd51,	reg_addr : 32'd921644},
'{step_type : REG_WRITE,	value : 32'd771,	reg_addr : 32'd917549},
'{step_type : REG_WRITE,	value : 32'd13107,	reg_addr : 32'd921645},
'{step_type : REG_WRITE,	value : 32'd51,	reg_addr : 32'd925740},
'{step_type : REG_WRITE,	value : 32'd51,	reg_addr : 32'd929836},
'{step_type : REG_WRITE,	value : 32'd771,	reg_addr : 32'd925741},
'{step_type : REG_WRITE,	value : 32'd13107,	reg_addr : 32'd929837},
'{step_type : REG_WRITE,	value : 32'd51,	reg_addr : 32'd933932},
'{step_type : REG_WRITE,	value : 32'd51,	reg_addr : 32'd938028},
'{step_type : REG_WRITE,	value : 32'd771,	reg_addr : 32'd933933},
'{step_type : REG_WRITE,	value : 32'd13107,	reg_addr : 32'd938029},
'{step_type : REG_WRITE,	value : 32'd51,	reg_addr : 32'd942124},
'{step_type : REG_WRITE,	value : 32'd51,	reg_addr : 32'd946220},
'{step_type : REG_WRITE,	value : 32'd771,	reg_addr : 32'd942125},
'{step_type : REG_WRITE,	value : 32'd13107,	reg_addr : 32'd946221},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd112},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd4208},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd8304},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd12400},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd16496},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd20592},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd28784},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd32880},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd36976},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd41072},
'{step_type : REG_WRITE,	value : 32'd255,	reg_addr : 32'd45168},
'{step_type : REG_WRITE,	value : 32'd119,	reg_addr : 32'd49264},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd917550},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd921646},
'{step_type : REG_WRITE,	value : 32'd13056,	reg_addr : 32'd917551},
'{step_type : REG_WRITE,	value : 32'd30464,	reg_addr : 32'd921647},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd925742},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd929838},
'{step_type : REG_WRITE,	value : 32'd13056,	reg_addr : 32'd925743},
'{step_type : REG_WRITE,	value : 32'd30464,	reg_addr : 32'd929839},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd933934},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd938030},
'{step_type : REG_WRITE,	value : 32'd13056,	reg_addr : 32'd933935},
'{step_type : REG_WRITE,	value : 32'd30464,	reg_addr : 32'd938031},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd942126},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd946222},
'{step_type : REG_WRITE,	value : 32'd13056,	reg_addr : 32'd942127},
'{step_type : REG_WRITE,	value : 32'd30464,	reg_addr : 32'd946223},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd121},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd4217},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd8313},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd12409},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd16505},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd20601},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd28793},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd32889},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd36985},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd41081},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd45177},
'{step_type : REG_WRITE,	value : 32'd48,	reg_addr : 32'd49273},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd917532},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd921628},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd925724},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd929820},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd933916},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd938012},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd942108},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd946204},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd109},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd4205},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd8301},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd12397},
'{step_type : REG_WRITE,	value : 32'd248,	reg_addr : 32'd16493},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd20589},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd28781},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd32877},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd36973},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd41069},
'{step_type : REG_WRITE,	value : 32'd248,	reg_addr : 32'd45165},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd49261},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917566},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921662},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925758},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929854},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd933950},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd938046},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942142},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946238},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65537},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69633},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73729},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd77825},
'{step_type : REG_WRITE,	value : 32'd91,	reg_addr : 32'd458816},
'{step_type : REG_WRITE,	value : 32'd15,	reg_addr : 32'd458817},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd65701},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd69797},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd73893},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd77989},
'{step_type : REG_WRITE,	value : 32'd12850,	reg_addr : 32'd66057},
'{step_type : REG_WRITE,	value : 32'd12850,	reg_addr : 32'd70153},
'{step_type : REG_WRITE,	value : 32'd12850,	reg_addr : 32'd74249},
'{step_type : REG_WRITE,	value : 32'd12850,	reg_addr : 32'd78345},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd66063},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd70159},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd74255},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd78351},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd131077},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd65544},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd69640},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd73736},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd77832},
'{step_type : REG_WRITE,	value : 32'd546,	reg_addr : 32'd458859},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd458854},
'{step_type : REG_WRITE,	value : 32'd546,	reg_addr : 32'd458987},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd458982},
'{step_type : REG_WRITE,	value : 32'd4108,	reg_addr : 32'd459061},
'{step_type : REG_WRITE,	value : 32'd4108,	reg_addr : 32'd459062},
'{step_type : REG_WRITE,	value : 32'd1052,	reg_addr : 32'd459063},
'{step_type : REG_WRITE,	value : 32'd6944,	reg_addr : 32'd459064},
'{step_type : REG_WRITE,	value : 32'd4124,	reg_addr : 32'd459065},
'{step_type : REG_WRITE,	value : 32'd4124,	reg_addr : 32'd459066},
'{step_type : REG_WRITE,	value : 32'd1068,	reg_addr : 32'd459067},
'{step_type : REG_WRITE,	value : 32'd12080,	reg_addr : 32'd459068},
'{step_type : REG_WRITE,	value : 32'd4100,	reg_addr : 32'd459069},
'{step_type : REG_WRITE,	value : 32'd4100,	reg_addr : 32'd459070},
'{step_type : REG_WRITE,	value : 32'd1044,	reg_addr : 32'd459071},
'{step_type : REG_WRITE,	value : 32'd4888,	reg_addr : 32'd459072},
'{step_type : REG_WRITE,	value : 32'd2107,	reg_addr : 32'd459052},
'{step_type : REG_WRITE,	value : 32'd2107,	reg_addr : 32'd459053},
'{step_type : REG_WRITE,	value : 32'd2107,	reg_addr : 32'd459056},
'{step_type : REG_WRITE,	value : 32'd2079,	reg_addr : 32'd459054},
'{step_type : REG_WRITE,	value : 32'd2079,	reg_addr : 32'd459055},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd196616},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd200712},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917523},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921619},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925715},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929811},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd933907},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd938003},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942099},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946195},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd1507},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd5603},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd9699},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd13795},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd17891},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd21987},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd30179},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd34275},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd38371},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd42467},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd46563},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd50659},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd919011},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd923107},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd927203},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd931299},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd935395},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd939491},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd943587},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd947683},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd1290},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd5386},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd9482},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd13578},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd17674},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd21770},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd29962},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd34058},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd38154},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd42250},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd46346},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd50442},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd67595},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd71691},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd75787},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd79883},
'{step_type : REG_WRITE,	value : 32'd4202,	reg_addr : 32'd198659},
'{step_type : REG_WRITE,	value : 32'd4202,	reg_addr : 32'd202755},
'{step_type : REG_WRITE,	value : 32'd4202,	reg_addr : 32'd67587},
'{step_type : REG_WRITE,	value : 32'd4202,	reg_addr : 32'd71683},
'{step_type : REG_WRITE,	value : 32'd4202,	reg_addr : 32'd75779},
'{step_type : REG_WRITE,	value : 32'd4202,	reg_addr : 32'd79875},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd1283},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd5379},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd9475},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd13571},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd17667},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd21763},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd29955},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd34051},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd38147},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd42243},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd46339},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd50435},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd68611},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd72707},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd76803},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd80899},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd272},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd4368},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd8464},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd12560},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd16656},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd20752},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd28944},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd33040},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd37136},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd41232},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd45328},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd49424},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd917776},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd921872},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd925968},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd930064},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd934160},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd938256},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd942352},
'{step_type : REG_WRITE,	value : 32'd31,	reg_addr : 32'd946448},
'{step_type : REG_WRITE,	value : 32'd19,	reg_addr : 32'd592104},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd592105},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd917506},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd921602},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd925698},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd929794},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd933890},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd937986},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd942082},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd946178},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65803},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69899},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73995},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd78091},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd99},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd4195},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd8291},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd12387},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd16483},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd20579},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd28771},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd32867},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd36963},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd41059},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd45155},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd49251},
'{step_type : REG_WRITE,	value : 32'd616,	reg_addr : 32'd591882},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd591883},
'{step_type : REG_WRITE,	value : 32'd616,	reg_addr : 32'd591893},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd591894},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd917603},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd917604},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd917639},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd921699},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd921700},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd921735},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd925795},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd925796},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd925831},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd929891},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd929892},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd929927},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd933987},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd933988},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd934023},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd938083},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd938084},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd938119},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd942179},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd942180},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd942215},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd946275},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd946276},
'{step_type : REG_WRITE,	value : 32'd104,	reg_addr : 32'd946311},
'{step_type : REG_WRITE,	value : 32'd7,	reg_addr : 32'd786560},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd917564},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd921660},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd925756},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd929852},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd933948},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd938044},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd942140},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd946236},
'{step_type : REG_WRITE,	value : 32'd83,	reg_addr : 32'd591895},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591896},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591897},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd196843},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd200939},
'{step_type : REG_WRITE,	value : 32'd1008,	reg_addr : 32'd393222},
'{step_type : REG_WRITE,	value : 32'd156,	reg_addr : 32'd65753},
'{step_type : REG_WRITE,	value : 32'd156,	reg_addr : 32'd69849},
'{step_type : REG_WRITE,	value : 32'd156,	reg_addr : 32'd73945},
'{step_type : REG_WRITE,	value : 32'd156,	reg_addr : 32'd78041},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd65575},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd69671},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd73767},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd77863},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd196642},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd200738},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd196825},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd196824},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd197080},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd197336},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd197592},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd197848},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd198104},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd198360},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd198872},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd199128},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd200921},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd200920},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd201176},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd201432},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd201688},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd201944},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd202200},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd202456},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd202968},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd203224},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd65536},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd69632},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd73728},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd77824},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd458765},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd65578},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd65579},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd69674},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd69675},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd73770},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd73771},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd77866},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd77867},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd65576},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd65577},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd69672},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd69673},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd73768},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd73769},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd77864},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd77865},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd65658},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd65659},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd65914},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd65915},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd66170},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd66171},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd66426},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd66427},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd66682},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd66683},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd66938},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd66939},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd67194},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd67195},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd67450},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd67451},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd67706},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd67707},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd69754},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd69755},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd70010},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd70011},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd70266},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd70267},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd70522},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd70523},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd70778},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd70779},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd71034},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd71035},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd71290},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd71291},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd71546},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd71547},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd71802},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd71803},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd73850},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd73851},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd74106},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd74107},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd74362},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd74363},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd74618},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd74619},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd74874},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd74875},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd75130},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd75131},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd75386},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd75387},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd75642},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd75643},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd75898},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd75899},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd77946},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd77947},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd78202},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd78203},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd78458},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd78459},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd78714},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd78715},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd78970},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd78971},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd79226},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd79227},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd79482},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd79483},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd79738},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd79739},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd79994},
'{step_type : REG_WRITE,	value : 32'd237,	reg_addr : 32'd79995},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd65656},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd65657},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd65912},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd65913},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd66168},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd66169},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd66424},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd66425},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd66680},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd66681},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd66936},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd66937},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd67192},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd67193},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd67448},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd67449},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd67704},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd67705},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd69752},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd69753},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd70008},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd70009},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd70264},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd70265},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd70520},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd70521},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd70776},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd70777},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd71032},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd71033},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd71288},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd71289},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd71544},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd71545},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd71800},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd71801},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd73848},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd73849},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd74104},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd74105},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd74360},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd74361},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd74616},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd74617},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd74872},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd74873},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd75128},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd75129},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd75384},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd75385},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd75640},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd75641},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd75896},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd75897},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd77944},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd77945},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd78200},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd78201},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd78456},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd78457},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd78712},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd78713},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd78968},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd78969},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd79224},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd79225},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd79480},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd79481},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd79736},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd79737},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd79992},
'{step_type : REG_WRITE,	value : 32'd953,	reg_addr : 32'd79993},
'{step_type : REG_WRITE,	value : 32'd793,	reg_addr : 32'd65568},
'{step_type : REG_WRITE,	value : 32'd793,	reg_addr : 32'd65569},
'{step_type : REG_WRITE,	value : 32'd793,	reg_addr : 32'd69664},
'{step_type : REG_WRITE,	value : 32'd793,	reg_addr : 32'd69665},
'{step_type : REG_WRITE,	value : 32'd793,	reg_addr : 32'd73760},
'{step_type : REG_WRITE,	value : 32'd793,	reg_addr : 32'd73761},
'{step_type : REG_WRITE,	value : 32'd793,	reg_addr : 32'd77856},
'{step_type : REG_WRITE,	value : 32'd793,	reg_addr : 32'd77857},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd65552},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd65553},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd65554},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd65555},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd65808},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd65809},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd65810},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd65811},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66064},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66065},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66066},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66067},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66320},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66321},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66322},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66323},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66576},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66577},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66578},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66579},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66832},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66833},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66834},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd66835},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67088},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67089},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67090},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67091},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67344},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67345},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67346},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67347},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67600},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67601},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67602},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd67603},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd69648},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd69649},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd69650},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd69651},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd69904},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd69905},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd69906},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd69907},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70160},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70161},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70162},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70163},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70416},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70417},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70418},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70419},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70672},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70673},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70674},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70675},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70928},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70929},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70930},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd70931},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71184},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71185},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71186},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71187},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71440},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71441},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71442},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71443},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71696},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71697},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71698},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd71699},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd73744},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd73745},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd73746},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd73747},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74000},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74001},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74002},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74003},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74256},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74257},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74258},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74259},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74512},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74513},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74514},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74515},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74768},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74769},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74770},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd74771},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75024},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75025},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75026},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75027},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75280},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75281},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75282},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75283},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75536},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75537},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75538},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75539},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75792},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75793},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75794},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd75795},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd77840},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd77841},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd77842},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd77843},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78096},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78097},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78098},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78099},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78352},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78353},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78354},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78355},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78608},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78609},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78610},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78611},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78864},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78865},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78866},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd78867},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79120},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79121},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79122},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79123},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79376},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79377},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79378},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79379},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79632},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79633},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79634},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79635},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79888},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79889},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79890},
'{step_type : REG_WRITE,	value : 32'd299,	reg_addr : 32'd79891},
'{step_type : REG_WRITE,	value : 32'd204,	reg_addr : 32'd65548},
'{step_type : REG_WRITE,	value : 32'd204,	reg_addr : 32'd65549},
'{step_type : REG_WRITE,	value : 32'd408,	reg_addr : 32'd65556},
'{step_type : REG_WRITE,	value : 32'd408,	reg_addr : 32'd65557},
'{step_type : REG_WRITE,	value : 32'd204,	reg_addr : 32'd69644},
'{step_type : REG_WRITE,	value : 32'd204,	reg_addr : 32'd69645},
'{step_type : REG_WRITE,	value : 32'd408,	reg_addr : 32'd69652},
'{step_type : REG_WRITE,	value : 32'd408,	reg_addr : 32'd69653},
'{step_type : REG_WRITE,	value : 32'd204,	reg_addr : 32'd73740},
'{step_type : REG_WRITE,	value : 32'd204,	reg_addr : 32'd73741},
'{step_type : REG_WRITE,	value : 32'd408,	reg_addr : 32'd73748},
'{step_type : REG_WRITE,	value : 32'd408,	reg_addr : 32'd73749},
'{step_type : REG_WRITE,	value : 32'd204,	reg_addr : 32'd77836},
'{step_type : REG_WRITE,	value : 32'd204,	reg_addr : 32'd77837},
'{step_type : REG_WRITE,	value : 32'd408,	reg_addr : 32'd77844},
'{step_type : REG_WRITE,	value : 32'd408,	reg_addr : 32'd77845},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd458871},
'{step_type : REG_WRITE,	value : 32'd102,	reg_addr : 32'd131185},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd99},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd4195},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd8291},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd12387},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd16483},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd20579},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd28771},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd32867},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd36963},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd41059},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd45155},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd49251},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd917603},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd917604},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd917639},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd921699},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd921700},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd921735},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd925795},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd925796},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd925831},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd929891},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd929892},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd929927},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd933987},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd933988},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd934023},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd938083},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd938084},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd938119},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd942179},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd942180},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd942215},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd946275},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd946276},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd946311},
'{step_type : REG_WRITE,	value : 32'd610,	reg_addr : 32'd591882},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd591883},
'{step_type : REG_WRITE,	value : 32'd610,	reg_addr : 32'd591893},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd591894},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd65887},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd69983},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd74079},
'{step_type : REG_WRITE,	value : 32'd98,	reg_addr : 32'd78175},
'{step_type : REG_WRITE,	value : 32'd16,	reg_addr : 32'd393225},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd66208},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd66209},
'{step_type : REG_WRITE,	value : 32'd10,	reg_addr : 32'd66210},
'{step_type : REG_WRITE,	value : 32'd62,	reg_addr : 32'd66211},
'{step_type : REG_WRITE,	value : 32'd114,	reg_addr : 32'd66212},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd70304},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd70305},
'{step_type : REG_WRITE,	value : 32'd10,	reg_addr : 32'd70306},
'{step_type : REG_WRITE,	value : 32'd62,	reg_addr : 32'd70307},
'{step_type : REG_WRITE,	value : 32'd114,	reg_addr : 32'd70308},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd74400},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd74401},
'{step_type : REG_WRITE,	value : 32'd10,	reg_addr : 32'd74402},
'{step_type : REG_WRITE,	value : 32'd62,	reg_addr : 32'd74403},
'{step_type : REG_WRITE,	value : 32'd114,	reg_addr : 32'd74404},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd78496},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd78497},
'{step_type : REG_WRITE,	value : 32'd10,	reg_addr : 32'd78498},
'{step_type : REG_WRITE,	value : 32'd62,	reg_addr : 32'd78499},
'{step_type : REG_WRITE,	value : 32'd114,	reg_addr : 32'd78500},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd66221},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd70317},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd74413},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd78509},
'{step_type : REG_WRITE,	value : 32'd76,	reg_addr : 32'd66223},
'{step_type : REG_WRITE,	value : 32'd76,	reg_addr : 32'd70319},
'{step_type : REG_WRITE,	value : 32'd76,	reg_addr : 32'd74415},
'{step_type : REG_WRITE,	value : 32'd76,	reg_addr : 32'd78511},
'{step_type : REG_WRITE,	value : 32'd38657,	reg_addr : 32'd591879},
'{step_type : REG_WRITE,	value : 32'd46721,	reg_addr : 32'd591880},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd65599},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65599},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd69695},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69695},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd73791},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73791},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd77887},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd77887},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd721680},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd721681},
'{step_type : REG_WRITE,	value : 32'd11606,	reg_addr : 32'd393224},
'{step_type : REG_WRITE,	value : 32'd1008,	reg_addr : 32'd393222},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd196629},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd200725},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65660},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69756},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73852},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd77948},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd459073},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd720897},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591884},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd65575},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd69671},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd73767},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd77863},
'{step_type : REG_WRITE,	value : 32'd8,	reg_addr : 32'd66063},
'{step_type : REG_WRITE,	value : 32'd8,	reg_addr : 32'd70159},
'{step_type : REG_WRITE,	value : 32'd8,	reg_addr : 32'd74255},
'{step_type : REG_WRITE,	value : 32'd8,	reg_addr : 32'd78351},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd917567},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd917645},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd921663},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd921741},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd925759},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd925837},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd929855},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd929933},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd933951},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd934029},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd938047},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd938125},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd942143},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd942221},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd946239},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd946317},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd592131},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd458866},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd591886},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd458867},
'{step_type : REG_WRITE,	value : 32'd3,	reg_addr : 32'd591887},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd851968},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266240},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266241},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266242},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266243},
'{step_type : REG_WRITE,	value : 32'd49192,	reg_addr : 32'd267348},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267349},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267350},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267351},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267352},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267353},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267354},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267355},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267356},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267357},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267358},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267359},
'{step_type : REG_WRITE,	value : 32'd51288,	reg_addr : 32'd267360},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267361},
'{step_type : REG_WRITE,	value : 32'd57480,	reg_addr : 32'd267362},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267363},
'{step_type : REG_WRITE,	value : 32'd57400,	reg_addr : 32'd267364},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267365},
'{step_type : REG_WRITE,	value : 32'd51288,	reg_addr : 32'd267366},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267367},
'{step_type : REG_WRITE,	value : 32'd49288,	reg_addr : 32'd267368},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267369},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267370},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267371},
'{step_type : REG_WRITE,	value : 32'd49192,	reg_addr : 32'd267372},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267373},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267374},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267375},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267376},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267377},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267378},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267379},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267380},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267381},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267382},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267383},
'{step_type : REG_WRITE,	value : 32'd51288,	reg_addr : 32'd267384},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267385},
'{step_type : REG_WRITE,	value : 32'd57864,	reg_addr : 32'd267386},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267387},
'{step_type : REG_WRITE,	value : 32'd57400,	reg_addr : 32'd267388},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267389},
'{step_type : REG_WRITE,	value : 32'd51288,	reg_addr : 32'd267390},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267391},
'{step_type : REG_WRITE,	value : 32'd49672,	reg_addr : 32'd267392},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267393},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267394},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267395},
'{step_type : REG_WRITE,	value : 32'd49216,	reg_addr : 32'd267396},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267397},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267398},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267399},
'{step_type : REG_WRITE,	value : 32'd49256,	reg_addr : 32'd267400},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267401},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267402},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267403},
'{step_type : REG_WRITE,	value : 32'd52824,	reg_addr : 32'd267404},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267405},
'{step_type : REG_WRITE,	value : 32'd49672,	reg_addr : 32'd267406},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267407},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267408},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267409},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267410},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267411},
'{step_type : REG_WRITE,	value : 32'd17264,	reg_addr : 32'd267412},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267413},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267414},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267415},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267416},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267417},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267418},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267419},
'{step_type : REG_WRITE,	value : 32'd33648,	reg_addr : 32'd267420},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267421},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267422},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267423},
'{step_type : REG_WRITE,	value : 32'd53976,	reg_addr : 32'd267424},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267425},
'{step_type : REG_WRITE,	value : 32'd57352,	reg_addr : 32'd267426},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267427},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267428},
'{step_type : REG_WRITE,	value : 32'd2063597568,	reg_addr : 32'd267429},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267430},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267431},
'{step_type : REG_WRITE,	value : 32'd49392,	reg_addr : 32'd267432},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267433},
'{step_type : REG_WRITE,	value : 32'd53208,	reg_addr : 32'd267434},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267435},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267436},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267437},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267438},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267439},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267440},
'{step_type : REG_WRITE,	value : 32'd989855744,	reg_addr : 32'd267441},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267442},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267443},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267444},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267445},
'{step_type : REG_WRITE,	value : 32'd53336,	reg_addr : 32'd267446},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267447},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267448},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267449},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267450},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267451},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267452},
'{step_type : REG_WRITE,	value : 32'd989855744,	reg_addr : 32'd267453},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267454},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267455},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267456},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267457},
'{step_type : REG_WRITE,	value : 32'd53464,	reg_addr : 32'd267458},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267459},
'{step_type : REG_WRITE,	value : 32'd49288,	reg_addr : 32'd267460},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267461},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267462},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267463},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267464},
'{step_type : REG_WRITE,	value : 32'd989855744,	reg_addr : 32'd267465},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267466},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267467},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267468},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267469},
'{step_type : REG_WRITE,	value : 32'd53592,	reg_addr : 32'd267470},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267471},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267472},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267473},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267474},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267475},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267476},
'{step_type : REG_WRITE,	value : 32'd1795162112,	reg_addr : 32'd267477},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267478},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267479},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267480},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267481},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267482},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267483},
'{step_type : REG_WRITE,	value : 32'd218120236,	reg_addr : 32'd267484},
'{step_type : REG_WRITE,	value : 32'd67108865,	reg_addr : 32'd267485},
'{step_type : REG_WRITE,	value : 32'd134234192,	reg_addr : 32'd267486},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267487},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267488},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267489},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267490},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267491},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267492},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267493},
'{step_type : REG_WRITE,	value : 32'd134430800,	reg_addr : 32'd267494},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267495},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267496},
'{step_type : REG_WRITE,	value : 32'd520093696,	reg_addr : 32'd267497},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267498},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267499},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267500},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267501},
'{step_type : REG_WRITE,	value : 32'd16508,	reg_addr : 32'd267502},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267503},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267504},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267505},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267506},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267507},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267508},
'{step_type : REG_WRITE,	value : 32'd67108865,	reg_addr : 32'd267509},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267510},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267511},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267512},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267513},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267514},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267515},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267516},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267517},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267518},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267519},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267520},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267521},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267522},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267523},
'{step_type : REG_WRITE,	value : 32'd218136620,	reg_addr : 32'd267524},
'{step_type : REG_WRITE,	value : 32'd68157441,	reg_addr : 32'd267525},
'{step_type : REG_WRITE,	value : 32'd134250576,	reg_addr : 32'd267526},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267527},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267528},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267529},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267530},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267531},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267532},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267533},
'{step_type : REG_WRITE,	value : 32'd134447184,	reg_addr : 32'd267534},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267535},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267536},
'{step_type : REG_WRITE,	value : 32'd520093696,	reg_addr : 32'd267537},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267538},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267539},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267540},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267541},
'{step_type : REG_WRITE,	value : 32'd32892,	reg_addr : 32'd267542},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267543},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267544},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267545},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267546},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267547},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267548},
'{step_type : REG_WRITE,	value : 32'd67108865,	reg_addr : 32'd267549},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267550},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267551},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267552},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267553},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267554},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267555},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267556},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267557},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267558},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267559},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267560},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267561},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267562},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267563},
'{step_type : REG_WRITE,	value : 32'd218120236,	reg_addr : 32'd267564},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267565},
'{step_type : REG_WRITE,	value : 32'd134234192,	reg_addr : 32'd267566},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267567},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267568},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267569},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267570},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267571},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267572},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267573},
'{step_type : REG_WRITE,	value : 32'd134430800,	reg_addr : 32'd267574},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267575},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267576},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267577},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267578},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267579},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267580},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267581},
'{step_type : REG_WRITE,	value : 32'd134430800,	reg_addr : 32'd267582},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267583},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267584},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267585},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267586},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267587},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267588},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267589},
'{step_type : REG_WRITE,	value : 32'd134234192,	reg_addr : 32'd267590},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267591},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267592},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267593},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267594},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267595},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267596},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267597},
'{step_type : REG_WRITE,	value : 32'd16508,	reg_addr : 32'd267598},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267599},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267600},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267601},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267602},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267603},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267604},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267605},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267606},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267607},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267608},
'{step_type : REG_WRITE,	value : 32'd1526726656,	reg_addr : 32'd267609},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267610},
'{step_type : REG_WRITE,	value : 32'd469762048,	reg_addr : 32'd267611},
'{step_type : REG_WRITE,	value : 32'd218136620,	reg_addr : 32'd267612},
'{step_type : REG_WRITE,	value : 32'd1048577,	reg_addr : 32'd267613},
'{step_type : REG_WRITE,	value : 32'd134250576,	reg_addr : 32'd267614},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267615},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267616},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267617},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267618},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267619},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267620},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267621},
'{step_type : REG_WRITE,	value : 32'd134447184,	reg_addr : 32'd267622},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267623},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267624},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267625},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267626},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267627},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267628},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267629},
'{step_type : REG_WRITE,	value : 32'd134447184,	reg_addr : 32'd267630},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267631},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267632},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267633},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267634},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267635},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267636},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267637},
'{step_type : REG_WRITE,	value : 32'd134250576,	reg_addr : 32'd267638},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267639},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267640},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267641},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267642},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267643},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267644},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267645},
'{step_type : REG_WRITE,	value : 32'd32892,	reg_addr : 32'd267646},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267647},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267648},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267649},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267650},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267651},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267652},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267653},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267654},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267655},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267656},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd267657},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267658},
'{step_type : REG_WRITE,	value : 32'd671088640,	reg_addr : 32'd267659},
'{step_type : REG_WRITE,	value : 32'd218120236,	reg_addr : 32'd267660},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267661},
'{step_type : REG_WRITE,	value : 32'd134435224,	reg_addr : 32'd267662},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267663},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267664},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267665},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267666},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267667},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267668},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267669},
'{step_type : REG_WRITE,	value : 32'd134435352,	reg_addr : 32'd267670},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267671},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267672},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267673},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267674},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267675},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267676},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267677},
'{step_type : REG_WRITE,	value : 32'd16508,	reg_addr : 32'd267678},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267679},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267680},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267681},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267682},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267683},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267684},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267685},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267686},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267687},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267688},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267689},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267690},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267691},
'{step_type : REG_WRITE,	value : 32'd218136620,	reg_addr : 32'd267692},
'{step_type : REG_WRITE,	value : 32'd1048577,	reg_addr : 32'd267693},
'{step_type : REG_WRITE,	value : 32'd134451608,	reg_addr : 32'd267694},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267695},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267696},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267697},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267698},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267699},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267700},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267701},
'{step_type : REG_WRITE,	value : 32'd134451736,	reg_addr : 32'd267702},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267703},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267704},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267705},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267706},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267707},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267708},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267709},
'{step_type : REG_WRITE,	value : 32'd32892,	reg_addr : 32'd267710},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267711},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267712},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267713},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267714},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267715},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267716},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267717},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267718},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267719},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267720},
'{step_type : REG_WRITE,	value : 32'd989855744,	reg_addr : 32'd267721},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267722},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267723},
'{step_type : REG_WRITE,	value : 32'd53976,	reg_addr : 32'd267724},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267725},
'{step_type : REG_WRITE,	value : 32'd57352,	reg_addr : 32'd267726},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267727},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267728},
'{step_type : REG_WRITE,	value : 32'd2063597568,	reg_addr : 32'd267729},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267730},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267731},
'{step_type : REG_WRITE,	value : 32'd49392,	reg_addr : 32'd267732},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267733},
'{step_type : REG_WRITE,	value : 32'd53208,	reg_addr : 32'd267734},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267735},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267736},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267737},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267738},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267739},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267740},
'{step_type : REG_WRITE,	value : 32'd989855744,	reg_addr : 32'd267741},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267742},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267743},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267744},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267745},
'{step_type : REG_WRITE,	value : 32'd53336,	reg_addr : 32'd267746},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267747},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267748},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267749},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267750},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267751},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267752},
'{step_type : REG_WRITE,	value : 32'd989855744,	reg_addr : 32'd267753},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267754},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267755},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267756},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267757},
'{step_type : REG_WRITE,	value : 32'd53464,	reg_addr : 32'd267758},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267759},
'{step_type : REG_WRITE,	value : 32'd49288,	reg_addr : 32'd267760},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267761},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267762},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267763},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267764},
'{step_type : REG_WRITE,	value : 32'd989855744,	reg_addr : 32'd267765},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267766},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267767},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267768},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267769},
'{step_type : REG_WRITE,	value : 32'd53592,	reg_addr : 32'd267770},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267771},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267772},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267773},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267774},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267775},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267776},
'{step_type : REG_WRITE,	value : 32'd1795162112,	reg_addr : 32'd267777},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267778},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267779},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267780},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267781},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267782},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267783},
'{step_type : REG_WRITE,	value : 32'd218120236,	reg_addr : 32'd267784},
'{step_type : REG_WRITE,	value : 32'd67108865,	reg_addr : 32'd267785},
'{step_type : REG_WRITE,	value : 32'd134234192,	reg_addr : 32'd267786},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267787},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267788},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267789},
'{step_type : REG_WRITE,	value : 32'd134430800,	reg_addr : 32'd267790},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267791},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267792},
'{step_type : REG_WRITE,	value : 32'd1325400064,	reg_addr : 32'd267793},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267794},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267795},
'{step_type : REG_WRITE,	value : 32'd16508,	reg_addr : 32'd267796},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267797},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267798},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267799},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267800},
'{step_type : REG_WRITE,	value : 32'd520093696,	reg_addr : 32'd267801},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267802},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267803},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267804},
'{step_type : REG_WRITE,	value : 32'd67108865,	reg_addr : 32'd267805},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267806},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267807},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267808},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267809},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267810},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267811},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267812},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267813},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267814},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267815},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267816},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267817},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267818},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267819},
'{step_type : REG_WRITE,	value : 32'd218136620,	reg_addr : 32'd267820},
'{step_type : REG_WRITE,	value : 32'd68157441,	reg_addr : 32'd267821},
'{step_type : REG_WRITE,	value : 32'd134250576,	reg_addr : 32'd267822},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267823},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267824},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267825},
'{step_type : REG_WRITE,	value : 32'd134447184,	reg_addr : 32'd267826},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267827},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267828},
'{step_type : REG_WRITE,	value : 32'd1325400064,	reg_addr : 32'd267829},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267830},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267831},
'{step_type : REG_WRITE,	value : 32'd32892,	reg_addr : 32'd267832},
'{step_type : REG_WRITE,	value : 32'd68157440,	reg_addr : 32'd267833},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267834},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267835},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267836},
'{step_type : REG_WRITE,	value : 32'd520093696,	reg_addr : 32'd267837},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267838},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267839},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267840},
'{step_type : REG_WRITE,	value : 32'd67108865,	reg_addr : 32'd267841},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267842},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267843},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267844},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd267845},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267846},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267847},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267848},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267849},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267850},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267851},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267852},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267853},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267854},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267855},
'{step_type : REG_WRITE,	value : 32'd218120236,	reg_addr : 32'd267856},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267857},
'{step_type : REG_WRITE,	value : 32'd134234192,	reg_addr : 32'd267858},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267859},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267860},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267861},
'{step_type : REG_WRITE,	value : 32'd134430800,	reg_addr : 32'd267862},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267863},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267864},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267865},
'{step_type : REG_WRITE,	value : 32'd134430800,	reg_addr : 32'd267866},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267867},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267868},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267869},
'{step_type : REG_WRITE,	value : 32'd134234192,	reg_addr : 32'd267870},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267871},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267872},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd267873},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267874},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267875},
'{step_type : REG_WRITE,	value : 32'd16508,	reg_addr : 32'd267876},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267877},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267878},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267879},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267880},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267881},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267882},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267883},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267884},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267885},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267886},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267887},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267888},
'{step_type : REG_WRITE,	value : 32'd1526726656,	reg_addr : 32'd267889},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267890},
'{step_type : REG_WRITE,	value : 32'd469762048,	reg_addr : 32'd267891},
'{step_type : REG_WRITE,	value : 32'd218136620,	reg_addr : 32'd267892},
'{step_type : REG_WRITE,	value : 32'd1048577,	reg_addr : 32'd267893},
'{step_type : REG_WRITE,	value : 32'd134250576,	reg_addr : 32'd267894},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267895},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267896},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267897},
'{step_type : REG_WRITE,	value : 32'd134447184,	reg_addr : 32'd267898},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267899},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267900},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267901},
'{step_type : REG_WRITE,	value : 32'd134447184,	reg_addr : 32'd267902},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267903},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267904},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267905},
'{step_type : REG_WRITE,	value : 32'd134250576,	reg_addr : 32'd267906},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267907},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267908},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd267909},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267910},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267911},
'{step_type : REG_WRITE,	value : 32'd32892,	reg_addr : 32'd267912},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267913},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267914},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267915},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267916},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267917},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267918},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267919},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267920},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267921},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267922},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267923},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267924},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267925},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267926},
'{step_type : REG_WRITE,	value : 32'd671088640,	reg_addr : 32'd267927},
'{step_type : REG_WRITE,	value : 32'd218120236,	reg_addr : 32'd267928},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267929},
'{step_type : REG_WRITE,	value : 32'd134435224,	reg_addr : 32'd267930},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267931},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267932},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267933},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267934},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267935},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267936},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267937},
'{step_type : REG_WRITE,	value : 32'd134435352,	reg_addr : 32'd267938},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267939},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267940},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd267941},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267942},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267943},
'{step_type : REG_WRITE,	value : 32'd16508,	reg_addr : 32'd267944},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267945},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267946},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267947},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267948},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267949},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267950},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267951},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267952},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267953},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267954},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267955},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267956},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267957},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267958},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267959},
'{step_type : REG_WRITE,	value : 32'd218136620,	reg_addr : 32'd267960},
'{step_type : REG_WRITE,	value : 32'd1048577,	reg_addr : 32'd267961},
'{step_type : REG_WRITE,	value : 32'd134451608,	reg_addr : 32'd267962},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267963},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267964},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267965},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267966},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267967},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267968},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267969},
'{step_type : REG_WRITE,	value : 32'd134451736,	reg_addr : 32'd267970},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267971},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267972},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd267973},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267974},
'{step_type : REG_WRITE,	value : 32'd134217728,	reg_addr : 32'd267975},
'{step_type : REG_WRITE,	value : 32'd32892,	reg_addr : 32'd267976},
'{step_type : REG_WRITE,	value : 32'd1048576,	reg_addr : 32'd267977},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267978},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267979},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267980},
'{step_type : REG_WRITE,	value : 32'd452984832,	reg_addr : 32'd267981},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267982},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267983},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267984},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd267985},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267986},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267987},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267988},
'{step_type : REG_WRITE,	value : 32'd1795162112,	reg_addr : 32'd267989},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267990},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267991},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267992},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267993},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267994},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267995},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267996},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267997},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267998},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267999},
'{step_type : REG_WRITE,	value : 32'd1065006208,	reg_addr : 32'd278528},
'{step_type : REG_WRITE,	value : 32'd91168,	reg_addr : 32'd278529},
'{step_type : REG_WRITE,	value : 32'd1024,	reg_addr : 32'd278530},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278531},
'{step_type : REG_WRITE,	value : 32'd2147484800,	reg_addr : 32'd278532},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd278533},
'{step_type : REG_WRITE,	value : 32'd67111936,	reg_addr : 32'd278534},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278535},
'{step_type : REG_WRITE,	value : 32'd2214593664,	reg_addr : 32'd278536},
'{step_type : REG_WRITE,	value : 32'd3072,	reg_addr : 32'd278537},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278538},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278539},
'{step_type : REG_WRITE,	value : 32'd2214592640,	reg_addr : 32'd278540},
'{step_type : REG_WRITE,	value : 32'd3072,	reg_addr : 32'd278541},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278542},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278543},
'{step_type : REG_WRITE,	value : 32'd2147910144,	reg_addr : 32'd278544},
'{step_type : REG_WRITE,	value : 32'd16399,	reg_addr : 32'd278545},
'{step_type : REG_WRITE,	value : 32'd35136,	reg_addr : 32'd278546},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278547},
'{step_type : REG_WRITE,	value : 32'd2684355712,	reg_addr : 32'd278548},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd278549},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278550},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278551},
'{step_type : REG_WRITE,	value : 32'd2617253024,	reg_addr : 32'd278552},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278553},
'{step_type : REG_WRITE,	value : 32'd2818574464,	reg_addr : 32'd278554},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd278555},
'{step_type : REG_WRITE,	value : 32'd2147549312,	reg_addr : 32'd278556},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278557},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278558},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278559},
'{step_type : REG_WRITE,	value : 32'd2147550336,	reg_addr : 32'd278560},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278561},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278562},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278563},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd278564},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd278565},
'{step_type : REG_WRITE,	value : 32'd2684354688,	reg_addr : 32'd278566},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd278567},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd278568},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278569},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd278570},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278571},
'{step_type : REG_WRITE,	value : 32'd12320,	reg_addr : 32'd278572},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278573},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd278574},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278575},
'{step_type : REG_WRITE,	value : 32'd2818574464,	reg_addr : 32'd278576},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd278577},
'{step_type : REG_WRITE,	value : 32'd2147551360,	reg_addr : 32'd278578},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278579},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278580},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278581},
'{step_type : REG_WRITE,	value : 32'd2147552384,	reg_addr : 32'd278582},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278583},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278584},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278585},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd278586},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278587},
'{step_type : REG_WRITE,	value : 32'd11296,	reg_addr : 32'd278588},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278589},
'{step_type : REG_WRITE,	value : 32'd11296,	reg_addr : 32'd278590},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278591},
'{step_type : REG_WRITE,	value : 32'd11296,	reg_addr : 32'd278592},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278593},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd278594},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278595},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278596},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278597},
'{step_type : REG_WRITE,	value : 32'd2818573440,	reg_addr : 32'd278598},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278599},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278600},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278601},
'{step_type : REG_WRITE,	value : 32'd1073758720,	reg_addr : 32'd278602},
'{step_type : REG_WRITE,	value : 32'd16384,	reg_addr : 32'd278603},
'{step_type : REG_WRITE,	value : 32'd68928,	reg_addr : 32'd278604},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278605},
'{step_type : REG_WRITE,	value : 32'd3355457696,	reg_addr : 32'd278606},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278607},
'{step_type : REG_WRITE,	value : 32'd3422567584,	reg_addr : 32'd278608},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278609},
'{step_type : REG_WRITE,	value : 32'd2751463584,	reg_addr : 32'd278610},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd278611},
'{step_type : REG_WRITE,	value : 32'd2818579584,	reg_addr : 32'd278612},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd278613},
'{step_type : REG_WRITE,	value : 32'd2147815552,	reg_addr : 32'd278614},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278615},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278616},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278617},
'{step_type : REG_WRITE,	value : 32'd2147816576,	reg_addr : 32'd278618},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278619},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278620},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278621},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd278622},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd278623},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd278624},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278625},
'{step_type : REG_WRITE,	value : 32'd3422552192,	reg_addr : 32'd278626},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278627},
'{step_type : REG_WRITE,	value : 32'd2818579584,	reg_addr : 32'd278628},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd278629},
'{step_type : REG_WRITE,	value : 32'd2147817600,	reg_addr : 32'd278630},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278631},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278632},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278633},
'{step_type : REG_WRITE,	value : 32'd2147818624,	reg_addr : 32'd278634},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278635},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278636},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278637},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd278638},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd278639},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd278640},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278641},
'{step_type : REG_WRITE,	value : 32'd3355443328,	reg_addr : 32'd278642},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278643},
'{step_type : REG_WRITE,	value : 32'd3422567584,	reg_addr : 32'd278644},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278645},
'{step_type : REG_WRITE,	value : 32'd2818579584,	reg_addr : 32'd278646},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd278647},
'{step_type : REG_WRITE,	value : 32'd2147819648,	reg_addr : 32'd278648},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278649},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278650},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278651},
'{step_type : REG_WRITE,	value : 32'd2147820672,	reg_addr : 32'd278652},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278653},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278654},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278655},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd278656},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd278657},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd278658},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278659},
'{step_type : REG_WRITE,	value : 32'd3355457696,	reg_addr : 32'd278660},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278661},
'{step_type : REG_WRITE,	value : 32'd1409286289,	reg_addr : 32'd278662},
'{step_type : REG_WRITE,	value : 32'd102336,	reg_addr : 32'd278663},
'{step_type : REG_WRITE,	value : 32'd1409286289,	reg_addr : 32'd278664},
'{step_type : REG_WRITE,	value : 32'd85952,	reg_addr : 32'd278665},
'{step_type : REG_WRITE,	value : 32'd4026531985,	reg_addr : 32'd278666},
'{step_type : REG_WRITE,	value : 32'd100289,	reg_addr : 32'd278667},
'{step_type : REG_WRITE,	value : 32'd4026531985,	reg_addr : 32'd278668},
'{step_type : REG_WRITE,	value : 32'd83905,	reg_addr : 32'd278669},
'{step_type : REG_WRITE,	value : 32'd134219281,	reg_addr : 32'd278670},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd278671},
'{step_type : REG_WRITE,	value : 32'd80241,	reg_addr : 32'd278672},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278673},
'{step_type : REG_WRITE,	value : 32'd67111185,	reg_addr : 32'd278674},
'{step_type : REG_WRITE,	value : 32'd107552,	reg_addr : 32'd278675},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd278676},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278677},
'{step_type : REG_WRITE,	value : 32'd2577,	reg_addr : 32'd278678},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd278679},
'{step_type : REG_WRITE,	value : 32'd94545,	reg_addr : 32'd278680},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278681},
'{step_type : REG_WRITE,	value : 32'd82289,	reg_addr : 32'd278682},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278683},
'{step_type : REG_WRITE,	value : 32'd1553,	reg_addr : 32'd278684},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd278685},
'{step_type : REG_WRITE,	value : 32'd94577,	reg_addr : 32'd278686},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278687},
'{step_type : REG_WRITE,	value : 32'd603980945,	reg_addr : 32'd278688},
'{step_type : REG_WRITE,	value : 32'd123936,	reg_addr : 32'd278689},
'{step_type : REG_WRITE,	value : 32'd8657,	reg_addr : 32'd278690},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278691},
'{step_type : REG_WRITE,	value : 32'd4145,	reg_addr : 32'd278692},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278693},
'{step_type : REG_WRITE,	value : 32'd4145,	reg_addr : 32'd278694},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278695},
'{step_type : REG_WRITE,	value : 32'd11313,	reg_addr : 32'd278696},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278697},
'{step_type : REG_WRITE,	value : 32'd2818572433,	reg_addr : 32'd278698},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd278699},
'{step_type : REG_WRITE,	value : 32'd2147575953,	reg_addr : 32'd278700},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278701},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278702},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278703},
'{step_type : REG_WRITE,	value : 32'd2147576977,	reg_addr : 32'd278704},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278705},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278706},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278707},
'{step_type : REG_WRITE,	value : 32'd2129,	reg_addr : 32'd278708},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd278709},
'{step_type : REG_WRITE,	value : 32'd2147483793,	reg_addr : 32'd278710},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278711},
'{step_type : REG_WRITE,	value : 32'd2818572416,	reg_addr : 32'd278712},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278713},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278714},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278715},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278716},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278717},
'{step_type : REG_WRITE,	value : 32'd2818572416,	reg_addr : 32'd278718},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd278719},
'{step_type : REG_WRITE,	value : 32'd2147559552,	reg_addr : 32'd278720},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278721},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278722},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278723},
'{step_type : REG_WRITE,	value : 32'd2147560576,	reg_addr : 32'd278724},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278725},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278726},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278727},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd278728},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd278729},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd278730},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd278731},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278732},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278733},
'{step_type : REG_WRITE,	value : 32'd524800,	reg_addr : 32'd278734},
'{step_type : REG_WRITE,	value : 32'd16398,	reg_addr : 32'd278735},
'{step_type : REG_WRITE,	value : 32'd110912,	reg_addr : 32'd278736},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278737},
'{step_type : REG_WRITE,	value : 32'd131584,	reg_addr : 32'd278738},
'{step_type : REG_WRITE,	value : 32'd16398,	reg_addr : 32'd278739},
'{step_type : REG_WRITE,	value : 32'd110912,	reg_addr : 32'd278740},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278741},
'{step_type : REG_WRITE,	value : 32'd2147910144,	reg_addr : 32'd278742},
'{step_type : REG_WRITE,	value : 32'd16399,	reg_addr : 32'd278743},
'{step_type : REG_WRITE,	value : 32'd805309632,	reg_addr : 32'd278744},
'{step_type : REG_WRITE,	value : 32'd1988,	reg_addr : 32'd278745},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278746},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278747},
'{step_type : REG_WRITE,	value : 32'd1050112,	reg_addr : 32'd278748},
'{step_type : REG_WRITE,	value : 32'd16,	reg_addr : 32'd278749},
'{step_type : REG_WRITE,	value : 32'd738198720,	reg_addr : 32'd278750},
'{step_type : REG_WRITE,	value : 32'd960,	reg_addr : 32'd278751},
'{step_type : REG_WRITE,	value : 32'd2348820640,	reg_addr : 32'd278752},
'{step_type : REG_WRITE,	value : 32'd97217,	reg_addr : 32'd278753},
'{step_type : REG_WRITE,	value : 32'd2684355712,	reg_addr : 32'd278754},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd278755},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278756},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278757},
'{step_type : REG_WRITE,	value : 32'd2348815520,	reg_addr : 32'd278758},
'{step_type : REG_WRITE,	value : 32'd82881,	reg_addr : 32'd278759},
'{step_type : REG_WRITE,	value : 32'd2684354688,	reg_addr : 32'd278760},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd278761},
'{step_type : REG_WRITE,	value : 32'd2013267072,	reg_addr : 32'd278762},
'{step_type : REG_WRITE,	value : 32'd984,	reg_addr : 32'd278763},
'{step_type : REG_WRITE,	value : 32'd2080375936,	reg_addr : 32'd278764},
'{step_type : REG_WRITE,	value : 32'd2040,	reg_addr : 32'd278765},
'{step_type : REG_WRITE,	value : 32'd134217856,	reg_addr : 32'd278766},
'{step_type : REG_WRITE,	value : 32'd4064,	reg_addr : 32'd278767},
'{step_type : REG_WRITE,	value : 32'd134217856,	reg_addr : 32'd278768},
'{step_type : REG_WRITE,	value : 32'd2016,	reg_addr : 32'd278769},
'{step_type : REG_WRITE,	value : 32'd525824,	reg_addr : 32'd278770},
'{step_type : REG_WRITE,	value : 32'd8,	reg_addr : 32'd278771},
'{step_type : REG_WRITE,	value : 32'd1216,	reg_addr : 32'd278772},
'{step_type : REG_WRITE,	value : 32'd85956,	reg_addr : 32'd278773},
'{step_type : REG_WRITE,	value : 32'd1216,	reg_addr : 32'd278774},
'{step_type : REG_WRITE,	value : 32'd83908,	reg_addr : 32'd278775},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd278776},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278777},
'{step_type : REG_WRITE,	value : 32'd134218880,	reg_addr : 32'd278778},
'{step_type : REG_WRITE,	value : 32'd4064,	reg_addr : 32'd278779},
'{step_type : REG_WRITE,	value : 32'd134218880,	reg_addr : 32'd278780},
'{step_type : REG_WRITE,	value : 32'd2016,	reg_addr : 32'd278781},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd278782},
'{step_type : REG_WRITE,	value : 32'd85956,	reg_addr : 32'd278783},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd278784},
'{step_type : REG_WRITE,	value : 32'd83908,	reg_addr : 32'd278785},
'{step_type : REG_WRITE,	value : 32'd2013266048,	reg_addr : 32'd278786},
'{step_type : REG_WRITE,	value : 32'd984,	reg_addr : 32'd278787},
'{step_type : REG_WRITE,	value : 32'd2080374912,	reg_addr : 32'd278788},
'{step_type : REG_WRITE,	value : 32'd2040,	reg_addr : 32'd278789},
'{step_type : REG_WRITE,	value : 32'd2348821664,	reg_addr : 32'd278790},
'{step_type : REG_WRITE,	value : 32'd97217,	reg_addr : 32'd278791},
'{step_type : REG_WRITE,	value : 32'd2684355712,	reg_addr : 32'd278792},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd278793},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278794},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278795},
'{step_type : REG_WRITE,	value : 32'd2348816544,	reg_addr : 32'd278796},
'{step_type : REG_WRITE,	value : 32'd82881,	reg_addr : 32'd278797},
'{step_type : REG_WRITE,	value : 32'd2684354688,	reg_addr : 32'd278798},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd278799},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd278800},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278801},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd278802},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd278803},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd278804},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd278805},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd278806},
'{step_type : REG_WRITE,	value : 32'd192,	reg_addr : 32'd278807},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd278808},
'{step_type : REG_WRITE,	value : 32'd256,	reg_addr : 32'd278809},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd278810},
'{step_type : REG_WRITE,	value : 32'd320,	reg_addr : 32'd278811},
'{step_type : REG_WRITE,	value : 32'd2098688,	reg_addr : 32'd278812},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd278813},
'{step_type : REG_WRITE,	value : 32'd738197696,	reg_addr : 32'd278814},
'{step_type : REG_WRITE,	value : 32'd448,	reg_addr : 32'd278815},
'{step_type : REG_WRITE,	value : 32'd738197696,	reg_addr : 32'd278816},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd278817},
'{step_type : REG_WRITE,	value : 32'd738197696,	reg_addr : 32'd278818},
'{step_type : REG_WRITE,	value : 32'd576,	reg_addr : 32'd278819},
'{step_type : REG_WRITE,	value : 32'd738197696,	reg_addr : 32'd278820},
'{step_type : REG_WRITE,	value : 32'd640,	reg_addr : 32'd278821},
'{step_type : REG_WRITE,	value : 32'd738197696,	reg_addr : 32'd278822},
'{step_type : REG_WRITE,	value : 32'd704,	reg_addr : 32'd278823},
'{step_type : REG_WRITE,	value : 32'd738197696,	reg_addr : 32'd278824},
'{step_type : REG_WRITE,	value : 32'd768,	reg_addr : 32'd278825},
'{step_type : REG_WRITE,	value : 32'd3288336512,	reg_addr : 32'd278826},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd278827},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278828},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278829},
'{step_type : REG_WRITE,	value : 32'd201327744,	reg_addr : 32'd278830},
'{step_type : REG_WRITE,	value : 32'd4036,	reg_addr : 32'd278831},
'{step_type : REG_WRITE,	value : 32'd67117056,	reg_addr : 32'd278832},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278833},
'{step_type : REG_WRITE,	value : 32'd201327744,	reg_addr : 32'd278834},
'{step_type : REG_WRITE,	value : 32'd1988,	reg_addr : 32'd278835},
'{step_type : REG_WRITE,	value : 32'd67117056,	reg_addr : 32'd278836},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278837},
'{step_type : REG_WRITE,	value : 32'd201326720,	reg_addr : 32'd278838},
'{step_type : REG_WRITE,	value : 32'd4036,	reg_addr : 32'd278839},
'{step_type : REG_WRITE,	value : 32'd201326720,	reg_addr : 32'd278840},
'{step_type : REG_WRITE,	value : 32'd1988,	reg_addr : 32'd278841},
'{step_type : REG_WRITE,	value : 32'd3288334464,	reg_addr : 32'd278842},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd278843},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278844},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278845},
'{step_type : REG_WRITE,	value : 32'd3758097536,	reg_addr : 32'd278846},
'{step_type : REG_WRITE,	value : 32'd2051,	reg_addr : 32'd278847},
'{step_type : REG_WRITE,	value : 32'd67117056,	reg_addr : 32'd278848},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278849},
'{step_type : REG_WRITE,	value : 32'd67110400,	reg_addr : 32'd278850},
'{step_type : REG_WRITE,	value : 32'd1024,	reg_addr : 32'd278851},
'{step_type : REG_WRITE,	value : 32'd643455168,	reg_addr : 32'd278852},
'{step_type : REG_WRITE,	value : 32'd100296,	reg_addr : 32'd278853},
'{step_type : REG_WRITE,	value : 32'd1476395136,	reg_addr : 32'd278854},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd278855},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278856},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278857},
'{step_type : REG_WRITE,	value : 32'd3758096512,	reg_addr : 32'd278858},
'{step_type : REG_WRITE,	value : 32'd2051,	reg_addr : 32'd278859},
'{step_type : REG_WRITE,	value : 32'd67117056,	reg_addr : 32'd278860},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278861},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278862},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278863},
'{step_type : REG_WRITE,	value : 32'd1342177408,	reg_addr : 32'd278864},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278865},
'{step_type : REG_WRITE,	value : 32'd1073742976,	reg_addr : 32'd278866},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd278867},
'{step_type : REG_WRITE,	value : 32'd3288334464,	reg_addr : 32'd278868},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd278869},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd278870},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd278871},
'{step_type : REG_WRITE,	value : 32'd2350907520,	reg_addr : 32'd278872},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd278873},
'{step_type : REG_WRITE,	value : 32'd2098688,	reg_addr : 32'd278874},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd278875},
'{step_type : REG_WRITE,	value : 32'd2282487936,	reg_addr : 32'd278876},
'{step_type : REG_WRITE,	value : 32'd3074,	reg_addr : 32'd278877},
'{step_type : REG_WRITE,	value : 32'd2282488000,	reg_addr : 32'd278878},
'{step_type : REG_WRITE,	value : 32'd3138,	reg_addr : 32'd278879},
'{step_type : REG_WRITE,	value : 32'd612367488,	reg_addr : 32'd278880},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd278881},
'{step_type : REG_WRITE,	value : 32'd673184896,	reg_addr : 32'd278882},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd278883},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278884},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278885},
'{step_type : REG_WRITE,	value : 32'd2148270208,	reg_addr : 32'd278886},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd278887},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278888},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278889},
'{step_type : REG_WRITE,	value : 32'd2550137984,	reg_addr : 32'd278890},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd278891},
'{step_type : REG_WRITE,	value : 32'd671089792,	reg_addr : 32'd278892},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd278893},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd278894},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278895},
'{step_type : REG_WRITE,	value : 32'd2164259968,	reg_addr : 32'd278896},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd278897},
'{step_type : REG_WRITE,	value : 32'd805306496,	reg_addr : 32'd278898},
'{step_type : REG_WRITE,	value : 32'd1988,	reg_addr : 32'd278899},
'{step_type : REG_WRITE,	value : 32'd67072,	reg_addr : 32'd278900},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd278901},
'{step_type : REG_WRITE,	value : 32'd194880,	reg_addr : 32'd278902},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278903},
'{step_type : REG_WRITE,	value : 32'd2147910144,	reg_addr : 32'd278904},
'{step_type : REG_WRITE,	value : 32'd16399,	reg_addr : 32'd278905},
'{step_type : REG_WRITE,	value : 32'd195936,	reg_addr : 32'd278906},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278907},
'{step_type : REG_WRITE,	value : 32'd105920,	reg_addr : 32'd278908},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278909},
'{step_type : REG_WRITE,	value : 32'd3758097536,	reg_addr : 32'd278910},
'{step_type : REG_WRITE,	value : 32'd2051,	reg_addr : 32'd278911},
'{step_type : REG_WRITE,	value : 32'd67116032,	reg_addr : 32'd278912},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278913},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd278914},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd278915},
'{step_type : REG_WRITE,	value : 32'd2281702528,	reg_addr : 32'd278916},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd278917},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd278918},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278919},
'{step_type : REG_WRITE,	value : 32'd1543504000,	reg_addr : 32'd278920},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd278921},
'{step_type : REG_WRITE,	value : 32'd33555968,	reg_addr : 32'd278922},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd278923},
'{step_type : REG_WRITE,	value : 32'd738201792,	reg_addr : 32'd278924},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd278925},
'{step_type : REG_WRITE,	value : 32'd738203776,	reg_addr : 32'd278926},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd278927},
'{step_type : REG_WRITE,	value : 32'd402659456,	reg_addr : 32'd278928},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd278929},
'{step_type : REG_WRITE,	value : 32'd469768320,	reg_addr : 32'd278930},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd278931},
'{step_type : REG_WRITE,	value : 32'd536877184,	reg_addr : 32'd278932},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd278933},
'{step_type : REG_WRITE,	value : 32'd603986048,	reg_addr : 32'd278934},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd278935},
'{step_type : REG_WRITE,	value : 32'd671094912,	reg_addr : 32'd278936},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd278937},
'{step_type : REG_WRITE,	value : 32'd131584,	reg_addr : 32'd278938},
'{step_type : REG_WRITE,	value : 32'd16398,	reg_addr : 32'd278939},
'{step_type : REG_WRITE,	value : 32'd223552,	reg_addr : 32'd278940},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278941},
'{step_type : REG_WRITE,	value : 32'd1073759744,	reg_addr : 32'd278942},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278943},
'{step_type : REG_WRITE,	value : 32'd218432,	reg_addr : 32'd278944},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278945},
'{step_type : REG_WRITE,	value : 32'd67111168,	reg_addr : 32'd278946},
'{step_type : REG_WRITE,	value : 32'd107552,	reg_addr : 32'd278947},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd278948},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278949},
'{step_type : REG_WRITE,	value : 32'd1073760768,	reg_addr : 32'd278950},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278951},
'{step_type : REG_WRITE,	value : 32'd201330912,	reg_addr : 32'd278952},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd278953},
'{step_type : REG_WRITE,	value : 32'd201326784,	reg_addr : 32'd278954},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd278955},
'{step_type : REG_WRITE,	value : 32'd67110016,	reg_addr : 32'd278956},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd278957},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278958},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278959},
'{step_type : REG_WRITE,	value : 32'd134218880,	reg_addr : 32'd278960},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd278961},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd278962},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278963},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278964},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278965},
'{step_type : REG_WRITE,	value : 32'd2617248945,	reg_addr : 32'd278966},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278967},
'{step_type : REG_WRITE,	value : 32'd2617249969,	reg_addr : 32'd278968},
'{step_type : REG_WRITE,	value : 32'd7171,	reg_addr : 32'd278969},
'{step_type : REG_WRITE,	value : 32'd603979921,	reg_addr : 32'd278970},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278971},
'{step_type : REG_WRITE,	value : 32'd81,	reg_addr : 32'd278972},
'{step_type : REG_WRITE,	value : 32'd16384,	reg_addr : 32'd278973},
'{step_type : REG_WRITE,	value : 32'd233777,	reg_addr : 32'd278974},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278975},
'{step_type : REG_WRITE,	value : 32'd1073748481,	reg_addr : 32'd278976},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278977},
'{step_type : REG_WRITE,	value : 32'd233825,	reg_addr : 32'd278978},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278979},
'{step_type : REG_WRITE,	value : 32'd603979905,	reg_addr : 32'd278980},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd278981},
'{step_type : REG_WRITE,	value : 32'd65,	reg_addr : 32'd278982},
'{step_type : REG_WRITE,	value : 32'd16384,	reg_addr : 32'd278983},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278984},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278985},
'{step_type : REG_WRITE,	value : 32'd2214594816,	reg_addr : 32'd278986},
'{step_type : REG_WRITE,	value : 32'd9244,	reg_addr : 32'd278987},
'{step_type : REG_WRITE,	value : 32'd3221307904,	reg_addr : 32'd278988},
'{step_type : REG_WRITE,	value : 32'd49153,	reg_addr : 32'd278989},
'{step_type : REG_WRITE,	value : 32'd239936,	reg_addr : 32'd278990},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278991},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd278992},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278993},
'{step_type : REG_WRITE,	value : 32'd738199712,	reg_addr : 32'd278994},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd278995},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd278996},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd278997},
'{step_type : REG_WRITE,	value : 32'd1073742976,	reg_addr : 32'd278998},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd278999},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279000},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279001},
'{step_type : REG_WRITE,	value : 32'd67108992,	reg_addr : 32'd279002},
'{step_type : REG_WRITE,	value : 32'd11264,	reg_addr : 32'd279003},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279004},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279005},
'{step_type : REG_WRITE,	value : 32'd131584,	reg_addr : 32'd279006},
'{step_type : REG_WRITE,	value : 32'd16398,	reg_addr : 32'd279007},
'{step_type : REG_WRITE,	value : 32'd278848,	reg_addr : 32'd279008},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279009},
'{step_type : REG_WRITE,	value : 32'd1073759744,	reg_addr : 32'd279010},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279011},
'{step_type : REG_WRITE,	value : 32'd67110080,	reg_addr : 32'd279012},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279013},
'{step_type : REG_WRITE,	value : 32'd134218944,	reg_addr : 32'd279014},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279015},
'{step_type : REG_WRITE,	value : 32'd278848,	reg_addr : 32'd279016},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279017},
'{step_type : REG_WRITE,	value : 32'd134217856,	reg_addr : 32'd279018},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279019},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279020},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279021},
'{step_type : REG_WRITE,	value : 32'd67108992,	reg_addr : 32'd279022},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279023},
'{step_type : REG_WRITE,	value : 32'd129,	reg_addr : 32'd279024},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279025},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279026},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279027},
'{step_type : REG_WRITE,	value : 32'd2281702528,	reg_addr : 32'd279028},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279029},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279030},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279031},
'{step_type : REG_WRITE,	value : 32'd201328896,	reg_addr : 32'd279032},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279033},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279034},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279035},
'{step_type : REG_WRITE,	value : 32'd68096,	reg_addr : 32'd279036},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd279037},
'{step_type : REG_WRITE,	value : 32'd269632,	reg_addr : 32'd279038},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279039},
'{step_type : REG_WRITE,	value : 32'd201329792,	reg_addr : 32'd279040},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279041},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd279042},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279043},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd279044},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279045},
'{step_type : REG_WRITE,	value : 32'd201328768,	reg_addr : 32'd279046},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279047},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd279048},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279049},
'{step_type : REG_WRITE,	value : 32'd201326720,	reg_addr : 32'd279050},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279051},
'{step_type : REG_WRITE,	value : 32'd279840,	reg_addr : 32'd279052},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279053},
'{step_type : REG_WRITE,	value : 32'd201333888,	reg_addr : 32'd279054},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279055},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd279056},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279057},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd279058},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279059},
'{step_type : REG_WRITE,	value : 32'd201332864,	reg_addr : 32'd279060},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279061},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd279062},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279063},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd279064},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279065},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd279066},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279067},
'{step_type : REG_WRITE,	value : 32'd201330816,	reg_addr : 32'd279068},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279069},
'{step_type : REG_WRITE,	value : 32'd279840,	reg_addr : 32'd279070},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279071},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd279072},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279073},
'{step_type : REG_WRITE,	value : 32'd2098688,	reg_addr : 32'd279074},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd279075},
'{step_type : REG_WRITE,	value : 32'd302432,	reg_addr : 32'd279076},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279077},
'{step_type : REG_WRITE,	value : 32'd402653312,	reg_addr : 32'd279078},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279079},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279080},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279081},
'{step_type : REG_WRITE,	value : 32'd536871040,	reg_addr : 32'd279082},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279083},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279084},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279085},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279086},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279087},
'{step_type : REG_WRITE,	value : 32'd738199680,	reg_addr : 32'd279088},
'{step_type : REG_WRITE,	value : 32'd14337,	reg_addr : 32'd279089},
'{step_type : REG_WRITE,	value : 32'd738201728,	reg_addr : 32'd279090},
'{step_type : REG_WRITE,	value : 32'd14401,	reg_addr : 32'd279091},
'{step_type : REG_WRITE,	value : 32'd738199680,	reg_addr : 32'd279092},
'{step_type : REG_WRITE,	value : 32'd14465,	reg_addr : 32'd279093},
'{step_type : REG_WRITE,	value : 32'd738201728,	reg_addr : 32'd279094},
'{step_type : REG_WRITE,	value : 32'd14529,	reg_addr : 32'd279095},
'{step_type : REG_WRITE,	value : 32'd738199680,	reg_addr : 32'd279096},
'{step_type : REG_WRITE,	value : 32'd14593,	reg_addr : 32'd279097},
'{step_type : REG_WRITE,	value : 32'd738201728,	reg_addr : 32'd279098},
'{step_type : REG_WRITE,	value : 32'd14657,	reg_addr : 32'd279099},
'{step_type : REG_WRITE,	value : 32'd738199680,	reg_addr : 32'd279100},
'{step_type : REG_WRITE,	value : 32'd14721,	reg_addr : 32'd279101},
'{step_type : REG_WRITE,	value : 32'd738201728,	reg_addr : 32'd279102},
'{step_type : REG_WRITE,	value : 32'd14785,	reg_addr : 32'd279103},
'{step_type : REG_WRITE,	value : 32'd33555968,	reg_addr : 32'd279104},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd279105},
'{step_type : REG_WRITE,	value : 32'd738201792,	reg_addr : 32'd279106},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279107},
'{step_type : REG_WRITE,	value : 32'd1476395136,	reg_addr : 32'd279108},
'{step_type : REG_WRITE,	value : 32'd975,	reg_addr : 32'd279109},
'{step_type : REG_WRITE,	value : 32'd1543504000,	reg_addr : 32'd279110},
'{step_type : REG_WRITE,	value : 32'd975,	reg_addr : 32'd279111},
'{step_type : REG_WRITE,	value : 32'd1543506048,	reg_addr : 32'd279112},
'{step_type : REG_WRITE,	value : 32'd207,	reg_addr : 32'd279113},
'{step_type : REG_WRITE,	value : 32'd1543506048,	reg_addr : 32'd279114},
'{step_type : REG_WRITE,	value : 32'd655,	reg_addr : 32'd279115},
'{step_type : REG_WRITE,	value : 32'd338208,	reg_addr : 32'd279116},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279117},
'{step_type : REG_WRITE,	value : 32'd402653312,	reg_addr : 32'd279118},
'{step_type : REG_WRITE,	value : 32'd14337,	reg_addr : 32'd279119},
'{step_type : REG_WRITE,	value : 32'd402653312,	reg_addr : 32'd279120},
'{step_type : REG_WRITE,	value : 32'd14401,	reg_addr : 32'd279121},
'{step_type : REG_WRITE,	value : 32'd402653312,	reg_addr : 32'd279122},
'{step_type : REG_WRITE,	value : 32'd14465,	reg_addr : 32'd279123},
'{step_type : REG_WRITE,	value : 32'd402653312,	reg_addr : 32'd279124},
'{step_type : REG_WRITE,	value : 32'd14529,	reg_addr : 32'd279125},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279126},
'{step_type : REG_WRITE,	value : 32'd14337,	reg_addr : 32'd279127},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279128},
'{step_type : REG_WRITE,	value : 32'd14401,	reg_addr : 32'd279129},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279130},
'{step_type : REG_WRITE,	value : 32'd14465,	reg_addr : 32'd279131},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279132},
'{step_type : REG_WRITE,	value : 32'd14529,	reg_addr : 32'd279133},
'{step_type : REG_WRITE,	value : 32'd536871040,	reg_addr : 32'd279134},
'{step_type : REG_WRITE,	value : 32'd14337,	reg_addr : 32'd279135},
'{step_type : REG_WRITE,	value : 32'd536871040,	reg_addr : 32'd279136},
'{step_type : REG_WRITE,	value : 32'd14401,	reg_addr : 32'd279137},
'{step_type : REG_WRITE,	value : 32'd536871040,	reg_addr : 32'd279138},
'{step_type : REG_WRITE,	value : 32'd14465,	reg_addr : 32'd279139},
'{step_type : REG_WRITE,	value : 32'd536871040,	reg_addr : 32'd279140},
'{step_type : REG_WRITE,	value : 32'd14529,	reg_addr : 32'd279141},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279142},
'{step_type : REG_WRITE,	value : 32'd14337,	reg_addr : 32'd279143},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279144},
'{step_type : REG_WRITE,	value : 32'd14401,	reg_addr : 32'd279145},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279146},
'{step_type : REG_WRITE,	value : 32'd14465,	reg_addr : 32'd279147},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279148},
'{step_type : REG_WRITE,	value : 32'd14529,	reg_addr : 32'd279149},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279150},
'{step_type : REG_WRITE,	value : 32'd14401,	reg_addr : 32'd279151},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279152},
'{step_type : REG_WRITE,	value : 32'd14529,	reg_addr : 32'd279153},
'{step_type : REG_WRITE,	value : 32'd738199680,	reg_addr : 32'd279154},
'{step_type : REG_WRITE,	value : 32'd14337,	reg_addr : 32'd279155},
'{step_type : REG_WRITE,	value : 32'd738201728,	reg_addr : 32'd279156},
'{step_type : REG_WRITE,	value : 32'd14401,	reg_addr : 32'd279157},
'{step_type : REG_WRITE,	value : 32'd738199680,	reg_addr : 32'd279158},
'{step_type : REG_WRITE,	value : 32'd14465,	reg_addr : 32'd279159},
'{step_type : REG_WRITE,	value : 32'd738201728,	reg_addr : 32'd279160},
'{step_type : REG_WRITE,	value : 32'd14529,	reg_addr : 32'd279161},
'{step_type : REG_WRITE,	value : 32'd33555968,	reg_addr : 32'd279162},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd279163},
'{step_type : REG_WRITE,	value : 32'd738201792,	reg_addr : 32'd279164},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279165},
'{step_type : REG_WRITE,	value : 32'd1476395136,	reg_addr : 32'd279166},
'{step_type : REG_WRITE,	value : 32'd15,	reg_addr : 32'd279167},
'{step_type : REG_WRITE,	value : 32'd1543504000,	reg_addr : 32'd279168},
'{step_type : REG_WRITE,	value : 32'd15,	reg_addr : 32'd279169},
'{step_type : REG_WRITE,	value : 32'd1476395136,	reg_addr : 32'd279170},
'{step_type : REG_WRITE,	value : 32'd79,	reg_addr : 32'd279171},
'{step_type : REG_WRITE,	value : 32'd1543504000,	reg_addr : 32'd279172},
'{step_type : REG_WRITE,	value : 32'd79,	reg_addr : 32'd279173},
'{step_type : REG_WRITE,	value : 32'd1476395136,	reg_addr : 32'd279174},
'{step_type : REG_WRITE,	value : 32'd143,	reg_addr : 32'd279175},
'{step_type : REG_WRITE,	value : 32'd1543504000,	reg_addr : 32'd279176},
'{step_type : REG_WRITE,	value : 32'd143,	reg_addr : 32'd279177},
'{step_type : REG_WRITE,	value : 32'd1476395136,	reg_addr : 32'd279178},
'{step_type : REG_WRITE,	value : 32'd207,	reg_addr : 32'd279179},
'{step_type : REG_WRITE,	value : 32'd1476395136,	reg_addr : 32'd279180},
'{step_type : REG_WRITE,	value : 32'd271,	reg_addr : 32'd279181},
'{step_type : REG_WRITE,	value : 32'd1543504000,	reg_addr : 32'd279182},
'{step_type : REG_WRITE,	value : 32'd271,	reg_addr : 32'd279183},
'{step_type : REG_WRITE,	value : 32'd1476395136,	reg_addr : 32'd279184},
'{step_type : REG_WRITE,	value : 32'd335,	reg_addr : 32'd279185},
'{step_type : REG_WRITE,	value : 32'd1543504000,	reg_addr : 32'd279186},
'{step_type : REG_WRITE,	value : 32'd335,	reg_addr : 32'd279187},
'{step_type : REG_WRITE,	value : 32'd536871040,	reg_addr : 32'd279188},
'{step_type : REG_WRITE,	value : 32'd11212,	reg_addr : 32'd279189},
'{step_type : REG_WRITE,	value : 32'd342321,	reg_addr : 32'd279190},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279191},
'{step_type : REG_WRITE,	value : 32'd1073748480,	reg_addr : 32'd279192},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279193},
'{step_type : REG_WRITE,	value : 32'd342368,	reg_addr : 32'd279194},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279195},
'{step_type : REG_WRITE,	value : 32'd67121312,	reg_addr : 32'd279196},
'{step_type : REG_WRITE,	value : 32'd11264,	reg_addr : 32'd279197},
'{step_type : REG_WRITE,	value : 32'd2281701504,	reg_addr : 32'd279198},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279199},
'{step_type : REG_WRITE,	value : 32'd1545600128,	reg_addr : 32'd279200},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279201},
'{step_type : REG_WRITE,	value : 32'd8390144,	reg_addr : 32'd279202},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd279203},
'{step_type : REG_WRITE,	value : 32'd3154118912,	reg_addr : 32'd279204},
'{step_type : REG_WRITE,	value : 32'd93196,	reg_addr : 32'd279205},
'{step_type : REG_WRITE,	value : 32'd67109056,	reg_addr : 32'd279206},
'{step_type : REG_WRITE,	value : 32'd9252,	reg_addr : 32'd279207},
'{step_type : REG_WRITE,	value : 32'd67141856,	reg_addr : 32'd279208},
'{step_type : REG_WRITE,	value : 32'd9252,	reg_addr : 32'd279209},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd279210},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279211},
'{step_type : REG_WRITE,	value : 32'd2550144181,	reg_addr : 32'd279212},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279213},
'{step_type : REG_WRITE,	value : 32'd2617254069,	reg_addr : 32'd279214},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279215},
'{step_type : REG_WRITE,	value : 32'd2550136981,	reg_addr : 32'd279216},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279217},
'{step_type : REG_WRITE,	value : 32'd2617245845,	reg_addr : 32'd279218},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279219},
'{step_type : REG_WRITE,	value : 32'd1073741973,	reg_addr : 32'd279220},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279221},
'{step_type : REG_WRITE,	value : 32'd1541,	reg_addr : 32'd279222},
'{step_type : REG_WRITE,	value : 32'd8192,	reg_addr : 32'd279223},
'{step_type : REG_WRITE,	value : 32'd1073742021,	reg_addr : 32'd279224},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279225},
'{step_type : REG_WRITE,	value : 32'd2147484869,	reg_addr : 32'd279226},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279227},
'{step_type : REG_WRITE,	value : 32'd2147483845,	reg_addr : 32'd279228},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279229},
'{step_type : REG_WRITE,	value : 32'd67109093,	reg_addr : 32'd279230},
'{step_type : REG_WRITE,	value : 32'd11264,	reg_addr : 32'd279231},
'{step_type : REG_WRITE,	value : 32'd3154116837,	reg_addr : 32'd279232},
'{step_type : REG_WRITE,	value : 32'd93196,	reg_addr : 32'd279233},
'{step_type : REG_WRITE,	value : 32'd67108864,	reg_addr : 32'd279234},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279235},
'{step_type : REG_WRITE,	value : 32'd2617115877,	reg_addr : 32'd279236},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279237},
'{step_type : REG_WRITE,	value : 32'd2684224741,	reg_addr : 32'd279238},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279239},
'{step_type : REG_WRITE,	value : 32'd2617114853,	reg_addr : 32'd279240},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279241},
'{step_type : REG_WRITE,	value : 32'd2684223717,	reg_addr : 32'd279242},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279243},
'{step_type : REG_WRITE,	value : 32'd1073743077,	reg_addr : 32'd279244},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279245},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279246},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279247},
'{step_type : REG_WRITE,	value : 32'd3154118821,	reg_addr : 32'd279248},
'{step_type : REG_WRITE,	value : 32'd93196,	reg_addr : 32'd279249},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd279250},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279251},
'{step_type : REG_WRITE,	value : 32'd3892513920,	reg_addr : 32'd279252},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279253},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279254},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279255},
'{step_type : REG_WRITE,	value : 32'd3892314240,	reg_addr : 32'd279256},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279257},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd279258},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279259},
'{step_type : REG_WRITE,	value : 32'd2281701504,	reg_addr : 32'd279260},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279261},
'{step_type : REG_WRITE,	value : 32'd67111936,	reg_addr : 32'd279262},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279263},
'{step_type : REG_WRITE,	value : 32'd52352,	reg_addr : 32'd279264},
'{step_type : REG_WRITE,	value : 32'd2056,	reg_addr : 32'd279265},
'{step_type : REG_WRITE,	value : 32'd469763200,	reg_addr : 32'd279266},
'{step_type : REG_WRITE,	value : 32'd4033,	reg_addr : 32'd279267},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279268},
'{step_type : REG_WRITE,	value : 32'd4033,	reg_addr : 32'd279269},
'{step_type : REG_WRITE,	value : 32'd469763200,	reg_addr : 32'd279270},
'{step_type : REG_WRITE,	value : 32'd1985,	reg_addr : 32'd279271},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279272},
'{step_type : REG_WRITE,	value : 32'd1985,	reg_addr : 32'd279273},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd279274},
'{step_type : REG_WRITE,	value : 32'd2056,	reg_addr : 32'd279275},
'{step_type : REG_WRITE,	value : 32'd1342177408,	reg_addr : 32'd279276},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279277},
'{step_type : REG_WRITE,	value : 32'd3087008896,	reg_addr : 32'd279278},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279279},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279280},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279281},
'{step_type : REG_WRITE,	value : 32'd263680,	reg_addr : 32'd279282},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd279283},
'{step_type : REG_WRITE,	value : 32'd1501561056,	reg_addr : 32'd279284},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd279285},
'{step_type : REG_WRITE,	value : 32'd671089792,	reg_addr : 32'd279286},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279287},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279288},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279289},
'{step_type : REG_WRITE,	value : 32'd3758096512,	reg_addr : 32'd279290},
'{step_type : REG_WRITE,	value : 32'd2051,	reg_addr : 32'd279291},
'{step_type : REG_WRITE,	value : 32'd67113984,	reg_addr : 32'd279292},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279293},
'{step_type : REG_WRITE,	value : 32'd2281703552,	reg_addr : 32'd279294},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279295},
'{step_type : REG_WRITE,	value : 32'd3104,	reg_addr : 32'd279296},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279297},
'{step_type : REG_WRITE,	value : 32'd1073759744,	reg_addr : 32'd279298},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279299},
'{step_type : REG_WRITE,	value : 32'd396640,	reg_addr : 32'd279300},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279301},
'{step_type : REG_WRITE,	value : 32'd469764224,	reg_addr : 32'd279302},
'{step_type : REG_WRITE,	value : 32'd4033,	reg_addr : 32'd279303},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279304},
'{step_type : REG_WRITE,	value : 32'd4033,	reg_addr : 32'd279305},
'{step_type : REG_WRITE,	value : 32'd469764224,	reg_addr : 32'd279306},
'{step_type : REG_WRITE,	value : 32'd1985,	reg_addr : 32'd279307},
'{step_type : REG_WRITE,	value : 32'd469762176,	reg_addr : 32'd279308},
'{step_type : REG_WRITE,	value : 32'd1985,	reg_addr : 32'd279309},
'{step_type : REG_WRITE,	value : 32'd67124224,	reg_addr : 32'd279310},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279311},
'{step_type : REG_WRITE,	value : 32'd263680,	reg_addr : 32'd279312},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd279313},
'{step_type : REG_WRITE,	value : 32'd404800,	reg_addr : 32'd279314},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279315},
'{step_type : REG_WRITE,	value : 32'd113088,	reg_addr : 32'd279316},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279317},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279318},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279319},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279320},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279321},
'{step_type : REG_WRITE,	value : 32'd2550136960,	reg_addr : 32'd279322},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279323},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279324},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279325},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279326},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279327},
'{step_type : REG_WRITE,	value : 32'd2285633664,	reg_addr : 32'd279328},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279329},
'{step_type : REG_WRITE,	value : 32'd2147746304,	reg_addr : 32'd279330},
'{step_type : REG_WRITE,	value : 32'd16399,	reg_addr : 32'd279331},
'{step_type : REG_WRITE,	value : 32'd419136,	reg_addr : 32'd279332},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279333},
'{step_type : REG_WRITE,	value : 32'd524800,	reg_addr : 32'd279334},
'{step_type : REG_WRITE,	value : 32'd16398,	reg_addr : 32'd279335},
'{step_type : REG_WRITE,	value : 32'd419136,	reg_addr : 32'd279336},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279337},
'{step_type : REG_WRITE,	value : 32'd3825206400,	reg_addr : 32'd279338},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279339},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279340},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279341},
'{step_type : REG_WRITE,	value : 32'd3825205376,	reg_addr : 32'd279342},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279343},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279344},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279345},
'{step_type : REG_WRITE,	value : 32'd3892513921,	reg_addr : 32'd279346},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279347},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279348},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279349},
'{step_type : REG_WRITE,	value : 32'd3892314241,	reg_addr : 32'd279350},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279351},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279352},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279353},
'{step_type : REG_WRITE,	value : 32'd1073748481,	reg_addr : 32'd279354},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279355},
'{step_type : REG_WRITE,	value : 32'd430401,	reg_addr : 32'd279356},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279357},
'{step_type : REG_WRITE,	value : 32'd2684355713,	reg_addr : 32'd279358},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd279359},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279360},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279361},
'{step_type : REG_WRITE,	value : 32'd1073754625,	reg_addr : 32'd279362},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279363},
'{step_type : REG_WRITE,	value : 32'd438593,	reg_addr : 32'd279364},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279365},
'{step_type : REG_WRITE,	value : 32'd430433,	reg_addr : 32'd279366},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279367},
'{step_type : REG_WRITE,	value : 32'd7201,	reg_addr : 32'd279368},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279369},
'{step_type : REG_WRITE,	value : 32'd2684354689,	reg_addr : 32'd279370},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd279371},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279372},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279373},
'{step_type : REG_WRITE,	value : 32'd132609,	reg_addr : 32'd279374},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd279375},
'{step_type : REG_WRITE,	value : 32'd3892513985,	reg_addr : 32'd279376},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279377},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279378},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279379},
'{step_type : REG_WRITE,	value : 32'd3892314305,	reg_addr : 32'd279380},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279381},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279382},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279383},
'{step_type : REG_WRITE,	value : 32'd2684354689,	reg_addr : 32'd279384},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd279385},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279386},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279387},
'{step_type : REG_WRITE,	value : 32'd3892513937,	reg_addr : 32'd279388},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279389},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279390},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279391},
'{step_type : REG_WRITE,	value : 32'd3892314257,	reg_addr : 32'd279392},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279393},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279394},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279395},
'{step_type : REG_WRITE,	value : 32'd2818573440,	reg_addr : 32'd279396},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279397},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279398},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279399},
'{step_type : REG_WRITE,	value : 32'd402653313,	reg_addr : 32'd279400},
'{step_type : REG_WRITE,	value : 32'd123936,	reg_addr : 32'd279401},
'{step_type : REG_WRITE,	value : 32'd1073767953,	reg_addr : 32'd279402},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279403},
'{step_type : REG_WRITE,	value : 32'd450897,	reg_addr : 32'd279404},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279405},
'{step_type : REG_WRITE,	value : 32'd8657,	reg_addr : 32'd279406},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279407},
'{step_type : REG_WRITE,	value : 32'd2684355729,	reg_addr : 32'd279408},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd279409},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279410},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279411},
'{step_type : REG_WRITE,	value : 32'd1409294513,	reg_addr : 32'd279412},
'{step_type : REG_WRITE,	value : 32'd85952,	reg_addr : 32'd279413},
'{step_type : REG_WRITE,	value : 32'd4026541233,	reg_addr : 32'd279414},
'{step_type : REG_WRITE,	value : 32'd83905,	reg_addr : 32'd279415},
'{step_type : REG_WRITE,	value : 32'd2684354705,	reg_addr : 32'd279416},
'{step_type : REG_WRITE,	value : 32'd9248,	reg_addr : 32'd279417},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd279418},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279419},
'{step_type : REG_WRITE,	value : 32'd2818572416,	reg_addr : 32'd279420},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279421},
'{step_type : REG_WRITE,	value : 32'd2147561600,	reg_addr : 32'd279422},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279423},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279424},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279425},
'{step_type : REG_WRITE,	value : 32'd2147562624,	reg_addr : 32'd279426},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279427},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279428},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279429},
'{step_type : REG_WRITE,	value : 32'd67116032,	reg_addr : 32'd279430},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279431},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279432},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279433},
'{step_type : REG_WRITE,	value : 32'd1056,	reg_addr : 32'd279434},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279435},
'{step_type : REG_WRITE,	value : 32'd2818572416,	reg_addr : 32'd279436},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279437},
'{step_type : REG_WRITE,	value : 32'd2147563648,	reg_addr : 32'd279438},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279439},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279440},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279441},
'{step_type : REG_WRITE,	value : 32'd2147564672,	reg_addr : 32'd279442},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279443},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279444},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279445},
'{step_type : REG_WRITE,	value : 32'd67116032,	reg_addr : 32'd279446},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279447},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279448},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279449},
'{step_type : REG_WRITE,	value : 32'd1056,	reg_addr : 32'd279450},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279451},
'{step_type : REG_WRITE,	value : 32'd2818572416,	reg_addr : 32'd279452},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279453},
'{step_type : REG_WRITE,	value : 32'd2147565696,	reg_addr : 32'd279454},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279455},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279456},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279457},
'{step_type : REG_WRITE,	value : 32'd2147566720,	reg_addr : 32'd279458},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279459},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279460},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279461},
'{step_type : REG_WRITE,	value : 32'd67116032,	reg_addr : 32'd279462},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279463},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279464},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279465},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd279466},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279467},
'{step_type : REG_WRITE,	value : 32'd536871046,	reg_addr : 32'd279468},
'{step_type : REG_WRITE,	value : 32'd116676,	reg_addr : 32'd279469},
'{step_type : REG_WRITE,	value : 32'd2650801280,	reg_addr : 32'd279470},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279471},
'{step_type : REG_WRITE,	value : 32'd3288727680,	reg_addr : 32'd279472},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279473},
'{step_type : REG_WRITE,	value : 32'd3556770944,	reg_addr : 32'd279474},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279475},
'{step_type : REG_WRITE,	value : 32'd3825206400,	reg_addr : 32'd279476},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279477},
'{step_type : REG_WRITE,	value : 32'd2617258112,	reg_addr : 32'd279478},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279479},
'{step_type : REG_WRITE,	value : 32'd2080374912,	reg_addr : 32'd279480},
'{step_type : REG_WRITE,	value : 32'd116673,	reg_addr : 32'd279481},
'{step_type : REG_WRITE,	value : 32'd2281704576,	reg_addr : 32'd279482},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279483},
'{step_type : REG_WRITE,	value : 32'd1677724800,	reg_addr : 32'd279484},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279485},
'{step_type : REG_WRITE,	value : 32'd2415921280,	reg_addr : 32'd279486},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279487},
'{step_type : REG_WRITE,	value : 32'd3960470656,	reg_addr : 32'd279488},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279489},
'{step_type : REG_WRITE,	value : 32'd3959423104,	reg_addr : 32'd279490},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279491},
'{step_type : REG_WRITE,	value : 32'd4160749696,	reg_addr : 32'd279492},
'{step_type : REG_WRITE,	value : 32'd2046,	reg_addr : 32'd279493},
'{step_type : REG_WRITE,	value : 32'd4160750720,	reg_addr : 32'd279494},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279495},
'{step_type : REG_WRITE,	value : 32'd4160750720,	reg_addr : 32'd279496},
'{step_type : REG_WRITE,	value : 32'd2002,	reg_addr : 32'd279497},
'{step_type : REG_WRITE,	value : 32'd2818576512,	reg_addr : 32'd279498},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279499},
'{step_type : REG_WRITE,	value : 32'd2147567744,	reg_addr : 32'd279500},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279501},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279502},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279503},
'{step_type : REG_WRITE,	value : 32'd2147568768,	reg_addr : 32'd279504},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279505},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279506},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279507},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd279508},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd279509},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279510},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279511},
'{step_type : REG_WRITE,	value : 32'd4160749696,	reg_addr : 32'd279512},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279513},
'{step_type : REG_WRITE,	value : 32'd4160749696,	reg_addr : 32'd279514},
'{step_type : REG_WRITE,	value : 32'd2002,	reg_addr : 32'd279515},
'{step_type : REG_WRITE,	value : 32'd3960470656,	reg_addr : 32'd279516},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279517},
'{step_type : REG_WRITE,	value : 32'd3959423104,	reg_addr : 32'd279518},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279519},
'{step_type : REG_WRITE,	value : 32'd4160750720,	reg_addr : 32'd279520},
'{step_type : REG_WRITE,	value : 32'd1990,	reg_addr : 32'd279521},
'{step_type : REG_WRITE,	value : 32'd4160750720,	reg_addr : 32'd279522},
'{step_type : REG_WRITE,	value : 32'd2006,	reg_addr : 32'd279523},
'{step_type : REG_WRITE,	value : 32'd2818576512,	reg_addr : 32'd279524},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279525},
'{step_type : REG_WRITE,	value : 32'd2147569792,	reg_addr : 32'd279526},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279527},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279528},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279529},
'{step_type : REG_WRITE,	value : 32'd2147570816,	reg_addr : 32'd279530},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279531},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279532},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279533},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd279534},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd279535},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279536},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279537},
'{step_type : REG_WRITE,	value : 32'd4160749696,	reg_addr : 32'd279538},
'{step_type : REG_WRITE,	value : 32'd1990,	reg_addr : 32'd279539},
'{step_type : REG_WRITE,	value : 32'd4160749696,	reg_addr : 32'd279540},
'{step_type : REG_WRITE,	value : 32'd2006,	reg_addr : 32'd279541},
'{step_type : REG_WRITE,	value : 32'd1677723776,	reg_addr : 32'd279542},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279543},
'{step_type : REG_WRITE,	value : 32'd5152,	reg_addr : 32'd279544},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279545},
'{step_type : REG_WRITE,	value : 32'd3288335488,	reg_addr : 32'd279546},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd279547},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279548},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279549},
'{step_type : REG_WRITE,	value : 32'd3288334464,	reg_addr : 32'd279550},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd279551},
'{step_type : REG_WRITE,	value : 32'd67110400,	reg_addr : 32'd279552},
'{step_type : REG_WRITE,	value : 32'd1024,	reg_addr : 32'd279553},
'{step_type : REG_WRITE,	value : 32'd617138368,	reg_addr : 32'd279554},
'{step_type : REG_WRITE,	value : 32'd83912,	reg_addr : 32'd279555},
'{step_type : REG_WRITE,	value : 32'd2147484800,	reg_addr : 32'd279556},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279557},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279558},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279559},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279560},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279561},
'{step_type : REG_WRITE,	value : 32'd2415919232,	reg_addr : 32'd279562},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279563},
'{step_type : REG_WRITE,	value : 32'd2550140032,	reg_addr : 32'd279564},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279565},
'{step_type : REG_WRITE,	value : 32'd2818576512,	reg_addr : 32'd279566},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279567},
'{step_type : REG_WRITE,	value : 32'd2147571840,	reg_addr : 32'd279568},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279569},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279570},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279571},
'{step_type : REG_WRITE,	value : 32'd2147572864,	reg_addr : 32'd279572},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279573},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279574},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279575},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd279576},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd279577},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279578},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279579},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279580},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279581},
'{step_type : REG_WRITE,	value : 32'd2550136960,	reg_addr : 32'd279582},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279583},
'{step_type : REG_WRITE,	value : 32'd2281701504,	reg_addr : 32'd279584},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279585},
'{step_type : REG_WRITE,	value : 32'd1677721728,	reg_addr : 32'd279586},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279587},
'{step_type : REG_WRITE,	value : 32'd2080375936,	reg_addr : 32'd279588},
'{step_type : REG_WRITE,	value : 32'd116673,	reg_addr : 32'd279589},
'{step_type : REG_WRITE,	value : 32'd3825206400,	reg_addr : 32'd279590},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279591},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279592},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279593},
'{step_type : REG_WRITE,	value : 32'd3825205376,	reg_addr : 32'd279594},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279595},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279596},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279597},
'{step_type : REG_WRITE,	value : 32'd6176,	reg_addr : 32'd279598},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279599},
'{step_type : REG_WRITE,	value : 32'd2415920256,	reg_addr : 32'd279600},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279601},
'{step_type : REG_WRITE,	value : 32'd2818576512,	reg_addr : 32'd279602},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279603},
'{step_type : REG_WRITE,	value : 32'd2147573888,	reg_addr : 32'd279604},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279605},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279606},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279607},
'{step_type : REG_WRITE,	value : 32'd2147574912,	reg_addr : 32'd279608},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279609},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279610},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279611},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd279612},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd279613},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279614},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279615},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279616},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279617},
'{step_type : REG_WRITE,	value : 32'd2147484800,	reg_addr : 32'd279618},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279619},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279620},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279621},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279622},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279623},
'{step_type : REG_WRITE,	value : 32'd2415919232,	reg_addr : 32'd279624},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279625},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279626},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279627},
'{step_type : REG_WRITE,	value : 32'd3825206400,	reg_addr : 32'd279628},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279629},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279630},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279631},
'{step_type : REG_WRITE,	value : 32'd3825205376,	reg_addr : 32'd279632},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279633},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279634},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279635},
'{step_type : REG_WRITE,	value : 32'd2818572416,	reg_addr : 32'd279636},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279637},
'{step_type : REG_WRITE,	value : 32'd1342178432,	reg_addr : 32'd279638},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279639},
'{step_type : REG_WRITE,	value : 32'd536872070,	reg_addr : 32'd279640},
'{step_type : REG_WRITE,	value : 32'd116676,	reg_addr : 32'd279641},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd279642},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279643},
'{step_type : REG_WRITE,	value : 32'd2147517952,	reg_addr : 32'd279644},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279645},
'{step_type : REG_WRITE,	value : 32'd581984,	reg_addr : 32'd279646},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279647},
'{step_type : REG_WRITE,	value : 32'd2147484800,	reg_addr : 32'd279648},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279649},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279650},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279651},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279652},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279653},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279654},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279655},
'{step_type : REG_WRITE,	value : 32'd3825206400,	reg_addr : 32'd279656},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279657},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279658},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279659},
'{step_type : REG_WRITE,	value : 32'd3825205376,	reg_addr : 32'd279660},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279661},
'{step_type : REG_WRITE,	value : 32'd2818572416,	reg_addr : 32'd279662},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279663},
'{step_type : REG_WRITE,	value : 32'd3087007872,	reg_addr : 32'd279664},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279665},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279666},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279667},
'{step_type : REG_WRITE,	value : 32'd4224,	reg_addr : 32'd279668},
'{step_type : REG_WRITE,	value : 32'd13250,	reg_addr : 32'd279669},
'{step_type : REG_WRITE,	value : 32'd1342178432,	reg_addr : 32'd279670},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279671},
'{step_type : REG_WRITE,	value : 32'd3019899008,	reg_addr : 32'd279672},
'{step_type : REG_WRITE,	value : 32'd9216,	reg_addr : 32'd279673},
'{step_type : REG_WRITE,	value : 32'd2281702529,	reg_addr : 32'd279674},
'{step_type : REG_WRITE,	value : 32'd3072,	reg_addr : 32'd279675},
'{step_type : REG_WRITE,	value : 32'd603980928,	reg_addr : 32'd279676},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279677},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd279678},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279679},
'{step_type : REG_WRITE,	value : 32'd1073742976,	reg_addr : 32'd279680},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279681},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd279682},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279683},
'{step_type : REG_WRITE,	value : 32'd2348810368,	reg_addr : 32'd279684},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279685},
'{step_type : REG_WRITE,	value : 32'd2098688,	reg_addr : 32'd279686},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd279687},
'{step_type : REG_WRITE,	value : 32'd2282487936,	reg_addr : 32'd279688},
'{step_type : REG_WRITE,	value : 32'd3074,	reg_addr : 32'd279689},
'{step_type : REG_WRITE,	value : 32'd2282488000,	reg_addr : 32'd279690},
'{step_type : REG_WRITE,	value : 32'd3138,	reg_addr : 32'd279691},
'{step_type : REG_WRITE,	value : 32'd612367488,	reg_addr : 32'd279692},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279693},
'{step_type : REG_WRITE,	value : 32'd673184896,	reg_addr : 32'd279694},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279695},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279696},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279697},
'{step_type : REG_WRITE,	value : 32'd2550137984,	reg_addr : 32'd279698},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279699},
'{step_type : REG_WRITE,	value : 32'd671089792,	reg_addr : 32'd279700},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279701},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279702},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279703},
'{step_type : REG_WRITE,	value : 32'd2164259968,	reg_addr : 32'd279704},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279705},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279706},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279707},
'{step_type : REG_WRITE,	value : 32'd3758097536,	reg_addr : 32'd279708},
'{step_type : REG_WRITE,	value : 32'd2051,	reg_addr : 32'd279709},
'{step_type : REG_WRITE,	value : 32'd67117056,	reg_addr : 32'd279710},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279711},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279712},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279713},
'{step_type : REG_WRITE,	value : 32'd1342177408,	reg_addr : 32'd279714},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279715},
'{step_type : REG_WRITE,	value : 32'd1152,	reg_addr : 32'd279716},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279717},
'{step_type : REG_WRITE,	value : 32'd201326720,	reg_addr : 32'd279718},
'{step_type : REG_WRITE,	value : 32'd6144,	reg_addr : 32'd279719},
'{step_type : REG_WRITE,	value : 32'd1543504000,	reg_addr : 32'd279720},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279721},
'{step_type : REG_WRITE,	value : 32'd67108992,	reg_addr : 32'd279722},
'{step_type : REG_WRITE,	value : 32'd11264,	reg_addr : 32'd279723},
'{step_type : REG_WRITE,	value : 32'd33555968,	reg_addr : 32'd279724},
'{step_type : REG_WRITE,	value : 32'd512,	reg_addr : 32'd279725},
'{step_type : REG_WRITE,	value : 32'd738201792,	reg_addr : 32'd279726},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279727},
'{step_type : REG_WRITE,	value : 32'd738203776,	reg_addr : 32'd279728},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279729},
'{step_type : REG_WRITE,	value : 32'd402659456,	reg_addr : 32'd279730},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279731},
'{step_type : REG_WRITE,	value : 32'd469768320,	reg_addr : 32'd279732},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279733},
'{step_type : REG_WRITE,	value : 32'd536877184,	reg_addr : 32'd279734},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279735},
'{step_type : REG_WRITE,	value : 32'd603986048,	reg_addr : 32'd279736},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279737},
'{step_type : REG_WRITE,	value : 32'd671094912,	reg_addr : 32'd279738},
'{step_type : REG_WRITE,	value : 32'd15297,	reg_addr : 32'd279739},
'{step_type : REG_WRITE,	value : 32'd536873088,	reg_addr : 32'd279740},
'{step_type : REG_WRITE,	value : 32'd11212,	reg_addr : 32'd279741},
'{step_type : REG_WRITE,	value : 32'd67121312,	reg_addr : 32'd279742},
'{step_type : REG_WRITE,	value : 32'd11264,	reg_addr : 32'd279743},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279744},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279745},
'{step_type : REG_WRITE,	value : 32'd3019900032,	reg_addr : 32'd279746},
'{step_type : REG_WRITE,	value : 32'd9216,	reg_addr : 32'd279747},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd279748},
'{step_type : REG_WRITE,	value : 32'd16384,	reg_addr : 32'd279749},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd279750},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279751},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd279752},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279753},
'{step_type : REG_WRITE,	value : 32'd2281704576,	reg_addr : 32'd279754},
'{step_type : REG_WRITE,	value : 32'd3072,	reg_addr : 32'd279755},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279756},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279757},
'{step_type : REG_WRITE,	value : 32'd67111936,	reg_addr : 32'd279758},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279759},
'{step_type : REG_WRITE,	value : 32'd2281702528,	reg_addr : 32'd279760},
'{step_type : REG_WRITE,	value : 32'd2050,	reg_addr : 32'd279761},
'{step_type : REG_WRITE,	value : 32'd480,	reg_addr : 32'd279762},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279763},
'{step_type : REG_WRITE,	value : 32'd6272,	reg_addr : 32'd279764},
'{step_type : REG_WRITE,	value : 32'd13250,	reg_addr : 32'd279765},
'{step_type : REG_WRITE,	value : 32'd2497,	reg_addr : 32'd279766},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279767},
'{step_type : REG_WRITE,	value : 32'd2617249041,	reg_addr : 32'd279768},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279769},
'{step_type : REG_WRITE,	value : 32'd67112977,	reg_addr : 32'd279770},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279771},
'{step_type : REG_WRITE,	value : 32'd2617250065,	reg_addr : 32'd279772},
'{step_type : REG_WRITE,	value : 32'd7171,	reg_addr : 32'd279773},
'{step_type : REG_WRITE,	value : 32'd67112977,	reg_addr : 32'd279774},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279775},
'{step_type : REG_WRITE,	value : 32'd2617245841,	reg_addr : 32'd279776},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279777},
'{step_type : REG_WRITE,	value : 32'd2617245841,	reg_addr : 32'd279778},
'{step_type : REG_WRITE,	value : 32'd7171,	reg_addr : 32'd279779},
'{step_type : REG_WRITE,	value : 32'd649505,	reg_addr : 32'd279780},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279781},
'{step_type : REG_WRITE,	value : 32'd3087008896,	reg_addr : 32'd279782},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279783},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279784},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279785},
'{step_type : REG_WRITE,	value : 32'd2147910144,	reg_addr : 32'd279786},
'{step_type : REG_WRITE,	value : 32'd16399,	reg_addr : 32'd279787},
'{step_type : REG_WRITE,	value : 32'd647488,	reg_addr : 32'd279788},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279789},
'{step_type : REG_WRITE,	value : 32'd36288,	reg_addr : 32'd279790},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279791},
'{step_type : REG_WRITE,	value : 32'd97728,	reg_addr : 32'd279792},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279793},
'{step_type : REG_WRITE,	value : 32'd172480,	reg_addr : 32'd279794},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279795},
'{step_type : REG_WRITE,	value : 32'd224704,	reg_addr : 32'd279796},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279797},
'{step_type : REG_WRITE,	value : 32'd234944,	reg_addr : 32'd279798},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279799},
'{step_type : REG_WRITE,	value : 32'd241088,	reg_addr : 32'd279800},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279801},
'{step_type : REG_WRITE,	value : 32'd375232,	reg_addr : 32'd279802},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279803},
'{step_type : REG_WRITE,	value : 32'd1610727552,	reg_addr : 32'd279804},
'{step_type : REG_WRITE,	value : 32'd9253,	reg_addr : 32'd279805},
'{step_type : REG_WRITE,	value : 32'd524800,	reg_addr : 32'd279806},
'{step_type : REG_WRITE,	value : 32'd16398,	reg_addr : 32'd279807},
'{step_type : REG_WRITE,	value : 32'd665920,	reg_addr : 32'd279808},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279809},
'{step_type : REG_WRITE,	value : 32'd658737,	reg_addr : 32'd279810},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279811},
'{step_type : REG_WRITE,	value : 32'd457152,	reg_addr : 32'd279812},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279813},
'{step_type : REG_WRITE,	value : 32'd2147517952,	reg_addr : 32'd279814},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279815},
'{step_type : REG_WRITE,	value : 32'd665920,	reg_addr : 32'd279816},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279817},
'{step_type : REG_WRITE,	value : 32'd481730,	reg_addr : 32'd279818},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279819},
'{step_type : REG_WRITE,	value : 32'd2147910144,	reg_addr : 32'd279820},
'{step_type : REG_WRITE,	value : 32'd16399,	reg_addr : 32'd279821},
'{step_type : REG_WRITE,	value : 32'd3288335552,	reg_addr : 32'd279822},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd279823},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279824},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279825},
'{step_type : REG_WRITE,	value : 32'd3288334528,	reg_addr : 32'd279826},
'{step_type : REG_WRITE,	value : 32'd1984,	reg_addr : 32'd279827},
'{step_type : REG_WRITE,	value : 32'd1073767953,	reg_addr : 32'd279828},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279829},
'{step_type : REG_WRITE,	value : 32'd684369,	reg_addr : 32'd279830},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279831},
'{step_type : REG_WRITE,	value : 32'd2147910161,	reg_addr : 32'd279832},
'{step_type : REG_WRITE,	value : 32'd16399,	reg_addr : 32'd279833},
'{step_type : REG_WRITE,	value : 32'd684369,	reg_addr : 32'd279834},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279835},
'{step_type : REG_WRITE,	value : 32'd524817,	reg_addr : 32'd279836},
'{step_type : REG_WRITE,	value : 32'd16398,	reg_addr : 32'd279837},
'{step_type : REG_WRITE,	value : 32'd674129,	reg_addr : 32'd279838},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279839},
'{step_type : REG_WRITE,	value : 32'd2147517969,	reg_addr : 32'd279840},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279841},
'{step_type : REG_WRITE,	value : 32'd677233,	reg_addr : 32'd279842},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279843},
'{step_type : REG_WRITE,	value : 32'd4145,	reg_addr : 32'd279844},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279845},
'{step_type : REG_WRITE,	value : 32'd4145,	reg_addr : 32'd279846},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279847},
'{step_type : REG_WRITE,	value : 32'd11313,	reg_addr : 32'd279848},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279849},
'{step_type : REG_WRITE,	value : 32'd2818572433,	reg_addr : 32'd279850},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279851},
'{step_type : REG_WRITE,	value : 32'd2147575953,	reg_addr : 32'd279852},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279853},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279854},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279855},
'{step_type : REG_WRITE,	value : 32'd2147576977,	reg_addr : 32'd279856},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279857},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279858},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279859},
'{step_type : REG_WRITE,	value : 32'd2129,	reg_addr : 32'd279860},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd279861},
'{step_type : REG_WRITE,	value : 32'd2147483793,	reg_addr : 32'd279862},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279863},
'{step_type : REG_WRITE,	value : 32'd603979921,	reg_addr : 32'd279864},
'{step_type : REG_WRITE,	value : 32'd123936,	reg_addr : 32'd279865},
'{step_type : REG_WRITE,	value : 32'd571840,	reg_addr : 32'd279866},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279867},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279868},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279869},
'{step_type : REG_WRITE,	value : 32'd590272,	reg_addr : 32'd279870},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279871},
'{step_type : REG_WRITE,	value : 32'd603980928,	reg_addr : 32'd279872},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279873},
'{step_type : REG_WRITE,	value : 32'd1024,	reg_addr : 32'd279874},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279875},
'{step_type : REG_WRITE,	value : 32'd1342177408,	reg_addr : 32'd279876},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279877},
'{step_type : REG_WRITE,	value : 32'd2617249024,	reg_addr : 32'd279878},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279879},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279880},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279881},
'{step_type : REG_WRITE,	value : 32'd2617250048,	reg_addr : 32'd279882},
'{step_type : REG_WRITE,	value : 32'd7171,	reg_addr : 32'd279883},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279884},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279885},
'{step_type : REG_WRITE,	value : 32'd2617245824,	reg_addr : 32'd279886},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279887},
'{step_type : REG_WRITE,	value : 32'd2617245824,	reg_addr : 32'd279888},
'{step_type : REG_WRITE,	value : 32'd7171,	reg_addr : 32'd279889},
'{step_type : REG_WRITE,	value : 32'd6272,	reg_addr : 32'd279890},
'{step_type : REG_WRITE,	value : 32'd13250,	reg_addr : 32'd279891},
'{step_type : REG_WRITE,	value : 32'd3087008896,	reg_addr : 32'd279892},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd279893},
'{step_type : REG_WRITE,	value : 32'd67111936,	reg_addr : 32'd279894},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279895},
'{step_type : REG_WRITE,	value : 32'd603980945,	reg_addr : 32'd279896},
'{step_type : REG_WRITE,	value : 32'd123936,	reg_addr : 32'd279897},
'{step_type : REG_WRITE,	value : 32'd2818572416,	reg_addr : 32'd279898},
'{step_type : REG_WRITE,	value : 32'd7174,	reg_addr : 32'd279899},
'{step_type : REG_WRITE,	value : 32'd2147559552,	reg_addr : 32'd279900},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279901},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279902},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279903},
'{step_type : REG_WRITE,	value : 32'd2147560576,	reg_addr : 32'd279904},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279905},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279906},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279907},
'{step_type : REG_WRITE,	value : 32'd2112,	reg_addr : 32'd279908},
'{step_type : REG_WRITE,	value : 32'd24576,	reg_addr : 32'd279909},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279910},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd279911},
'{step_type : REG_WRITE,	value : 32'd738197632,	reg_addr : 32'd279912},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279913},
'{step_type : REG_WRITE,	value : 32'd2350907520,	reg_addr : 32'd279914},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279915},
'{step_type : REG_WRITE,	value : 32'd2098688,	reg_addr : 32'd279916},
'{step_type : REG_WRITE,	value : 32'd32,	reg_addr : 32'd279917},
'{step_type : REG_WRITE,	value : 32'd2285633664,	reg_addr : 32'd279918},
'{step_type : REG_WRITE,	value : 32'd3074,	reg_addr : 32'd279919},
'{step_type : REG_WRITE,	value : 32'd2285633728,	reg_addr : 32'd279920},
'{step_type : REG_WRITE,	value : 32'd3138,	reg_addr : 32'd279921},
'{step_type : REG_WRITE,	value : 32'd2550137984,	reg_addr : 32'd279922},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279923},
'{step_type : REG_WRITE,	value : 32'd671089792,	reg_addr : 32'd279924},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279925},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279926},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279927},
'{step_type : REG_WRITE,	value : 32'd2164259968,	reg_addr : 32'd279928},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279929},
'{step_type : REG_WRITE,	value : 32'd612367488,	reg_addr : 32'd279930},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279931},
'{step_type : REG_WRITE,	value : 32'd673184896,	reg_addr : 32'd279932},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279933},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd279934},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279935},
'{step_type : REG_WRITE,	value : 32'd3758097536,	reg_addr : 32'd279936},
'{step_type : REG_WRITE,	value : 32'd2051,	reg_addr : 32'd279937},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279938},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279939},
'{step_type : REG_WRITE,	value : 32'd8390144,	reg_addr : 32'd279940},
'{step_type : REG_WRITE,	value : 32'd128,	reg_addr : 32'd279941},
'{step_type : REG_WRITE,	value : 32'd67109056,	reg_addr : 32'd279942},
'{step_type : REG_WRITE,	value : 32'd9252,	reg_addr : 32'd279943},
'{step_type : REG_WRITE,	value : 32'd67141856,	reg_addr : 32'd279944},
'{step_type : REG_WRITE,	value : 32'd9252,	reg_addr : 32'd279945},
'{step_type : REG_WRITE,	value : 32'd1073743074,	reg_addr : 32'd279946},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279947},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279948},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279949},
'{step_type : REG_WRITE,	value : 32'd1073742050,	reg_addr : 32'd279950},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279951},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279952},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279953},
'{step_type : REG_WRITE,	value : 32'd2147484896,	reg_addr : 32'd279954},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279955},
'{step_type : REG_WRITE,	value : 32'd2147483872,	reg_addr : 32'd279956},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279957},
'{step_type : REG_WRITE,	value : 32'd1541,	reg_addr : 32'd279958},
'{step_type : REG_WRITE,	value : 32'd8192,	reg_addr : 32'd279959},
'{step_type : REG_WRITE,	value : 32'd1073743042,	reg_addr : 32'd279960},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279961},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279962},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279963},
'{step_type : REG_WRITE,	value : 32'd1073742018,	reg_addr : 32'd279964},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279965},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279966},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279967},
'{step_type : REG_WRITE,	value : 32'd2147484864,	reg_addr : 32'd279968},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279969},
'{step_type : REG_WRITE,	value : 32'd2147483840,	reg_addr : 32'd279970},
'{step_type : REG_WRITE,	value : 32'd11276,	reg_addr : 32'd279971},
'{step_type : REG_WRITE,	value : 32'd67111936,	reg_addr : 32'd279972},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279973},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279974},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd279975},
'{step_type : REG_WRITE,	value : 32'd268435968,	reg_addr : 32'd279976},
'{step_type : REG_WRITE,	value : 32'd20480,	reg_addr : 32'd279977},
'{step_type : REG_WRITE,	value : 32'd744768,	reg_addr : 32'd279978},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279979},
'{step_type : REG_WRITE,	value : 32'd64,	reg_addr : 32'd279980},
'{step_type : REG_WRITE,	value : 32'd16384,	reg_addr : 32'd279981},
'{step_type : REG_WRITE,	value : 32'd671089792,	reg_addr : 32'd279982},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279983},
'{step_type : REG_WRITE,	value : 32'd67112960,	reg_addr : 32'd279984},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279985},
'{step_type : REG_WRITE,	value : 32'd3758096512,	reg_addr : 32'd279986},
'{step_type : REG_WRITE,	value : 32'd2051,	reg_addr : 32'd279987},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd279988},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd279989},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279990},
'{step_type : REG_WRITE,	value : 32'd4032,	reg_addr : 32'd279991},
'{step_type : REG_WRITE,	value : 32'd2147483776,	reg_addr : 32'd279992},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279993},
'{step_type : REG_WRITE,	value : 32'd2550136960,	reg_addr : 32'd279994},
'{step_type : REG_WRITE,	value : 32'd4034,	reg_addr : 32'd279995},
'{step_type : REG_WRITE,	value : 32'd603979904,	reg_addr : 32'd279996},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279997},
'{step_type : REG_WRITE,	value : 32'd671088768,	reg_addr : 32'd279998},
'{step_type : REG_WRITE,	value : 32'd1986,	reg_addr : 32'd279999},
'{step_type : REG_WRITE,	value : 32'd3825206400,	reg_addr : 32'd280000},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd280001},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd280002},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280003},
'{step_type : REG_WRITE,	value : 32'd3825205376,	reg_addr : 32'd280004},
'{step_type : REG_WRITE,	value : 32'd2049,	reg_addr : 32'd280005},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd280006},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280007},
'{step_type : REG_WRITE,	value : 32'd2818573440,	reg_addr : 32'd280008},
'{step_type : REG_WRITE,	value : 32'd7172,	reg_addr : 32'd280009},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd280010},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280011},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd280012},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280013},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd280014},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280015},
'{step_type : REG_WRITE,	value : 32'd4128,	reg_addr : 32'd280016},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280017},
'{step_type : REG_WRITE,	value : 32'd3892513920,	reg_addr : 32'd280018},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd280019},
'{step_type : REG_WRITE,	value : 32'd67110912,	reg_addr : 32'd280020},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280021},
'{step_type : REG_WRITE,	value : 32'd3892314240,	reg_addr : 32'd280022},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd280023},
'{step_type : REG_WRITE,	value : 32'd67109888,	reg_addr : 32'd280024},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280025},
'{step_type : REG_WRITE,	value : 32'd2617248928,	reg_addr : 32'd280026},
'{step_type : REG_WRITE,	value : 32'd7169,	reg_addr : 32'd280027},
'{step_type : REG_WRITE,	value : 32'd2617249952,	reg_addr : 32'd280028},
'{step_type : REG_WRITE,	value : 32'd7171,	reg_addr : 32'd280029},
'{step_type : REG_WRITE,	value : 32'd658720,	reg_addr : 32'd280030},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd280031},
'{step_type : REG_WRITE,	value : 32'd1536,	reg_addr : 32'd852199},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459146},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd459556},
'{step_type : REG_WRITE,	value : 32'd25,	reg_addr : 32'd459557},
'{step_type : REG_WRITE,	value : 32'd46,	reg_addr : 32'd459558},
'{step_type : REG_WRITE,	value : 32'd67,	reg_addr : 32'd459559},
'{step_type : REG_WRITE,	value : 32'd91,	reg_addr : 32'd459560},
'{step_type : REG_WRITE,	value : 32'd112,	reg_addr : 32'd459561},
'{step_type : REG_WRITE,	value : 32'd133,	reg_addr : 32'd459562},
'{step_type : REG_WRITE,	value : 32'd157,	reg_addr : 32'd459563},
'{step_type : REG_WRITE,	value : 32'd178,	reg_addr : 32'd459564},
'{step_type : REG_WRITE,	value : 32'd199,	reg_addr : 32'd459565},
'{step_type : REG_WRITE,	value : 32'd223,	reg_addr : 32'd459566},
'{step_type : REG_WRITE,	value : 32'd244,	reg_addr : 32'd459567},
'{step_type : REG_WRITE,	value : 32'd265,	reg_addr : 32'd459568},
'{step_type : REG_WRITE,	value : 32'd275,	reg_addr : 32'd459569},
'{step_type : REG_WRITE,	value : 32'd277,	reg_addr : 32'd459570},
'{step_type : REG_WRITE,	value : 32'd281,	reg_addr : 32'd459571},
'{step_type : REG_WRITE,	value : 32'd283,	reg_addr : 32'd459572},
'{step_type : REG_WRITE,	value : 32'd287,	reg_addr : 32'd459573},
'{step_type : REG_WRITE,	value : 32'd289,	reg_addr : 32'd459574},
'{step_type : REG_WRITE,	value : 32'd290,	reg_addr : 32'd459575},
'{step_type : REG_WRITE,	value : 32'd291,	reg_addr : 32'd459577},
'{step_type : REG_WRITE,	value : 32'd293,	reg_addr : 32'd459578},
'{step_type : REG_WRITE,	value : 32'd295,	reg_addr : 32'd459579},
'{step_type : REG_WRITE,	value : 32'd296,	reg_addr : 32'd459580},
'{step_type : REG_WRITE,	value : 32'd321,	reg_addr : 32'd459581},
'{step_type : REG_WRITE,	value : 32'd331,	reg_addr : 32'd459582},
'{step_type : REG_WRITE,	value : 32'd355,	reg_addr : 32'd459583},
'{step_type : REG_WRITE,	value : 32'd371,	reg_addr : 32'd459600},
'{step_type : REG_WRITE,	value : 32'd395,	reg_addr : 32'd459601},
'{step_type : REG_WRITE,	value : 32'd404,	reg_addr : 32'd459602},
'{step_type : REG_WRITE,	value : 32'd422,	reg_addr : 32'd459603},
'{step_type : REG_WRITE,	value : 32'd24,	reg_addr : 32'd459659},
'{step_type : REG_WRITE,	value : 32'd45,	reg_addr : 32'd459660},
'{step_type : REG_WRITE,	value : 32'd66,	reg_addr : 32'd459661},
'{step_type : REG_WRITE,	value : 32'd90,	reg_addr : 32'd459662},
'{step_type : REG_WRITE,	value : 32'd111,	reg_addr : 32'd459663},
'{step_type : REG_WRITE,	value : 32'd132,	reg_addr : 32'd459664},
'{step_type : REG_WRITE,	value : 32'd156,	reg_addr : 32'd459665},
'{step_type : REG_WRITE,	value : 32'd177,	reg_addr : 32'd459666},
'{step_type : REG_WRITE,	value : 32'd198,	reg_addr : 32'd459667},
'{step_type : REG_WRITE,	value : 32'd222,	reg_addr : 32'd459668},
'{step_type : REG_WRITE,	value : 32'd243,	reg_addr : 32'd459669},
'{step_type : REG_WRITE,	value : 32'd264,	reg_addr : 32'd459670},
'{step_type : REG_WRITE,	value : 32'd274,	reg_addr : 32'd459671},
'{step_type : REG_WRITE,	value : 32'd276,	reg_addr : 32'd459672},
'{step_type : REG_WRITE,	value : 32'd280,	reg_addr : 32'd459673},
'{step_type : REG_WRITE,	value : 32'd282,	reg_addr : 32'd459674},
'{step_type : REG_WRITE,	value : 32'd286,	reg_addr : 32'd459675},
'{step_type : REG_WRITE,	value : 32'd288,	reg_addr : 32'd459676},
'{step_type : REG_WRITE,	value : 32'd289,	reg_addr : 32'd459677},
'{step_type : REG_WRITE,	value : 32'd290,	reg_addr : 32'd459678},
'{step_type : REG_WRITE,	value : 32'd292,	reg_addr : 32'd459680},
'{step_type : REG_WRITE,	value : 32'd294,	reg_addr : 32'd459681},
'{step_type : REG_WRITE,	value : 32'd295,	reg_addr : 32'd459682},
'{step_type : REG_WRITE,	value : 32'd320,	reg_addr : 32'd459683},
'{step_type : REG_WRITE,	value : 32'd330,	reg_addr : 32'd459684},
'{step_type : REG_WRITE,	value : 32'd354,	reg_addr : 32'd459685},
'{step_type : REG_WRITE,	value : 32'd370,	reg_addr : 32'd459686},
'{step_type : REG_WRITE,	value : 32'd394,	reg_addr : 32'd459703},
'{step_type : REG_WRITE,	value : 32'd403,	reg_addr : 32'd459704},
'{step_type : REG_WRITE,	value : 32'd421,	reg_addr : 32'd459705},
'{step_type : REG_WRITE,	value : 32'd438,	reg_addr : 32'd459706},
'{step_type : REG_WRITE,	value : 32'd1038,	reg_addr : 32'd459264},
'{step_type : REG_WRITE,	value : 32'd1103,	reg_addr : 32'd459266},
'{step_type : REG_WRITE,	value : 32'd192,	reg_addr : 32'd459268},
'{step_type : REG_WRITE,	value : 32'd582,	reg_addr : 32'd459269},
'{step_type : REG_WRITE,	value : 32'd257,	reg_addr : 32'd459270},
'{step_type : REG_WRITE,	value : 32'd647,	reg_addr : 32'd459271},
'{step_type : REG_WRITE,	value : 32'd322,	reg_addr : 32'd459272},
'{step_type : REG_WRITE,	value : 32'd712,	reg_addr : 32'd459273},
'{step_type : REG_WRITE,	value : 32'd18,	reg_addr : 32'd459274},
'{step_type : REG_WRITE,	value : 32'd844,	reg_addr : 32'd459275},
'{step_type : REG_WRITE,	value : 32'd21,	reg_addr : 32'd459276},
'{step_type : REG_WRITE,	value : 32'd22,	reg_addr : 32'd459278},
'{step_type : REG_WRITE,	value : 32'd23,	reg_addr : 32'd459280},
'{step_type : REG_WRITE,	value : 32'd44,	reg_addr : 32'd459282},
'{step_type : REG_WRITE,	value : 32'd24,	reg_addr : 32'd459283},
'{step_type : REG_WRITE,	value : 32'd45,	reg_addr : 32'd459284},
'{step_type : REG_WRITE,	value : 32'd25,	reg_addr : 32'd459285},
'{step_type : REG_WRITE,	value : 32'd46,	reg_addr : 32'd459286},
'{step_type : REG_WRITE,	value : 32'd26,	reg_addr : 32'd459287},
'{step_type : REG_WRITE,	value : 32'd47,	reg_addr : 32'd459288},
'{step_type : REG_WRITE,	value : 32'd27,	reg_addr : 32'd459289},
'{step_type : REG_WRITE,	value : 32'd19,	reg_addr : 32'd459290},
'{step_type : REG_WRITE,	value : 32'd618,	reg_addr : 32'd589852},
'{step_type : REG_WRITE,	value : 32'd618,	reg_addr : 32'd589853},
'{step_type : REG_WRITE,	value : 32'd618,	reg_addr : 32'd589854},
'{step_type : REG_WRITE,	value : 32'd618,	reg_addr : 32'd589855},
'{step_type : REG_WRITE,	value : 32'd674,	reg_addr : 32'd589856},
'{step_type : REG_WRITE,	value : 32'd618,	reg_addr : 32'd589857},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd589858},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd589859},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd589860},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd589861},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd589862},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd589863},
'{step_type : REG_WRITE,	value : 32'd671,	reg_addr : 32'd589867},
'{step_type : REG_WRITE,	value : 32'd2,	reg_addr : 32'd459077},
'{step_type : REG_WRITE,	value : 32'd51672,	reg_addr : 32'd266244},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266245},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266246},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266247},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266248},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266249},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266250},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266251},
'{step_type : REG_WRITE,	value : 32'd51544,	reg_addr : 32'd266252},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266253},
'{step_type : REG_WRITE,	value : 32'd53000,	reg_addr : 32'd266254},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266255},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266256},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266257},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266258},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266259},
'{step_type : REG_WRITE,	value : 32'd49368,	reg_addr : 32'd266260},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266261},
'{step_type : REG_WRITE,	value : 32'd55368,	reg_addr : 32'd266262},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266263},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266264},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266265},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266266},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266267},
'{step_type : REG_WRITE,	value : 32'd49496,	reg_addr : 32'd266268},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266269},
'{step_type : REG_WRITE,	value : 32'd56776,	reg_addr : 32'd266270},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266271},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266272},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266273},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266274},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266275},
'{step_type : REG_WRITE,	value : 32'd49624,	reg_addr : 32'd266276},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266277},
'{step_type : REG_WRITE,	value : 32'd49928,	reg_addr : 32'd266278},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266279},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266280},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266281},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266282},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266283},
'{step_type : REG_WRITE,	value : 32'd50520,	reg_addr : 32'd266284},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266285},
'{step_type : REG_WRITE,	value : 32'd60424,	reg_addr : 32'd266286},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266287},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266288},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266289},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266290},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266291},
'{step_type : REG_WRITE,	value : 32'd50648,	reg_addr : 32'd266292},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266293},
'{step_type : REG_WRITE,	value : 32'd55944,	reg_addr : 32'd266294},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266295},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266296},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266297},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266298},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266299},
'{step_type : REG_WRITE,	value : 32'd18648,	reg_addr : 32'd266300},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266301},
'{step_type : REG_WRITE,	value : 32'd23816,	reg_addr : 32'd266302},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266303},
'{step_type : REG_WRITE,	value : 32'd35032,	reg_addr : 32'd266304},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266305},
'{step_type : REG_WRITE,	value : 32'd40200,	reg_addr : 32'd266306},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266307},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266308},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266309},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266310},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266311},
'{step_type : REG_WRITE,	value : 32'd51800,	reg_addr : 32'd266312},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266313},
'{step_type : REG_WRITE,	value : 32'd49416,	reg_addr : 32'd266314},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266315},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266316},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266317},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266318},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266319},
'{step_type : REG_WRITE,	value : 32'd52056,	reg_addr : 32'd266320},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266321},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266322},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266323},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266324},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266325},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266326},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266327},
'{step_type : REG_WRITE,	value : 32'd54488,	reg_addr : 32'd266328},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266329},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266330},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266331},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266332},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266333},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266334},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266335},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266336},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266337},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266338},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266339},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266340},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266341},
'{step_type : REG_WRITE,	value : 32'd22408,	reg_addr : 32'd266342},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266343},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266344},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266345},
'{step_type : REG_WRITE,	value : 32'd38792,	reg_addr : 32'd266346},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266347},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266348},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266349},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266350},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266351},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266352},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266353},
'{step_type : REG_WRITE,	value : 32'd22472,	reg_addr : 32'd266354},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266355},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266356},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266357},
'{step_type : REG_WRITE,	value : 32'd38792,	reg_addr : 32'd266358},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266359},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266360},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266361},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266362},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266363},
'{step_type : REG_WRITE,	value : 32'd18264,	reg_addr : 32'd266364},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266365},
'{step_type : REG_WRITE,	value : 32'd18824,	reg_addr : 32'd266366},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266367},
'{step_type : REG_WRITE,	value : 32'd34648,	reg_addr : 32'd266368},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266369},
'{step_type : REG_WRITE,	value : 32'd35208,	reg_addr : 32'd266370},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266371},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266372},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266373},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266374},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266375},
'{step_type : REG_WRITE,	value : 32'd18392,	reg_addr : 32'd266376},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266377},
'{step_type : REG_WRITE,	value : 32'd26376,	reg_addr : 32'd266378},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266379},
'{step_type : REG_WRITE,	value : 32'd34776,	reg_addr : 32'd266380},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266381},
'{step_type : REG_WRITE,	value : 32'd42760,	reg_addr : 32'd266382},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266383},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266384},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266385},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266386},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266387},
'{step_type : REG_WRITE,	value : 32'd19544,	reg_addr : 32'd266388},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266389},
'{step_type : REG_WRITE,	value : 32'd18760,	reg_addr : 32'd266390},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266391},
'{step_type : REG_WRITE,	value : 32'd35928,	reg_addr : 32'd266392},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266393},
'{step_type : REG_WRITE,	value : 32'd35144,	reg_addr : 32'd266394},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266395},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266396},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266397},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266398},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266399},
'{step_type : REG_WRITE,	value : 32'd20312,	reg_addr : 32'd266400},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266401},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd266402},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266403},
'{step_type : REG_WRITE,	value : 32'd36696,	reg_addr : 32'd266404},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266405},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd266406},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266407},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266408},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266409},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266410},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266411},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266412},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266413},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266414},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266415},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266416},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266417},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266418},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266419},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266420},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266421},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266422},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266423},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266424},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266425},
'{step_type : REG_WRITE,	value : 32'd22408,	reg_addr : 32'd266426},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266427},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266428},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266429},
'{step_type : REG_WRITE,	value : 32'd38792,	reg_addr : 32'd266430},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266431},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266432},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266433},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266434},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266435},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266436},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266437},
'{step_type : REG_WRITE,	value : 32'd22408,	reg_addr : 32'd266438},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266439},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266440},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266441},
'{step_type : REG_WRITE,	value : 32'd38792,	reg_addr : 32'd266442},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266443},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266444},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266445},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266446},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266447},
'{step_type : REG_WRITE,	value : 32'd18264,	reg_addr : 32'd266448},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266449},
'{step_type : REG_WRITE,	value : 32'd18824,	reg_addr : 32'd266450},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266451},
'{step_type : REG_WRITE,	value : 32'd34648,	reg_addr : 32'd266452},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266453},
'{step_type : REG_WRITE,	value : 32'd35208,	reg_addr : 32'd266454},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266455},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266456},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266457},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266458},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266459},
'{step_type : REG_WRITE,	value : 32'd18392,	reg_addr : 32'd266460},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266461},
'{step_type : REG_WRITE,	value : 32'd26376,	reg_addr : 32'd266462},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266463},
'{step_type : REG_WRITE,	value : 32'd34776,	reg_addr : 32'd266464},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266465},
'{step_type : REG_WRITE,	value : 32'd42760,	reg_addr : 32'd266466},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266467},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266468},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266469},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266470},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266471},
'{step_type : REG_WRITE,	value : 32'd19544,	reg_addr : 32'd266472},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266473},
'{step_type : REG_WRITE,	value : 32'd18760,	reg_addr : 32'd266474},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266475},
'{step_type : REG_WRITE,	value : 32'd35928,	reg_addr : 32'd266476},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266477},
'{step_type : REG_WRITE,	value : 32'd35144,	reg_addr : 32'd266478},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266479},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266480},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266481},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266482},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266483},
'{step_type : REG_WRITE,	value : 32'd20312,	reg_addr : 32'd266484},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266485},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd266486},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266487},
'{step_type : REG_WRITE,	value : 32'd36696,	reg_addr : 32'd266488},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266489},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd266490},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266491},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266492},
'{step_type : REG_WRITE,	value : 32'd1258291200,	reg_addr : 32'd266493},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266494},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266495},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266496},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266497},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266498},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266499},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266500},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266501},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266502},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266503},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266504},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266505},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266506},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266507},
'{step_type : REG_WRITE,	value : 32'd51672,	reg_addr : 32'd266508},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266509},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266510},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266511},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266512},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266513},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266514},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266515},
'{step_type : REG_WRITE,	value : 32'd51544,	reg_addr : 32'd266516},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266517},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266518},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266519},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266520},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266521},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266522},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266523},
'{step_type : REG_WRITE,	value : 32'd49368,	reg_addr : 32'd266524},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266525},
'{step_type : REG_WRITE,	value : 32'd59400,	reg_addr : 32'd266526},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266527},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266528},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266529},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266530},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266531},
'{step_type : REG_WRITE,	value : 32'd49496,	reg_addr : 32'd266532},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266533},
'{step_type : REG_WRITE,	value : 32'd60040,	reg_addr : 32'd266534},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266535},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266536},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266537},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266538},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266539},
'{step_type : REG_WRITE,	value : 32'd49624,	reg_addr : 32'd266540},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266541},
'{step_type : REG_WRITE,	value : 32'd50952,	reg_addr : 32'd266542},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266543},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266544},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266545},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266546},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266547},
'{step_type : REG_WRITE,	value : 32'd50520,	reg_addr : 32'd266548},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266549},
'{step_type : REG_WRITE,	value : 32'd59912,	reg_addr : 32'd266550},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266551},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266552},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266553},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266554},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266555},
'{step_type : REG_WRITE,	value : 32'd50648,	reg_addr : 32'd266556},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266557},
'{step_type : REG_WRITE,	value : 32'd57864,	reg_addr : 32'd266558},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266559},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266560},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266561},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266562},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266563},
'{step_type : REG_WRITE,	value : 32'd18648,	reg_addr : 32'd266564},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266565},
'{step_type : REG_WRITE,	value : 32'd16968,	reg_addr : 32'd266566},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266567},
'{step_type : REG_WRITE,	value : 32'd35032,	reg_addr : 32'd266568},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266569},
'{step_type : REG_WRITE,	value : 32'd38472,	reg_addr : 32'd266570},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266571},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266572},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266573},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266574},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266575},
'{step_type : REG_WRITE,	value : 32'd51800,	reg_addr : 32'd266576},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266577},
'{step_type : REG_WRITE,	value : 32'd49416,	reg_addr : 32'd266578},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266579},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266580},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266581},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266582},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266583},
'{step_type : REG_WRITE,	value : 32'd52056,	reg_addr : 32'd266584},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266585},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266586},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266587},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266588},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266589},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266590},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266591},
'{step_type : REG_WRITE,	value : 32'd54488,	reg_addr : 32'd266592},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266593},
'{step_type : REG_WRITE,	value : 32'd61448,	reg_addr : 32'd266594},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266595},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266596},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266597},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266598},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266599},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266600},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266601},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266602},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266603},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266604},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266605},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266606},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266607},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266608},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266609},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266610},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266611},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266612},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266613},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266614},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266615},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266616},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266617},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266618},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266619},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266620},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266621},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266622},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266623},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266624},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266625},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266626},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266627},
'{step_type : REG_WRITE,	value : 32'd18264,	reg_addr : 32'd266628},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266629},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266630},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266631},
'{step_type : REG_WRITE,	value : 32'd34648,	reg_addr : 32'd266632},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266633},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266634},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266635},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266636},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266637},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266638},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266639},
'{step_type : REG_WRITE,	value : 32'd18392,	reg_addr : 32'd266640},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266641},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266642},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266643},
'{step_type : REG_WRITE,	value : 32'd34776,	reg_addr : 32'd266644},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266645},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266646},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266647},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266648},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266649},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266650},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266651},
'{step_type : REG_WRITE,	value : 32'd19544,	reg_addr : 32'd266652},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266653},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd266654},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266655},
'{step_type : REG_WRITE,	value : 32'd35928,	reg_addr : 32'd266656},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266657},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd266658},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266659},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266660},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266661},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266662},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266663},
'{step_type : REG_WRITE,	value : 32'd20312,	reg_addr : 32'd266664},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266665},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd266666},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266667},
'{step_type : REG_WRITE,	value : 32'd36696,	reg_addr : 32'd266668},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266669},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd266670},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266671},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266672},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266673},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266674},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266675},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266676},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266677},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266678},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266679},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266680},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266681},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266682},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266683},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266684},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266685},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266686},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266687},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266688},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266689},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266690},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266691},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266692},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266693},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266694},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266695},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266696},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266697},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266698},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266699},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266700},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266701},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266702},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266703},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266704},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266705},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266706},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266707},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266708},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266709},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266710},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266711},
'{step_type : REG_WRITE,	value : 32'd18264,	reg_addr : 32'd266712},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266713},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266714},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266715},
'{step_type : REG_WRITE,	value : 32'd34648,	reg_addr : 32'd266716},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266717},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266718},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266719},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266720},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266721},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266722},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266723},
'{step_type : REG_WRITE,	value : 32'd18392,	reg_addr : 32'd266724},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266725},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266726},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266727},
'{step_type : REG_WRITE,	value : 32'd34776,	reg_addr : 32'd266728},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266729},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266730},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266731},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266732},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266733},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266734},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266735},
'{step_type : REG_WRITE,	value : 32'd19544,	reg_addr : 32'd266736},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266737},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd266738},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266739},
'{step_type : REG_WRITE,	value : 32'd35928,	reg_addr : 32'd266740},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266741},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd266742},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266743},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266744},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266745},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266746},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266747},
'{step_type : REG_WRITE,	value : 32'd20312,	reg_addr : 32'd266748},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266749},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd266750},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266751},
'{step_type : REG_WRITE,	value : 32'd36696,	reg_addr : 32'd266752},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266753},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd266754},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266755},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266756},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266757},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266758},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266759},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266760},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266761},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266762},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266763},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266764},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266765},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266766},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266767},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266768},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266769},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266770},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266771},
'{step_type : REG_WRITE,	value : 32'd51672,	reg_addr : 32'd266772},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266773},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266774},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266775},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266776},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266777},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266778},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266779},
'{step_type : REG_WRITE,	value : 32'd51544,	reg_addr : 32'd266780},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266781},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266782},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266783},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266784},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266785},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266786},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266787},
'{step_type : REG_WRITE,	value : 32'd49368,	reg_addr : 32'd266788},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266789},
'{step_type : REG_WRITE,	value : 32'd59400,	reg_addr : 32'd266790},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266791},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266792},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266793},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266794},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266795},
'{step_type : REG_WRITE,	value : 32'd49496,	reg_addr : 32'd266796},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266797},
'{step_type : REG_WRITE,	value : 32'd60040,	reg_addr : 32'd266798},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266799},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266800},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266801},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266802},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266803},
'{step_type : REG_WRITE,	value : 32'd49624,	reg_addr : 32'd266804},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266805},
'{step_type : REG_WRITE,	value : 32'd50952,	reg_addr : 32'd266806},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266807},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266808},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266809},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266810},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266811},
'{step_type : REG_WRITE,	value : 32'd50520,	reg_addr : 32'd266812},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266813},
'{step_type : REG_WRITE,	value : 32'd59912,	reg_addr : 32'd266814},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266815},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266816},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266817},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266818},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266819},
'{step_type : REG_WRITE,	value : 32'd50648,	reg_addr : 32'd266820},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266821},
'{step_type : REG_WRITE,	value : 32'd57864,	reg_addr : 32'd266822},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266823},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266824},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266825},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266826},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266827},
'{step_type : REG_WRITE,	value : 32'd18648,	reg_addr : 32'd266828},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266829},
'{step_type : REG_WRITE,	value : 32'd16968,	reg_addr : 32'd266830},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266831},
'{step_type : REG_WRITE,	value : 32'd35032,	reg_addr : 32'd266832},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266833},
'{step_type : REG_WRITE,	value : 32'd38472,	reg_addr : 32'd266834},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266835},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266836},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266837},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266838},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266839},
'{step_type : REG_WRITE,	value : 32'd51800,	reg_addr : 32'd266840},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266841},
'{step_type : REG_WRITE,	value : 32'd49416,	reg_addr : 32'd266842},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266843},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266844},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266845},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266846},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266847},
'{step_type : REG_WRITE,	value : 32'd52056,	reg_addr : 32'd266848},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266849},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd266850},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266851},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266852},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266853},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266854},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266855},
'{step_type : REG_WRITE,	value : 32'd54488,	reg_addr : 32'd266856},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266857},
'{step_type : REG_WRITE,	value : 32'd61448,	reg_addr : 32'd266858},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266859},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266860},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266861},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266862},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266863},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266864},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266865},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266866},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266867},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266868},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266869},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266870},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266871},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266872},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266873},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266874},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266875},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266876},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266877},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266878},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266879},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266880},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266881},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266882},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266883},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266884},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266885},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266886},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266887},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266888},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266889},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266890},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266891},
'{step_type : REG_WRITE,	value : 32'd18264,	reg_addr : 32'd266892},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266893},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266894},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266895},
'{step_type : REG_WRITE,	value : 32'd34648,	reg_addr : 32'd266896},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266897},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266898},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266899},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266900},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266901},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266902},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266903},
'{step_type : REG_WRITE,	value : 32'd18392,	reg_addr : 32'd266904},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266905},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266906},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266907},
'{step_type : REG_WRITE,	value : 32'd34776,	reg_addr : 32'd266908},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266909},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266910},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266911},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266912},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266913},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266914},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266915},
'{step_type : REG_WRITE,	value : 32'd19544,	reg_addr : 32'd266916},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266917},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd266918},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266919},
'{step_type : REG_WRITE,	value : 32'd35928,	reg_addr : 32'd266920},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266921},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd266922},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266923},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266924},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266925},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266926},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266927},
'{step_type : REG_WRITE,	value : 32'd20312,	reg_addr : 32'd266928},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266929},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd266930},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266931},
'{step_type : REG_WRITE,	value : 32'd36696,	reg_addr : 32'd266932},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266933},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd266934},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266935},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266936},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266937},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266938},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266939},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266940},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266941},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266942},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266943},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266944},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266945},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266946},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266947},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266948},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266949},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266950},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266951},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266952},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266953},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266954},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266955},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266956},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266957},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266958},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266959},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266960},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266961},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266962},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266963},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd266964},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266965},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266966},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266967},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd266968},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266969},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266970},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266971},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266972},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266973},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266974},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266975},
'{step_type : REG_WRITE,	value : 32'd18264,	reg_addr : 32'd266976},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266977},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266978},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266979},
'{step_type : REG_WRITE,	value : 32'd34648,	reg_addr : 32'd266980},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266981},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266982},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266983},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266984},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266985},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266986},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266987},
'{step_type : REG_WRITE,	value : 32'd18392,	reg_addr : 32'd266988},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266989},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd266990},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266991},
'{step_type : REG_WRITE,	value : 32'd34776,	reg_addr : 32'd266992},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266993},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd266994},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266995},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266996},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd266997},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266998},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd266999},
'{step_type : REG_WRITE,	value : 32'd19544,	reg_addr : 32'd267000},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267001},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd267002},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267003},
'{step_type : REG_WRITE,	value : 32'd35928,	reg_addr : 32'd267004},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267005},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd267006},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267007},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267008},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267009},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267010},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267011},
'{step_type : REG_WRITE,	value : 32'd20312,	reg_addr : 32'd267012},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267013},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd267014},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267015},
'{step_type : REG_WRITE,	value : 32'd36696,	reg_addr : 32'd267016},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267017},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd267018},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267019},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267020},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267021},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267022},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267023},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267024},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267025},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267026},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267027},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267028},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267029},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267030},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267031},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267032},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267033},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267034},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267035},
'{step_type : REG_WRITE,	value : 32'd51672,	reg_addr : 32'd267036},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267037},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267038},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267039},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267040},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267041},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267042},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267043},
'{step_type : REG_WRITE,	value : 32'd51544,	reg_addr : 32'd267044},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267045},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267046},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267047},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267048},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267049},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267050},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267051},
'{step_type : REG_WRITE,	value : 32'd49368,	reg_addr : 32'd267052},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267053},
'{step_type : REG_WRITE,	value : 32'd59400,	reg_addr : 32'd267054},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267055},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267056},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267057},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267058},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267059},
'{step_type : REG_WRITE,	value : 32'd49496,	reg_addr : 32'd267060},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267061},
'{step_type : REG_WRITE,	value : 32'd60040,	reg_addr : 32'd267062},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267063},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267064},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267065},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267066},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267067},
'{step_type : REG_WRITE,	value : 32'd49624,	reg_addr : 32'd267068},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267069},
'{step_type : REG_WRITE,	value : 32'd50952,	reg_addr : 32'd267070},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267071},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267072},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267073},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267074},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267075},
'{step_type : REG_WRITE,	value : 32'd50520,	reg_addr : 32'd267076},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267077},
'{step_type : REG_WRITE,	value : 32'd59912,	reg_addr : 32'd267078},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267079},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267080},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267081},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267082},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267083},
'{step_type : REG_WRITE,	value : 32'd50648,	reg_addr : 32'd267084},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267085},
'{step_type : REG_WRITE,	value : 32'd57864,	reg_addr : 32'd267086},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267087},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267088},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267089},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267090},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267091},
'{step_type : REG_WRITE,	value : 32'd18648,	reg_addr : 32'd267092},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267093},
'{step_type : REG_WRITE,	value : 32'd16968,	reg_addr : 32'd267094},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267095},
'{step_type : REG_WRITE,	value : 32'd35032,	reg_addr : 32'd267096},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267097},
'{step_type : REG_WRITE,	value : 32'd38472,	reg_addr : 32'd267098},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267099},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267100},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267101},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267102},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267103},
'{step_type : REG_WRITE,	value : 32'd51800,	reg_addr : 32'd267104},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267105},
'{step_type : REG_WRITE,	value : 32'd49416,	reg_addr : 32'd267106},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267107},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267108},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267109},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267110},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267111},
'{step_type : REG_WRITE,	value : 32'd52056,	reg_addr : 32'd267112},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267113},
'{step_type : REG_WRITE,	value : 32'd49160,	reg_addr : 32'd267114},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267115},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267116},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267117},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267118},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267119},
'{step_type : REG_WRITE,	value : 32'd54488,	reg_addr : 32'd267120},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267121},
'{step_type : REG_WRITE,	value : 32'd61448,	reg_addr : 32'd267122},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267123},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267124},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267125},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267126},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267127},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267128},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267129},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267130},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267131},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd267132},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267133},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd267134},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267135},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd267136},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267137},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd267138},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267139},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267140},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267141},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267142},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267143},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd267144},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267145},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd267146},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267147},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd267148},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267149},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd267150},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267151},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267152},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267153},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267154},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267155},
'{step_type : REG_WRITE,	value : 32'd18264,	reg_addr : 32'd267156},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267157},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd267158},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267159},
'{step_type : REG_WRITE,	value : 32'd34648,	reg_addr : 32'd267160},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267161},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd267162},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267163},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267164},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267165},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267166},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267167},
'{step_type : REG_WRITE,	value : 32'd18392,	reg_addr : 32'd267168},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267169},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd267170},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267171},
'{step_type : REG_WRITE,	value : 32'd34776,	reg_addr : 32'd267172},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267173},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd267174},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267175},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267176},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267177},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267178},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267179},
'{step_type : REG_WRITE,	value : 32'd19544,	reg_addr : 32'd267180},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267181},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd267182},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267183},
'{step_type : REG_WRITE,	value : 32'd35928,	reg_addr : 32'd267184},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267185},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd267186},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267187},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267188},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267189},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267190},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267191},
'{step_type : REG_WRITE,	value : 32'd20312,	reg_addr : 32'd267192},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267193},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd267194},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267195},
'{step_type : REG_WRITE,	value : 32'd36696,	reg_addr : 32'd267196},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267197},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd267198},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267199},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267200},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267201},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267202},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267203},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267204},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267205},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267206},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267207},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267208},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267209},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267210},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267211},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267212},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267213},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267214},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267215},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd267216},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267217},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd267218},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267219},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd267220},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267221},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd267222},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267223},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267224},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267225},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267226},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267227},
'{step_type : REG_WRITE,	value : 32'd18008,	reg_addr : 32'd267228},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267229},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd267230},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267231},
'{step_type : REG_WRITE,	value : 32'd34392,	reg_addr : 32'd267232},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267233},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd267234},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267235},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267236},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267237},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267238},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267239},
'{step_type : REG_WRITE,	value : 32'd18264,	reg_addr : 32'd267240},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267241},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd267242},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267243},
'{step_type : REG_WRITE,	value : 32'd34648,	reg_addr : 32'd267244},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267245},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd267246},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267247},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267248},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267249},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267250},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267251},
'{step_type : REG_WRITE,	value : 32'd18392,	reg_addr : 32'd267252},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267253},
'{step_type : REG_WRITE,	value : 32'd26632,	reg_addr : 32'd267254},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267255},
'{step_type : REG_WRITE,	value : 32'd34776,	reg_addr : 32'd267256},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267257},
'{step_type : REG_WRITE,	value : 32'd43016,	reg_addr : 32'd267258},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267259},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267260},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267261},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267262},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267263},
'{step_type : REG_WRITE,	value : 32'd19544,	reg_addr : 32'd267264},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267265},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd267266},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267267},
'{step_type : REG_WRITE,	value : 32'd35928,	reg_addr : 32'd267268},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267269},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd267270},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267271},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267272},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267273},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267274},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267275},
'{step_type : REG_WRITE,	value : 32'd20312,	reg_addr : 32'd267276},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267277},
'{step_type : REG_WRITE,	value : 32'd16392,	reg_addr : 32'd267278},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267279},
'{step_type : REG_WRITE,	value : 32'd36696,	reg_addr : 32'd267280},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267281},
'{step_type : REG_WRITE,	value : 32'd32776,	reg_addr : 32'd267282},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267283},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267284},
'{step_type : REG_WRITE,	value : 32'd721420288,	reg_addr : 32'd267285},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267286},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267287},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267288},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267289},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267290},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267291},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267292},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267293},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267294},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267295},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267296},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267297},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267298},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd267299},
'{step_type : REG_WRITE,	value : 32'd1024,	reg_addr : 32'd852199},
'{step_type : REG_WRITE,	value : 32'd22561,	reg_addr : 32'd786433},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591628},
'{step_type : REG_WRITE,	value : 32'd254,	reg_addr : 32'd591629},
'{step_type : REG_WRITE,	value : 32'd65535,	reg_addr : 32'd591630},
'{step_type : REG_WRITE,	value : 32'd61504,	reg_addr : 32'd591631},
'{step_type : REG_WRITE,	value : 32'd61504,	reg_addr : 32'd591632},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591633},
'{step_type : REG_WRITE,	value : 32'd65535,	reg_addr : 32'd591634},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591635},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591636},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591637},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591638},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591639},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591640},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591641},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591642},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd591643},
'{step_type : REG_WRITE,	value : 32'd2925,	reg_addr : 32'd458992},
'{step_type : REG_WRITE,	value : 32'd195,	reg_addr : 32'd458878},
'{step_type : REG_WRITE,	value : 32'd32767,	reg_addr : 32'd459247},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd196774},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd200870},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459176},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459048},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459057},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459058},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459059},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459060},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459074},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd459076},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd786560},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd851968},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd851968},
'{step_type : REG_WRITE,	value : 32'd7,	reg_addr : 32'd786560},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd720897},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd131079},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd196642},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd200738},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd16496},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd20592},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd45168},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd49264},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd1065072},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd1069168},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd1093744},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd1097840},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd2113648},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd2117744},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd2142320},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd2146416},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd3162224},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd3166320},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd3190896},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd3194992},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd655362},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd131237},
'{step_type : POLL,	value : 32'd2047,	reg_addr : 32'd65687},
'{step_type : POLL,	value : 32'd2047,	reg_addr : 32'd69783},
'{step_type : POLL,	value : 32'd2047,	reg_addr : 32'd73879},
'{step_type : POLL,	value : 32'd2047,	reg_addr : 32'd77975},
'{step_type : POLL,	value : 32'd9,	reg_addr : 32'd721667},
'{step_type : POLL,	value : 32'd38,	reg_addr : 32'd656130},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd721665},
'{step_type : POLL,	value : 32'd29,	reg_addr : 32'd721679},
'{step_type : POLL,	value : 32'd6272,	reg_addr : 32'd196782},
'{step_type : POLL,	value : 32'd6272,	reg_addr : 32'd196781},
'{step_type : POLL,	value : 32'd6272,	reg_addr : 32'd196780},
'{step_type : POLL,	value : 32'd6272,	reg_addr : 32'd200878},
'{step_type : POLL,	value : 32'd6272,	reg_addr : 32'd200877},
'{step_type : POLL,	value : 32'd6272,	reg_addr : 32'd200876},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd786566},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459035},
'{step_type : POLL,	value : 32'd2099,	reg_addr : 32'd65699},
'{step_type : POLL,	value : 32'd2099,	reg_addr : 32'd69795},
'{step_type : POLL,	value : 32'd2099,	reg_addr : 32'd73891},
'{step_type : POLL,	value : 32'd2099,	reg_addr : 32'd77987},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd786672},
'{step_type : POLL,	value : 32'd2,	reg_addr : 32'd786673},
'{step_type : POLL,	value : 32'd7,	reg_addr : 32'd786674},
'{step_type : POLL,	value : 32'd52,	reg_addr : 32'd786675},
'{step_type : POLL,	value : 32'd45,	reg_addr : 32'd591667},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd786676},
'{step_type : POLL,	value : 32'd61440,	reg_addr : 32'd786679},
'{step_type : POLL,	value : 32'd2560,	reg_addr : 32'd591671},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd591647},
'{step_type : POLL,	value : 32'd15,	reg_addr : 32'd591913},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917626},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd921722},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925818},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd929914},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934010},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd938106},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942202},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd946298},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1566},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd5662},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd9758},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd13854},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd17950},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd22046},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd30238},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd34334},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd38430},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd42526},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd46622},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd50718},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69151},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73247},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd77343},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd81439},
'{step_type : POLL,	value : 32'd61030,	reg_addr : 32'd198663},
'{step_type : POLL,	value : 32'd61030,	reg_addr : 32'd202759},
'{step_type : POLL,	value : 32'd61030,	reg_addr : 32'd67591},
'{step_type : POLL,	value : 32'd61030,	reg_addr : 32'd71687},
'{step_type : POLL,	value : 32'd61030,	reg_addr : 32'd75783},
'{step_type : POLL,	value : 32'd61030,	reg_addr : 32'd79879},
'{step_type : POLL,	value : 32'd16383,	reg_addr : 32'd196768},
'{step_type : POLL,	value : 32'd16383,	reg_addr : 32'd200864},
'{step_type : POLL,	value : 32'd8191,	reg_addr : 32'd65673},
'{step_type : POLL,	value : 32'd2047,	reg_addr : 32'd65674},
'{step_type : POLL,	value : 32'd8191,	reg_addr : 32'd69769},
'{step_type : POLL,	value : 32'd2047,	reg_addr : 32'd69770},
'{step_type : POLL,	value : 32'd8191,	reg_addr : 32'd73865},
'{step_type : POLL,	value : 32'd2047,	reg_addr : 32'd73866},
'{step_type : POLL,	value : 32'd8191,	reg_addr : 32'd77961},
'{step_type : POLL,	value : 32'd2047,	reg_addr : 32'd77962},
'{step_type : POLL,	value : 32'd15,	reg_addr : 32'd131078},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd131084},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd917517},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd921613},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd925709},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd929805},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd933901},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd937997},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd942093},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd946189},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd196647},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd63},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd4159},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd8255},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd12351},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd16447},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd20543},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd200743},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd28735},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd32831},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd36927},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd41023},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd45119},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd49215},
'{step_type : POLL,	value : 32'd49314,	reg_addr : 32'd591873},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591874},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd591878},
'{step_type : POLL,	value : 32'd16641,	reg_addr : 32'd656383},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd656139},
'{step_type : POLL,	value : 32'd11606,	reg_addr : 32'd393224},
'{step_type : POLL,	value : 32'd100,	reg_addr : 32'd592096},
'{step_type : POLL,	value : 32'd300,	reg_addr : 32'd592097},
'{step_type : POLL,	value : 32'd2000,	reg_addr : 32'd592098},
'{step_type : POLL,	value : 32'd88,	reg_addr : 32'd592099},
'{step_type : POLL,	value : 32'd20,	reg_addr : 32'd592100},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd592101},
'{step_type : POLL,	value : 32'd67,	reg_addr : 32'd592102},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd592103},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd592106},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd592107},
'{step_type : POLL,	value : 32'd10,	reg_addr : 32'd592108},
'{step_type : POLL,	value : 32'd78,	reg_addr : 32'd592109},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd131074},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd393280},
'{step_type : POLL,	value : 32'd2,	reg_addr : 32'd131072},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65787},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69883},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73979},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78075},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917515},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921611},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925707},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929803},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933899},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd937995},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942091},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946187},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd65572},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd69668},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd73764},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd77860},
'{step_type : POLL,	value : 32'd44,	reg_addr : 32'd65573},
'{step_type : POLL,	value : 32'd44,	reg_addr : 32'd69669},
'{step_type : POLL,	value : 32'd44,	reg_addr : 32'd73765},
'{step_type : POLL,	value : 32'd44,	reg_addr : 32'd77861},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65540},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65539},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69636},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69635},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73732},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73731},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd77828},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd77827},
'{step_type : POLL,	value : 32'd800,	reg_addr : 32'd720900},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd656140},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd65598},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd69694},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd73790},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd77886},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd131075},
'{step_type : POLL,	value : 32'd4369,	reg_addr : 32'd131083},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65800},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69896},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73992},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78088},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd458757},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd458767},
'{step_type : POLL,	value : 32'd4864,	reg_addr : 32'd65550},
'{step_type : POLL,	value : 32'd4864,	reg_addr : 32'd69646},
'{step_type : POLL,	value : 32'd4864,	reg_addr : 32'd73742},
'{step_type : POLL,	value : 32'd4864,	reg_addr : 32'd77838},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd131097},
'{step_type : POLL,	value : 32'd51,	reg_addr : 32'd917548},
'{step_type : POLL,	value : 32'd51,	reg_addr : 32'd921644},
'{step_type : POLL,	value : 32'd771,	reg_addr : 32'd917549},
'{step_type : POLL,	value : 32'd13107,	reg_addr : 32'd921645},
'{step_type : POLL,	value : 32'd51,	reg_addr : 32'd925740},
'{step_type : POLL,	value : 32'd51,	reg_addr : 32'd929836},
'{step_type : POLL,	value : 32'd771,	reg_addr : 32'd925741},
'{step_type : POLL,	value : 32'd13107,	reg_addr : 32'd929837},
'{step_type : POLL,	value : 32'd51,	reg_addr : 32'd933932},
'{step_type : POLL,	value : 32'd51,	reg_addr : 32'd938028},
'{step_type : POLL,	value : 32'd771,	reg_addr : 32'd933933},
'{step_type : POLL,	value : 32'd13107,	reg_addr : 32'd938029},
'{step_type : POLL,	value : 32'd51,	reg_addr : 32'd942124},
'{step_type : POLL,	value : 32'd51,	reg_addr : 32'd946220},
'{step_type : POLL,	value : 32'd771,	reg_addr : 32'd942125},
'{step_type : POLL,	value : 32'd13107,	reg_addr : 32'd946221},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd112},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd4208},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd8304},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd12400},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd28784},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd32880},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd36976},
'{step_type : POLL,	value : 32'd119,	reg_addr : 32'd41072},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd917550},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd921646},
'{step_type : POLL,	value : 32'd13056,	reg_addr : 32'd917551},
'{step_type : POLL,	value : 32'd30464,	reg_addr : 32'd921647},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd925742},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd929838},
'{step_type : POLL,	value : 32'd13056,	reg_addr : 32'd925743},
'{step_type : POLL,	value : 32'd30464,	reg_addr : 32'd929839},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd933934},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd938030},
'{step_type : POLL,	value : 32'd13056,	reg_addr : 32'd933935},
'{step_type : POLL,	value : 32'd30464,	reg_addr : 32'd938031},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd942126},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd946222},
'{step_type : POLL,	value : 32'd13056,	reg_addr : 32'd942127},
'{step_type : POLL,	value : 32'd30464,	reg_addr : 32'd946223},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd121},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd4217},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd8313},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd12409},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd16505},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd20601},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd28793},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd32889},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd36985},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd41081},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd45177},
'{step_type : POLL,	value : 32'd48,	reg_addr : 32'd49273},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd917532},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd921628},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd925724},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd929820},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd933916},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd938012},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd942108},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd946204},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd109},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd4205},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd8301},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd12397},
'{step_type : POLL,	value : 32'd248,	reg_addr : 32'd16493},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd20589},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd28781},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd32877},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd36973},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd41069},
'{step_type : POLL,	value : 32'd248,	reg_addr : 32'd45165},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd49261},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917566},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921662},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925758},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929854},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933950},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938046},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942142},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946238},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65537},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69633},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73729},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd77825},
'{step_type : POLL,	value : 32'd91,	reg_addr : 32'd458816},
'{step_type : POLL,	value : 32'd15,	reg_addr : 32'd458817},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd65701},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd69797},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd73893},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd77989},
'{step_type : POLL,	value : 32'd12850,	reg_addr : 32'd66057},
'{step_type : POLL,	value : 32'd12850,	reg_addr : 32'd70153},
'{step_type : POLL,	value : 32'd12850,	reg_addr : 32'd74249},
'{step_type : POLL,	value : 32'd12850,	reg_addr : 32'd78345},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd66063},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd70159},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd74255},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd78351},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd131077},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd65544},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd69640},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd73736},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd77832},
'{step_type : POLL,	value : 32'd546,	reg_addr : 32'd458859},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd458854},
'{step_type : POLL,	value : 32'd546,	reg_addr : 32'd458987},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd458982},
'{step_type : POLL,	value : 32'd4108,	reg_addr : 32'd459061},
'{step_type : POLL,	value : 32'd4108,	reg_addr : 32'd459062},
'{step_type : POLL,	value : 32'd1052,	reg_addr : 32'd459063},
'{step_type : POLL,	value : 32'd6944,	reg_addr : 32'd459064},
'{step_type : POLL,	value : 32'd4124,	reg_addr : 32'd459065},
'{step_type : POLL,	value : 32'd4124,	reg_addr : 32'd459066},
'{step_type : POLL,	value : 32'd1068,	reg_addr : 32'd459067},
'{step_type : POLL,	value : 32'd12080,	reg_addr : 32'd459068},
'{step_type : POLL,	value : 32'd4100,	reg_addr : 32'd459069},
'{step_type : POLL,	value : 32'd4100,	reg_addr : 32'd459070},
'{step_type : POLL,	value : 32'd1044,	reg_addr : 32'd459071},
'{step_type : POLL,	value : 32'd4888,	reg_addr : 32'd459072},
'{step_type : POLL,	value : 32'd2107,	reg_addr : 32'd459052},
'{step_type : POLL,	value : 32'd2107,	reg_addr : 32'd459053},
'{step_type : POLL,	value : 32'd2107,	reg_addr : 32'd459056},
'{step_type : POLL,	value : 32'd2079,	reg_addr : 32'd459054},
'{step_type : POLL,	value : 32'd2079,	reg_addr : 32'd459055},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd196616},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd200712},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917523},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921619},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925715},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929811},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933907},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938003},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942099},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946195},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd1507},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd5603},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd9699},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd13795},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd17891},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd21987},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd30179},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd34275},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd38371},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd42467},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd46563},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd50659},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd919011},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd923107},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd927203},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd931299},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd935395},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd939491},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd943587},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd947683},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1290},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd5386},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd9482},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd13578},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd17674},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd21770},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd29962},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd34058},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd38154},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd42250},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd46346},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd50442},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd67595},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd71691},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd75787},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd79883},
'{step_type : POLL,	value : 32'd4202,	reg_addr : 32'd198659},
'{step_type : POLL,	value : 32'd4202,	reg_addr : 32'd202755},
'{step_type : POLL,	value : 32'd4202,	reg_addr : 32'd67587},
'{step_type : POLL,	value : 32'd4202,	reg_addr : 32'd71683},
'{step_type : POLL,	value : 32'd4202,	reg_addr : 32'd75779},
'{step_type : POLL,	value : 32'd4202,	reg_addr : 32'd79875},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd1283},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd5379},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd9475},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd13571},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd17667},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd21763},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd29955},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd34051},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd38147},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd42243},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd46339},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd50435},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd68611},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd72707},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd76803},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd80899},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd272},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd4368},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd8464},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd12560},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd16656},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd20752},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd28944},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd33040},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd37136},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd41232},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd45328},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd49424},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd917776},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd921872},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd925968},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd930064},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd934160},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd938256},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd942352},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd946448},
'{step_type : POLL,	value : 32'd19,	reg_addr : 32'd592104},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd592105},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917506},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921602},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925698},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929794},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933890},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd937986},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942082},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946178},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65803},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69899},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73995},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78091},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd99},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd4195},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd8291},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd12387},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd16483},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd20579},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd28771},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd32867},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd36963},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd41059},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd45155},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd49251},
'{step_type : POLL,	value : 32'd610,	reg_addr : 32'd591882},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd591883},
'{step_type : POLL,	value : 32'd610,	reg_addr : 32'd591893},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd591894},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd917603},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd917604},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd917639},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd921699},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd921700},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd921735},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd925795},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd925796},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd925831},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd929891},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd929892},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd929927},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd933987},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd933988},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd934023},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd938083},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd938084},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd938119},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd942179},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd942180},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd942215},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd946275},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd946276},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd946311},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd917564},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd921660},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd925756},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd929852},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd933948},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd938044},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd942140},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd946236},
'{step_type : POLL,	value : 32'd83,	reg_addr : 32'd591895},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591896},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591897},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd196843},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd200939},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd721681},
'{step_type : POLL,	value : 32'd1008,	reg_addr : 32'd393222},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd196629},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd200725},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65660},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69756},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73852},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd77948},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd459073},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591884},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65575},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69671},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73767},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd77863},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd917567},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd917645},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd921663},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd921741},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd925759},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd925837},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd929855},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd929933},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd933951},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd934029},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd938047},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd938125},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd942143},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd942221},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd946239},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd946317},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd592131},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd458866},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd591886},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd458867},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd591887},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266240},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266241},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266242},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266243},
'{step_type : POLL,	value : 32'd49192,	reg_addr : 32'd267348},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267349},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267350},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267351},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267352},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267353},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267354},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267355},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267356},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267357},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267358},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267359},
'{step_type : POLL,	value : 32'd51288,	reg_addr : 32'd267360},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267361},
'{step_type : POLL,	value : 32'd57480,	reg_addr : 32'd267362},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267363},
'{step_type : POLL,	value : 32'd57400,	reg_addr : 32'd267364},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267365},
'{step_type : POLL,	value : 32'd51288,	reg_addr : 32'd267366},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267367},
'{step_type : POLL,	value : 32'd49288,	reg_addr : 32'd267368},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267369},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267370},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267371},
'{step_type : POLL,	value : 32'd49192,	reg_addr : 32'd267372},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267373},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267374},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267375},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267376},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267377},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267378},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267379},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267380},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267381},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267382},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267383},
'{step_type : POLL,	value : 32'd51288,	reg_addr : 32'd267384},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267385},
'{step_type : POLL,	value : 32'd57864,	reg_addr : 32'd267386},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267387},
'{step_type : POLL,	value : 32'd57400,	reg_addr : 32'd267388},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267389},
'{step_type : POLL,	value : 32'd51288,	reg_addr : 32'd267390},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267391},
'{step_type : POLL,	value : 32'd49672,	reg_addr : 32'd267392},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267393},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267394},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267395},
'{step_type : POLL,	value : 32'd49216,	reg_addr : 32'd267396},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267397},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267398},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267399},
'{step_type : POLL,	value : 32'd49256,	reg_addr : 32'd267400},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267401},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267402},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267403},
'{step_type : POLL,	value : 32'd52824,	reg_addr : 32'd267404},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267405},
'{step_type : POLL,	value : 32'd49672,	reg_addr : 32'd267406},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267407},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267408},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267409},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267410},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267411},
'{step_type : POLL,	value : 32'd17264,	reg_addr : 32'd267412},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267413},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267414},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267415},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267416},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267417},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267418},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267419},
'{step_type : POLL,	value : 32'd33648,	reg_addr : 32'd267420},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267421},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267422},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267423},
'{step_type : POLL,	value : 32'd53976,	reg_addr : 32'd267424},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267425},
'{step_type : POLL,	value : 32'd57352,	reg_addr : 32'd267426},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267427},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267428},
'{step_type : POLL,	value : 32'd2063597568,	reg_addr : 32'd267429},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267430},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267431},
'{step_type : POLL,	value : 32'd49392,	reg_addr : 32'd267432},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267433},
'{step_type : POLL,	value : 32'd53208,	reg_addr : 32'd267434},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267435},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267436},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267437},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267438},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267439},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267440},
'{step_type : POLL,	value : 32'd989855744,	reg_addr : 32'd267441},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267442},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267443},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267444},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267445},
'{step_type : POLL,	value : 32'd53336,	reg_addr : 32'd267446},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267447},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267448},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267449},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267450},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267451},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267452},
'{step_type : POLL,	value : 32'd989855744,	reg_addr : 32'd267453},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267454},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267455},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267456},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267457},
'{step_type : POLL,	value : 32'd53464,	reg_addr : 32'd267458},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267459},
'{step_type : POLL,	value : 32'd49288,	reg_addr : 32'd267460},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267461},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267462},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267463},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267464},
'{step_type : POLL,	value : 32'd989855744,	reg_addr : 32'd267465},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267466},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267467},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267468},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267469},
'{step_type : POLL,	value : 32'd53592,	reg_addr : 32'd267470},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267471},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267472},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267473},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267474},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267475},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267476},
'{step_type : POLL,	value : 32'd1795162112,	reg_addr : 32'd267477},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267478},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267479},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267480},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267481},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267482},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267483},
'{step_type : POLL,	value : 32'd218120236,	reg_addr : 32'd267484},
'{step_type : POLL,	value : 32'd67108865,	reg_addr : 32'd267485},
'{step_type : POLL,	value : 32'd134234192,	reg_addr : 32'd267486},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267487},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267488},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267489},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267490},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267491},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267492},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267493},
'{step_type : POLL,	value : 32'd134430800,	reg_addr : 32'd267494},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267495},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267496},
'{step_type : POLL,	value : 32'd520093696,	reg_addr : 32'd267497},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267498},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267499},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267500},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267501},
'{step_type : POLL,	value : 32'd16508,	reg_addr : 32'd267502},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267503},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267504},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267505},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267506},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267507},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267508},
'{step_type : POLL,	value : 32'd67108865,	reg_addr : 32'd267509},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267510},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267511},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267512},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267513},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267514},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267515},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267516},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267517},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267518},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267519},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267520},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267521},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267522},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267523},
'{step_type : POLL,	value : 32'd218136620,	reg_addr : 32'd267524},
'{step_type : POLL,	value : 32'd68157441,	reg_addr : 32'd267525},
'{step_type : POLL,	value : 32'd134250576,	reg_addr : 32'd267526},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267527},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267528},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267529},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267530},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267531},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267532},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267533},
'{step_type : POLL,	value : 32'd134447184,	reg_addr : 32'd267534},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267535},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267536},
'{step_type : POLL,	value : 32'd520093696,	reg_addr : 32'd267537},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267538},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267539},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267540},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267541},
'{step_type : POLL,	value : 32'd32892,	reg_addr : 32'd267542},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267543},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267544},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267545},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267546},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267547},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267548},
'{step_type : POLL,	value : 32'd67108865,	reg_addr : 32'd267549},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267550},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267551},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267552},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267553},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267554},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267555},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267556},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267557},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267558},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267559},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267560},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267561},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267562},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267563},
'{step_type : POLL,	value : 32'd218120236,	reg_addr : 32'd267564},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267565},
'{step_type : POLL,	value : 32'd134234192,	reg_addr : 32'd267566},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267567},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267568},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267569},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267570},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267571},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267572},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267573},
'{step_type : POLL,	value : 32'd134430800,	reg_addr : 32'd267574},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267575},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267576},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267577},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267578},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267579},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267580},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267581},
'{step_type : POLL,	value : 32'd134430800,	reg_addr : 32'd267582},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267583},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267584},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267585},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267586},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267587},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267588},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267589},
'{step_type : POLL,	value : 32'd134234192,	reg_addr : 32'd267590},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267591},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267592},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267593},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267594},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267595},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267596},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267597},
'{step_type : POLL,	value : 32'd16508,	reg_addr : 32'd267598},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267599},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267600},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267601},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267602},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267603},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267604},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267605},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267606},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267607},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267608},
'{step_type : POLL,	value : 32'd1526726656,	reg_addr : 32'd267609},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267610},
'{step_type : POLL,	value : 32'd469762048,	reg_addr : 32'd267611},
'{step_type : POLL,	value : 32'd218136620,	reg_addr : 32'd267612},
'{step_type : POLL,	value : 32'd1048577,	reg_addr : 32'd267613},
'{step_type : POLL,	value : 32'd134250576,	reg_addr : 32'd267614},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267615},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267616},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267617},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267618},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267619},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267620},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267621},
'{step_type : POLL,	value : 32'd134447184,	reg_addr : 32'd267622},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267623},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267624},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267625},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267626},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267627},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267628},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267629},
'{step_type : POLL,	value : 32'd134447184,	reg_addr : 32'd267630},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267631},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267632},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267633},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267634},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267635},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267636},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267637},
'{step_type : POLL,	value : 32'd134250576,	reg_addr : 32'd267638},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267639},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267640},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267641},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267642},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267643},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267644},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267645},
'{step_type : POLL,	value : 32'd32892,	reg_addr : 32'd267646},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267647},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267648},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267649},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267650},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267651},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267652},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267653},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267654},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267655},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267656},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd267657},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267658},
'{step_type : POLL,	value : 32'd671088640,	reg_addr : 32'd267659},
'{step_type : POLL,	value : 32'd218120236,	reg_addr : 32'd267660},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267661},
'{step_type : POLL,	value : 32'd134435224,	reg_addr : 32'd267662},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267663},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267664},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267665},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267666},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267667},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267668},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267669},
'{step_type : POLL,	value : 32'd134435352,	reg_addr : 32'd267670},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267671},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267672},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267673},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267674},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267675},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267676},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267677},
'{step_type : POLL,	value : 32'd16508,	reg_addr : 32'd267678},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267679},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267680},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267681},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267682},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267683},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267684},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267685},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267686},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267687},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267688},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267689},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267690},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267691},
'{step_type : POLL,	value : 32'd218136620,	reg_addr : 32'd267692},
'{step_type : POLL,	value : 32'd1048577,	reg_addr : 32'd267693},
'{step_type : POLL,	value : 32'd134451608,	reg_addr : 32'd267694},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267695},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267696},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267697},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267698},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267699},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267700},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267701},
'{step_type : POLL,	value : 32'd134451736,	reg_addr : 32'd267702},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267703},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267704},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267705},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267706},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267707},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267708},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267709},
'{step_type : POLL,	value : 32'd32892,	reg_addr : 32'd267710},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267711},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267712},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267713},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267714},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267715},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267716},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267717},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267718},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267719},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267720},
'{step_type : POLL,	value : 32'd989855744,	reg_addr : 32'd267721},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267722},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267723},
'{step_type : POLL,	value : 32'd53976,	reg_addr : 32'd267724},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267725},
'{step_type : POLL,	value : 32'd57352,	reg_addr : 32'd267726},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267727},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267728},
'{step_type : POLL,	value : 32'd2063597568,	reg_addr : 32'd267729},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267730},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267731},
'{step_type : POLL,	value : 32'd49392,	reg_addr : 32'd267732},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267733},
'{step_type : POLL,	value : 32'd53208,	reg_addr : 32'd267734},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267735},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267736},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267737},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267738},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267739},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267740},
'{step_type : POLL,	value : 32'd989855744,	reg_addr : 32'd267741},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267742},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267743},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267744},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267745},
'{step_type : POLL,	value : 32'd53336,	reg_addr : 32'd267746},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267747},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267748},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267749},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267750},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267751},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267752},
'{step_type : POLL,	value : 32'd989855744,	reg_addr : 32'd267753},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267754},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267755},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267756},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267757},
'{step_type : POLL,	value : 32'd53464,	reg_addr : 32'd267758},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267759},
'{step_type : POLL,	value : 32'd49288,	reg_addr : 32'd267760},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267761},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267762},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267763},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267764},
'{step_type : POLL,	value : 32'd989855744,	reg_addr : 32'd267765},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267766},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267767},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267768},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267769},
'{step_type : POLL,	value : 32'd53592,	reg_addr : 32'd267770},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267771},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267772},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267773},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267774},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267775},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267776},
'{step_type : POLL,	value : 32'd1795162112,	reg_addr : 32'd267777},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267778},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267779},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267780},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267781},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267782},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267783},
'{step_type : POLL,	value : 32'd218120236,	reg_addr : 32'd267784},
'{step_type : POLL,	value : 32'd67108865,	reg_addr : 32'd267785},
'{step_type : POLL,	value : 32'd134234192,	reg_addr : 32'd267786},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267787},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267788},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267789},
'{step_type : POLL,	value : 32'd134430800,	reg_addr : 32'd267790},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267791},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267792},
'{step_type : POLL,	value : 32'd1325400064,	reg_addr : 32'd267793},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267794},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267795},
'{step_type : POLL,	value : 32'd16508,	reg_addr : 32'd267796},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267797},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267798},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267799},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267800},
'{step_type : POLL,	value : 32'd520093696,	reg_addr : 32'd267801},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267802},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267803},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267804},
'{step_type : POLL,	value : 32'd67108865,	reg_addr : 32'd267805},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267806},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267807},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267808},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267809},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267810},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267811},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267812},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267813},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267814},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267815},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267816},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267817},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267818},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267819},
'{step_type : POLL,	value : 32'd218136620,	reg_addr : 32'd267820},
'{step_type : POLL,	value : 32'd68157441,	reg_addr : 32'd267821},
'{step_type : POLL,	value : 32'd134250576,	reg_addr : 32'd267822},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267823},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267824},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267825},
'{step_type : POLL,	value : 32'd134447184,	reg_addr : 32'd267826},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267827},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267828},
'{step_type : POLL,	value : 32'd1325400064,	reg_addr : 32'd267829},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267830},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267831},
'{step_type : POLL,	value : 32'd32892,	reg_addr : 32'd267832},
'{step_type : POLL,	value : 32'd68157440,	reg_addr : 32'd267833},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267834},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267835},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267836},
'{step_type : POLL,	value : 32'd520093696,	reg_addr : 32'd267837},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267838},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267839},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267840},
'{step_type : POLL,	value : 32'd67108865,	reg_addr : 32'd267841},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267842},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267843},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267844},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd267845},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267846},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267847},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267848},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267849},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267850},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267851},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267852},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267853},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267854},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267855},
'{step_type : POLL,	value : 32'd218120236,	reg_addr : 32'd267856},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267857},
'{step_type : POLL,	value : 32'd134234192,	reg_addr : 32'd267858},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267859},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267860},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267861},
'{step_type : POLL,	value : 32'd134430800,	reg_addr : 32'd267862},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267863},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267864},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267865},
'{step_type : POLL,	value : 32'd134430800,	reg_addr : 32'd267866},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267867},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267868},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267869},
'{step_type : POLL,	value : 32'd134234192,	reg_addr : 32'd267870},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267871},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267872},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd267873},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267874},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267875},
'{step_type : POLL,	value : 32'd16508,	reg_addr : 32'd267876},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267877},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267878},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267879},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267880},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267881},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267882},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267883},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267884},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267885},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267886},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267887},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267888},
'{step_type : POLL,	value : 32'd1526726656,	reg_addr : 32'd267889},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267890},
'{step_type : POLL,	value : 32'd469762048,	reg_addr : 32'd267891},
'{step_type : POLL,	value : 32'd218136620,	reg_addr : 32'd267892},
'{step_type : POLL,	value : 32'd1048577,	reg_addr : 32'd267893},
'{step_type : POLL,	value : 32'd134250576,	reg_addr : 32'd267894},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267895},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267896},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267897},
'{step_type : POLL,	value : 32'd134447184,	reg_addr : 32'd267898},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267899},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267900},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267901},
'{step_type : POLL,	value : 32'd134447184,	reg_addr : 32'd267902},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267903},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267904},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267905},
'{step_type : POLL,	value : 32'd134250576,	reg_addr : 32'd267906},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267907},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267908},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd267909},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267910},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267911},
'{step_type : POLL,	value : 32'd32892,	reg_addr : 32'd267912},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267913},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267914},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267915},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267916},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267917},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267918},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267919},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267920},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267921},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267922},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267923},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267924},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267925},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267926},
'{step_type : POLL,	value : 32'd671088640,	reg_addr : 32'd267927},
'{step_type : POLL,	value : 32'd218120236,	reg_addr : 32'd267928},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267929},
'{step_type : POLL,	value : 32'd134435224,	reg_addr : 32'd267930},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267931},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267932},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267933},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267934},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267935},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267936},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267937},
'{step_type : POLL,	value : 32'd134435352,	reg_addr : 32'd267938},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267939},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267940},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd267941},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267942},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267943},
'{step_type : POLL,	value : 32'd16508,	reg_addr : 32'd267944},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267945},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267946},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267947},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267948},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267949},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267950},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267951},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267952},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267953},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267954},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267955},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267956},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267957},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267958},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267959},
'{step_type : POLL,	value : 32'd218136620,	reg_addr : 32'd267960},
'{step_type : POLL,	value : 32'd1048577,	reg_addr : 32'd267961},
'{step_type : POLL,	value : 32'd134451608,	reg_addr : 32'd267962},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267963},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267964},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267965},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267966},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267967},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267968},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267969},
'{step_type : POLL,	value : 32'd134451736,	reg_addr : 32'd267970},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267971},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267972},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd267973},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267974},
'{step_type : POLL,	value : 32'd134217728,	reg_addr : 32'd267975},
'{step_type : POLL,	value : 32'd32892,	reg_addr : 32'd267976},
'{step_type : POLL,	value : 32'd1048576,	reg_addr : 32'd267977},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267978},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267979},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267980},
'{step_type : POLL,	value : 32'd452984832,	reg_addr : 32'd267981},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267982},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267983},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267984},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd267985},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267986},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267987},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267988},
'{step_type : POLL,	value : 32'd1795162112,	reg_addr : 32'd267989},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267990},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267991},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267992},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267993},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267994},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267995},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267996},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267997},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267998},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267999},
'{step_type : POLL,	value : 32'd1065006208,	reg_addr : 32'd278528},
'{step_type : POLL,	value : 32'd91168,	reg_addr : 32'd278529},
'{step_type : POLL,	value : 32'd1024,	reg_addr : 32'd278530},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278531},
'{step_type : POLL,	value : 32'd2147484800,	reg_addr : 32'd278532},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd278533},
'{step_type : POLL,	value : 32'd67111936,	reg_addr : 32'd278534},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278535},
'{step_type : POLL,	value : 32'd2214593664,	reg_addr : 32'd278536},
'{step_type : POLL,	value : 32'd3072,	reg_addr : 32'd278537},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278538},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278539},
'{step_type : POLL,	value : 32'd2214592640,	reg_addr : 32'd278540},
'{step_type : POLL,	value : 32'd3072,	reg_addr : 32'd278541},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278542},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278543},
'{step_type : POLL,	value : 32'd2147910144,	reg_addr : 32'd278544},
'{step_type : POLL,	value : 32'd16399,	reg_addr : 32'd278545},
'{step_type : POLL,	value : 32'd35136,	reg_addr : 32'd278546},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278547},
'{step_type : POLL,	value : 32'd2684355712,	reg_addr : 32'd278548},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd278549},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278550},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278551},
'{step_type : POLL,	value : 32'd2617253024,	reg_addr : 32'd278552},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278553},
'{step_type : POLL,	value : 32'd2818574464,	reg_addr : 32'd278554},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd278555},
'{step_type : POLL,	value : 32'd2147549312,	reg_addr : 32'd278556},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278557},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278558},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278559},
'{step_type : POLL,	value : 32'd2147550336,	reg_addr : 32'd278560},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278561},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278562},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278563},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd278564},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd278565},
'{step_type : POLL,	value : 32'd2684354688,	reg_addr : 32'd278566},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd278567},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd278568},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278569},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd278570},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278571},
'{step_type : POLL,	value : 32'd12320,	reg_addr : 32'd278572},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278573},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd278574},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278575},
'{step_type : POLL,	value : 32'd2818574464,	reg_addr : 32'd278576},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd278577},
'{step_type : POLL,	value : 32'd2147551360,	reg_addr : 32'd278578},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278579},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278580},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278581},
'{step_type : POLL,	value : 32'd2147552384,	reg_addr : 32'd278582},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278583},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278584},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278585},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd278586},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278587},
'{step_type : POLL,	value : 32'd11296,	reg_addr : 32'd278588},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278589},
'{step_type : POLL,	value : 32'd11296,	reg_addr : 32'd278590},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278591},
'{step_type : POLL,	value : 32'd11296,	reg_addr : 32'd278592},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278593},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd278594},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278595},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278596},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278597},
'{step_type : POLL,	value : 32'd2818573440,	reg_addr : 32'd278598},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278599},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278600},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278601},
'{step_type : POLL,	value : 32'd1073758720,	reg_addr : 32'd278602},
'{step_type : POLL,	value : 32'd16384,	reg_addr : 32'd278603},
'{step_type : POLL,	value : 32'd68928,	reg_addr : 32'd278604},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278605},
'{step_type : POLL,	value : 32'd3355457696,	reg_addr : 32'd278606},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278607},
'{step_type : POLL,	value : 32'd3422567584,	reg_addr : 32'd278608},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278609},
'{step_type : POLL,	value : 32'd2751463584,	reg_addr : 32'd278610},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd278611},
'{step_type : POLL,	value : 32'd2818579584,	reg_addr : 32'd278612},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd278613},
'{step_type : POLL,	value : 32'd2147815552,	reg_addr : 32'd278614},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278615},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278616},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278617},
'{step_type : POLL,	value : 32'd2147816576,	reg_addr : 32'd278618},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278619},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278620},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278621},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd278622},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd278623},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd278624},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278625},
'{step_type : POLL,	value : 32'd3422552192,	reg_addr : 32'd278626},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278627},
'{step_type : POLL,	value : 32'd2818579584,	reg_addr : 32'd278628},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd278629},
'{step_type : POLL,	value : 32'd2147817600,	reg_addr : 32'd278630},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278631},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278632},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278633},
'{step_type : POLL,	value : 32'd2147818624,	reg_addr : 32'd278634},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278635},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278636},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278637},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd278638},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd278639},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd278640},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278641},
'{step_type : POLL,	value : 32'd3355443328,	reg_addr : 32'd278642},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278643},
'{step_type : POLL,	value : 32'd3422567584,	reg_addr : 32'd278644},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278645},
'{step_type : POLL,	value : 32'd2818579584,	reg_addr : 32'd278646},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd278647},
'{step_type : POLL,	value : 32'd2147819648,	reg_addr : 32'd278648},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278649},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278650},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278651},
'{step_type : POLL,	value : 32'd2147820672,	reg_addr : 32'd278652},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278653},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278654},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278655},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd278656},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd278657},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd278658},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278659},
'{step_type : POLL,	value : 32'd3355457696,	reg_addr : 32'd278660},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278661},
'{step_type : POLL,	value : 32'd1409286289,	reg_addr : 32'd278662},
'{step_type : POLL,	value : 32'd102336,	reg_addr : 32'd278663},
'{step_type : POLL,	value : 32'd1409286289,	reg_addr : 32'd278664},
'{step_type : POLL,	value : 32'd85952,	reg_addr : 32'd278665},
'{step_type : POLL,	value : 32'd4026531985,	reg_addr : 32'd278666},
'{step_type : POLL,	value : 32'd100289,	reg_addr : 32'd278667},
'{step_type : POLL,	value : 32'd4026531985,	reg_addr : 32'd278668},
'{step_type : POLL,	value : 32'd83905,	reg_addr : 32'd278669},
'{step_type : POLL,	value : 32'd134219281,	reg_addr : 32'd278670},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd278671},
'{step_type : POLL,	value : 32'd80241,	reg_addr : 32'd278672},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278673},
'{step_type : POLL,	value : 32'd67111185,	reg_addr : 32'd278674},
'{step_type : POLL,	value : 32'd107552,	reg_addr : 32'd278675},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd278676},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278677},
'{step_type : POLL,	value : 32'd2577,	reg_addr : 32'd278678},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd278679},
'{step_type : POLL,	value : 32'd94545,	reg_addr : 32'd278680},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278681},
'{step_type : POLL,	value : 32'd82289,	reg_addr : 32'd278682},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278683},
'{step_type : POLL,	value : 32'd1553,	reg_addr : 32'd278684},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd278685},
'{step_type : POLL,	value : 32'd94577,	reg_addr : 32'd278686},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278687},
'{step_type : POLL,	value : 32'd603980945,	reg_addr : 32'd278688},
'{step_type : POLL,	value : 32'd123936,	reg_addr : 32'd278689},
'{step_type : POLL,	value : 32'd8657,	reg_addr : 32'd278690},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278691},
'{step_type : POLL,	value : 32'd4145,	reg_addr : 32'd278692},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278693},
'{step_type : POLL,	value : 32'd4145,	reg_addr : 32'd278694},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278695},
'{step_type : POLL,	value : 32'd11313,	reg_addr : 32'd278696},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278697},
'{step_type : POLL,	value : 32'd2818572433,	reg_addr : 32'd278698},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd278699},
'{step_type : POLL,	value : 32'd2147575953,	reg_addr : 32'd278700},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278701},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278702},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278703},
'{step_type : POLL,	value : 32'd2147576977,	reg_addr : 32'd278704},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278705},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278706},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278707},
'{step_type : POLL,	value : 32'd2129,	reg_addr : 32'd278708},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd278709},
'{step_type : POLL,	value : 32'd2147483793,	reg_addr : 32'd278710},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278711},
'{step_type : POLL,	value : 32'd2818572416,	reg_addr : 32'd278712},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278713},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278714},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278715},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278716},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278717},
'{step_type : POLL,	value : 32'd2818572416,	reg_addr : 32'd278718},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd278719},
'{step_type : POLL,	value : 32'd2147559552,	reg_addr : 32'd278720},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278721},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278722},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278723},
'{step_type : POLL,	value : 32'd2147560576,	reg_addr : 32'd278724},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278725},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278726},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278727},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd278728},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd278729},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd278730},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd278731},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278732},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278733},
'{step_type : POLL,	value : 32'd524800,	reg_addr : 32'd278734},
'{step_type : POLL,	value : 32'd16398,	reg_addr : 32'd278735},
'{step_type : POLL,	value : 32'd110912,	reg_addr : 32'd278736},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278737},
'{step_type : POLL,	value : 32'd131584,	reg_addr : 32'd278738},
'{step_type : POLL,	value : 32'd16398,	reg_addr : 32'd278739},
'{step_type : POLL,	value : 32'd110912,	reg_addr : 32'd278740},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278741},
'{step_type : POLL,	value : 32'd2147910144,	reg_addr : 32'd278742},
'{step_type : POLL,	value : 32'd16399,	reg_addr : 32'd278743},
'{step_type : POLL,	value : 32'd805309632,	reg_addr : 32'd278744},
'{step_type : POLL,	value : 32'd1988,	reg_addr : 32'd278745},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278746},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278747},
'{step_type : POLL,	value : 32'd1050112,	reg_addr : 32'd278748},
'{step_type : POLL,	value : 32'd16,	reg_addr : 32'd278749},
'{step_type : POLL,	value : 32'd738198720,	reg_addr : 32'd278750},
'{step_type : POLL,	value : 32'd960,	reg_addr : 32'd278751},
'{step_type : POLL,	value : 32'd2348820640,	reg_addr : 32'd278752},
'{step_type : POLL,	value : 32'd97217,	reg_addr : 32'd278753},
'{step_type : POLL,	value : 32'd2684355712,	reg_addr : 32'd278754},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd278755},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278756},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278757},
'{step_type : POLL,	value : 32'd2348815520,	reg_addr : 32'd278758},
'{step_type : POLL,	value : 32'd82881,	reg_addr : 32'd278759},
'{step_type : POLL,	value : 32'd2684354688,	reg_addr : 32'd278760},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd278761},
'{step_type : POLL,	value : 32'd2013267072,	reg_addr : 32'd278762},
'{step_type : POLL,	value : 32'd984,	reg_addr : 32'd278763},
'{step_type : POLL,	value : 32'd2080375936,	reg_addr : 32'd278764},
'{step_type : POLL,	value : 32'd2040,	reg_addr : 32'd278765},
'{step_type : POLL,	value : 32'd134217856,	reg_addr : 32'd278766},
'{step_type : POLL,	value : 32'd4064,	reg_addr : 32'd278767},
'{step_type : POLL,	value : 32'd134217856,	reg_addr : 32'd278768},
'{step_type : POLL,	value : 32'd2016,	reg_addr : 32'd278769},
'{step_type : POLL,	value : 32'd525824,	reg_addr : 32'd278770},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd278771},
'{step_type : POLL,	value : 32'd1216,	reg_addr : 32'd278772},
'{step_type : POLL,	value : 32'd85956,	reg_addr : 32'd278773},
'{step_type : POLL,	value : 32'd1216,	reg_addr : 32'd278774},
'{step_type : POLL,	value : 32'd83908,	reg_addr : 32'd278775},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd278776},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278777},
'{step_type : POLL,	value : 32'd134218880,	reg_addr : 32'd278778},
'{step_type : POLL,	value : 32'd4064,	reg_addr : 32'd278779},
'{step_type : POLL,	value : 32'd134218880,	reg_addr : 32'd278780},
'{step_type : POLL,	value : 32'd2016,	reg_addr : 32'd278781},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd278782},
'{step_type : POLL,	value : 32'd85956,	reg_addr : 32'd278783},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd278784},
'{step_type : POLL,	value : 32'd83908,	reg_addr : 32'd278785},
'{step_type : POLL,	value : 32'd2013266048,	reg_addr : 32'd278786},
'{step_type : POLL,	value : 32'd984,	reg_addr : 32'd278787},
'{step_type : POLL,	value : 32'd2080374912,	reg_addr : 32'd278788},
'{step_type : POLL,	value : 32'd2040,	reg_addr : 32'd278789},
'{step_type : POLL,	value : 32'd2348821664,	reg_addr : 32'd278790},
'{step_type : POLL,	value : 32'd97217,	reg_addr : 32'd278791},
'{step_type : POLL,	value : 32'd2684355712,	reg_addr : 32'd278792},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd278793},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278794},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278795},
'{step_type : POLL,	value : 32'd2348816544,	reg_addr : 32'd278796},
'{step_type : POLL,	value : 32'd82881,	reg_addr : 32'd278797},
'{step_type : POLL,	value : 32'd2684354688,	reg_addr : 32'd278798},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd278799},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd278800},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278801},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd278802},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd278803},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd278804},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd278805},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd278806},
'{step_type : POLL,	value : 32'd192,	reg_addr : 32'd278807},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd278808},
'{step_type : POLL,	value : 32'd256,	reg_addr : 32'd278809},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd278810},
'{step_type : POLL,	value : 32'd320,	reg_addr : 32'd278811},
'{step_type : POLL,	value : 32'd2098688,	reg_addr : 32'd278812},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd278813},
'{step_type : POLL,	value : 32'd738197696,	reg_addr : 32'd278814},
'{step_type : POLL,	value : 32'd448,	reg_addr : 32'd278815},
'{step_type : POLL,	value : 32'd738197696,	reg_addr : 32'd278816},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd278817},
'{step_type : POLL,	value : 32'd738197696,	reg_addr : 32'd278818},
'{step_type : POLL,	value : 32'd576,	reg_addr : 32'd278819},
'{step_type : POLL,	value : 32'd738197696,	reg_addr : 32'd278820},
'{step_type : POLL,	value : 32'd640,	reg_addr : 32'd278821},
'{step_type : POLL,	value : 32'd738197696,	reg_addr : 32'd278822},
'{step_type : POLL,	value : 32'd704,	reg_addr : 32'd278823},
'{step_type : POLL,	value : 32'd738197696,	reg_addr : 32'd278824},
'{step_type : POLL,	value : 32'd768,	reg_addr : 32'd278825},
'{step_type : POLL,	value : 32'd3288336512,	reg_addr : 32'd278826},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd278827},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278828},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278829},
'{step_type : POLL,	value : 32'd201327744,	reg_addr : 32'd278830},
'{step_type : POLL,	value : 32'd4036,	reg_addr : 32'd278831},
'{step_type : POLL,	value : 32'd67117056,	reg_addr : 32'd278832},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278833},
'{step_type : POLL,	value : 32'd201327744,	reg_addr : 32'd278834},
'{step_type : POLL,	value : 32'd1988,	reg_addr : 32'd278835},
'{step_type : POLL,	value : 32'd67117056,	reg_addr : 32'd278836},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278837},
'{step_type : POLL,	value : 32'd201326720,	reg_addr : 32'd278838},
'{step_type : POLL,	value : 32'd4036,	reg_addr : 32'd278839},
'{step_type : POLL,	value : 32'd201326720,	reg_addr : 32'd278840},
'{step_type : POLL,	value : 32'd1988,	reg_addr : 32'd278841},
'{step_type : POLL,	value : 32'd3288334464,	reg_addr : 32'd278842},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd278843},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278844},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278845},
'{step_type : POLL,	value : 32'd3758097536,	reg_addr : 32'd278846},
'{step_type : POLL,	value : 32'd2051,	reg_addr : 32'd278847},
'{step_type : POLL,	value : 32'd67117056,	reg_addr : 32'd278848},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278849},
'{step_type : POLL,	value : 32'd67110400,	reg_addr : 32'd278850},
'{step_type : POLL,	value : 32'd1024,	reg_addr : 32'd278851},
'{step_type : POLL,	value : 32'd643455168,	reg_addr : 32'd278852},
'{step_type : POLL,	value : 32'd100296,	reg_addr : 32'd278853},
'{step_type : POLL,	value : 32'd1476395136,	reg_addr : 32'd278854},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd278855},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278856},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278857},
'{step_type : POLL,	value : 32'd3758096512,	reg_addr : 32'd278858},
'{step_type : POLL,	value : 32'd2051,	reg_addr : 32'd278859},
'{step_type : POLL,	value : 32'd67117056,	reg_addr : 32'd278860},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278861},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278862},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278863},
'{step_type : POLL,	value : 32'd1342177408,	reg_addr : 32'd278864},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278865},
'{step_type : POLL,	value : 32'd1073742976,	reg_addr : 32'd278866},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd278867},
'{step_type : POLL,	value : 32'd3288334464,	reg_addr : 32'd278868},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd278869},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd278870},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd278871},
'{step_type : POLL,	value : 32'd2350907520,	reg_addr : 32'd278872},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd278873},
'{step_type : POLL,	value : 32'd2098688,	reg_addr : 32'd278874},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd278875},
'{step_type : POLL,	value : 32'd2282487936,	reg_addr : 32'd278876},
'{step_type : POLL,	value : 32'd3074,	reg_addr : 32'd278877},
'{step_type : POLL,	value : 32'd2282488000,	reg_addr : 32'd278878},
'{step_type : POLL,	value : 32'd3138,	reg_addr : 32'd278879},
'{step_type : POLL,	value : 32'd612367488,	reg_addr : 32'd278880},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd278881},
'{step_type : POLL,	value : 32'd673184896,	reg_addr : 32'd278882},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd278883},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278884},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278885},
'{step_type : POLL,	value : 32'd2148270208,	reg_addr : 32'd278886},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd278887},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278888},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278889},
'{step_type : POLL,	value : 32'd2550137984,	reg_addr : 32'd278890},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd278891},
'{step_type : POLL,	value : 32'd671089792,	reg_addr : 32'd278892},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd278893},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd278894},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278895},
'{step_type : POLL,	value : 32'd2164259968,	reg_addr : 32'd278896},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd278897},
'{step_type : POLL,	value : 32'd805306496,	reg_addr : 32'd278898},
'{step_type : POLL,	value : 32'd1988,	reg_addr : 32'd278899},
'{step_type : POLL,	value : 32'd67072,	reg_addr : 32'd278900},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd278901},
'{step_type : POLL,	value : 32'd194880,	reg_addr : 32'd278902},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278903},
'{step_type : POLL,	value : 32'd2147910144,	reg_addr : 32'd278904},
'{step_type : POLL,	value : 32'd16399,	reg_addr : 32'd278905},
'{step_type : POLL,	value : 32'd195936,	reg_addr : 32'd278906},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278907},
'{step_type : POLL,	value : 32'd105920,	reg_addr : 32'd278908},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278909},
'{step_type : POLL,	value : 32'd3758097536,	reg_addr : 32'd278910},
'{step_type : POLL,	value : 32'd2051,	reg_addr : 32'd278911},
'{step_type : POLL,	value : 32'd67116032,	reg_addr : 32'd278912},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278913},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd278914},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd278915},
'{step_type : POLL,	value : 32'd2281702528,	reg_addr : 32'd278916},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd278917},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd278918},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278919},
'{step_type : POLL,	value : 32'd1543504000,	reg_addr : 32'd278920},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd278921},
'{step_type : POLL,	value : 32'd33555968,	reg_addr : 32'd278922},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd278923},
'{step_type : POLL,	value : 32'd738201792,	reg_addr : 32'd278924},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd278925},
'{step_type : POLL,	value : 32'd738203776,	reg_addr : 32'd278926},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd278927},
'{step_type : POLL,	value : 32'd402659456,	reg_addr : 32'd278928},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd278929},
'{step_type : POLL,	value : 32'd469768320,	reg_addr : 32'd278930},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd278931},
'{step_type : POLL,	value : 32'd536877184,	reg_addr : 32'd278932},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd278933},
'{step_type : POLL,	value : 32'd603986048,	reg_addr : 32'd278934},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd278935},
'{step_type : POLL,	value : 32'd671094912,	reg_addr : 32'd278936},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd278937},
'{step_type : POLL,	value : 32'd131584,	reg_addr : 32'd278938},
'{step_type : POLL,	value : 32'd16398,	reg_addr : 32'd278939},
'{step_type : POLL,	value : 32'd223552,	reg_addr : 32'd278940},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278941},
'{step_type : POLL,	value : 32'd1073759744,	reg_addr : 32'd278942},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278943},
'{step_type : POLL,	value : 32'd218432,	reg_addr : 32'd278944},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278945},
'{step_type : POLL,	value : 32'd67111168,	reg_addr : 32'd278946},
'{step_type : POLL,	value : 32'd107552,	reg_addr : 32'd278947},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd278948},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278949},
'{step_type : POLL,	value : 32'd1073760768,	reg_addr : 32'd278950},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278951},
'{step_type : POLL,	value : 32'd201330912,	reg_addr : 32'd278952},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd278953},
'{step_type : POLL,	value : 32'd201326784,	reg_addr : 32'd278954},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd278955},
'{step_type : POLL,	value : 32'd67110016,	reg_addr : 32'd278956},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd278957},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278958},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278959},
'{step_type : POLL,	value : 32'd134218880,	reg_addr : 32'd278960},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd278961},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd278962},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278963},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278964},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278965},
'{step_type : POLL,	value : 32'd2617248945,	reg_addr : 32'd278966},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278967},
'{step_type : POLL,	value : 32'd2617249969,	reg_addr : 32'd278968},
'{step_type : POLL,	value : 32'd7171,	reg_addr : 32'd278969},
'{step_type : POLL,	value : 32'd603979921,	reg_addr : 32'd278970},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278971},
'{step_type : POLL,	value : 32'd81,	reg_addr : 32'd278972},
'{step_type : POLL,	value : 32'd16384,	reg_addr : 32'd278973},
'{step_type : POLL,	value : 32'd233777,	reg_addr : 32'd278974},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278975},
'{step_type : POLL,	value : 32'd1073748481,	reg_addr : 32'd278976},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278977},
'{step_type : POLL,	value : 32'd233825,	reg_addr : 32'd278978},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278979},
'{step_type : POLL,	value : 32'd603979905,	reg_addr : 32'd278980},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd278981},
'{step_type : POLL,	value : 32'd65,	reg_addr : 32'd278982},
'{step_type : POLL,	value : 32'd16384,	reg_addr : 32'd278983},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278984},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278985},
'{step_type : POLL,	value : 32'd2214594816,	reg_addr : 32'd278986},
'{step_type : POLL,	value : 32'd9244,	reg_addr : 32'd278987},
'{step_type : POLL,	value : 32'd3221307904,	reg_addr : 32'd278988},
'{step_type : POLL,	value : 32'd49153,	reg_addr : 32'd278989},
'{step_type : POLL,	value : 32'd239936,	reg_addr : 32'd278990},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278991},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd278992},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278993},
'{step_type : POLL,	value : 32'd738199712,	reg_addr : 32'd278994},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd278995},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd278996},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd278997},
'{step_type : POLL,	value : 32'd1073742976,	reg_addr : 32'd278998},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd278999},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279000},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279001},
'{step_type : POLL,	value : 32'd67108992,	reg_addr : 32'd279002},
'{step_type : POLL,	value : 32'd11264,	reg_addr : 32'd279003},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279004},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279005},
'{step_type : POLL,	value : 32'd131584,	reg_addr : 32'd279006},
'{step_type : POLL,	value : 32'd16398,	reg_addr : 32'd279007},
'{step_type : POLL,	value : 32'd278848,	reg_addr : 32'd279008},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279009},
'{step_type : POLL,	value : 32'd1073759744,	reg_addr : 32'd279010},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279011},
'{step_type : POLL,	value : 32'd67110080,	reg_addr : 32'd279012},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279013},
'{step_type : POLL,	value : 32'd134218944,	reg_addr : 32'd279014},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279015},
'{step_type : POLL,	value : 32'd278848,	reg_addr : 32'd279016},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279017},
'{step_type : POLL,	value : 32'd134217856,	reg_addr : 32'd279018},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279019},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279020},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279021},
'{step_type : POLL,	value : 32'd67108992,	reg_addr : 32'd279022},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279023},
'{step_type : POLL,	value : 32'd129,	reg_addr : 32'd279024},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279025},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279026},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279027},
'{step_type : POLL,	value : 32'd2281702528,	reg_addr : 32'd279028},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279029},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279030},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279031},
'{step_type : POLL,	value : 32'd201328896,	reg_addr : 32'd279032},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279033},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279034},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279035},
'{step_type : POLL,	value : 32'd68096,	reg_addr : 32'd279036},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd279037},
'{step_type : POLL,	value : 32'd269632,	reg_addr : 32'd279038},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279039},
'{step_type : POLL,	value : 32'd201329792,	reg_addr : 32'd279040},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279041},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd279042},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279043},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd279044},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279045},
'{step_type : POLL,	value : 32'd201328768,	reg_addr : 32'd279046},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279047},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd279048},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279049},
'{step_type : POLL,	value : 32'd201326720,	reg_addr : 32'd279050},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279051},
'{step_type : POLL,	value : 32'd279840,	reg_addr : 32'd279052},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279053},
'{step_type : POLL,	value : 32'd201333888,	reg_addr : 32'd279054},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279055},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd279056},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279057},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd279058},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279059},
'{step_type : POLL,	value : 32'd201332864,	reg_addr : 32'd279060},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279061},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd279062},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279063},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd279064},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279065},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd279066},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279067},
'{step_type : POLL,	value : 32'd201330816,	reg_addr : 32'd279068},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279069},
'{step_type : POLL,	value : 32'd279840,	reg_addr : 32'd279070},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279071},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd279072},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279073},
'{step_type : POLL,	value : 32'd2098688,	reg_addr : 32'd279074},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd279075},
'{step_type : POLL,	value : 32'd302432,	reg_addr : 32'd279076},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279077},
'{step_type : POLL,	value : 32'd402653312,	reg_addr : 32'd279078},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279079},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279080},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279081},
'{step_type : POLL,	value : 32'd536871040,	reg_addr : 32'd279082},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279083},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279084},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279085},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279086},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279087},
'{step_type : POLL,	value : 32'd738199680,	reg_addr : 32'd279088},
'{step_type : POLL,	value : 32'd14337,	reg_addr : 32'd279089},
'{step_type : POLL,	value : 32'd738201728,	reg_addr : 32'd279090},
'{step_type : POLL,	value : 32'd14401,	reg_addr : 32'd279091},
'{step_type : POLL,	value : 32'd738199680,	reg_addr : 32'd279092},
'{step_type : POLL,	value : 32'd14465,	reg_addr : 32'd279093},
'{step_type : POLL,	value : 32'd738201728,	reg_addr : 32'd279094},
'{step_type : POLL,	value : 32'd14529,	reg_addr : 32'd279095},
'{step_type : POLL,	value : 32'd738199680,	reg_addr : 32'd279096},
'{step_type : POLL,	value : 32'd14593,	reg_addr : 32'd279097},
'{step_type : POLL,	value : 32'd738201728,	reg_addr : 32'd279098},
'{step_type : POLL,	value : 32'd14657,	reg_addr : 32'd279099},
'{step_type : POLL,	value : 32'd738199680,	reg_addr : 32'd279100},
'{step_type : POLL,	value : 32'd14721,	reg_addr : 32'd279101},
'{step_type : POLL,	value : 32'd738201728,	reg_addr : 32'd279102},
'{step_type : POLL,	value : 32'd14785,	reg_addr : 32'd279103},
'{step_type : POLL,	value : 32'd33555968,	reg_addr : 32'd279104},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd279105},
'{step_type : POLL,	value : 32'd738201792,	reg_addr : 32'd279106},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279107},
'{step_type : POLL,	value : 32'd1476395136,	reg_addr : 32'd279108},
'{step_type : POLL,	value : 32'd975,	reg_addr : 32'd279109},
'{step_type : POLL,	value : 32'd1543504000,	reg_addr : 32'd279110},
'{step_type : POLL,	value : 32'd975,	reg_addr : 32'd279111},
'{step_type : POLL,	value : 32'd1543506048,	reg_addr : 32'd279112},
'{step_type : POLL,	value : 32'd207,	reg_addr : 32'd279113},
'{step_type : POLL,	value : 32'd1543506048,	reg_addr : 32'd279114},
'{step_type : POLL,	value : 32'd655,	reg_addr : 32'd279115},
'{step_type : POLL,	value : 32'd338208,	reg_addr : 32'd279116},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279117},
'{step_type : POLL,	value : 32'd402653312,	reg_addr : 32'd279118},
'{step_type : POLL,	value : 32'd14337,	reg_addr : 32'd279119},
'{step_type : POLL,	value : 32'd402653312,	reg_addr : 32'd279120},
'{step_type : POLL,	value : 32'd14401,	reg_addr : 32'd279121},
'{step_type : POLL,	value : 32'd402653312,	reg_addr : 32'd279122},
'{step_type : POLL,	value : 32'd14465,	reg_addr : 32'd279123},
'{step_type : POLL,	value : 32'd402653312,	reg_addr : 32'd279124},
'{step_type : POLL,	value : 32'd14529,	reg_addr : 32'd279125},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279126},
'{step_type : POLL,	value : 32'd14337,	reg_addr : 32'd279127},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279128},
'{step_type : POLL,	value : 32'd14401,	reg_addr : 32'd279129},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279130},
'{step_type : POLL,	value : 32'd14465,	reg_addr : 32'd279131},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279132},
'{step_type : POLL,	value : 32'd14529,	reg_addr : 32'd279133},
'{step_type : POLL,	value : 32'd536871040,	reg_addr : 32'd279134},
'{step_type : POLL,	value : 32'd14337,	reg_addr : 32'd279135},
'{step_type : POLL,	value : 32'd536871040,	reg_addr : 32'd279136},
'{step_type : POLL,	value : 32'd14401,	reg_addr : 32'd279137},
'{step_type : POLL,	value : 32'd536871040,	reg_addr : 32'd279138},
'{step_type : POLL,	value : 32'd14465,	reg_addr : 32'd279139},
'{step_type : POLL,	value : 32'd536871040,	reg_addr : 32'd279140},
'{step_type : POLL,	value : 32'd14529,	reg_addr : 32'd279141},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279142},
'{step_type : POLL,	value : 32'd14337,	reg_addr : 32'd279143},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279144},
'{step_type : POLL,	value : 32'd14401,	reg_addr : 32'd279145},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279146},
'{step_type : POLL,	value : 32'd14465,	reg_addr : 32'd279147},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279148},
'{step_type : POLL,	value : 32'd14529,	reg_addr : 32'd279149},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279150},
'{step_type : POLL,	value : 32'd14401,	reg_addr : 32'd279151},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279152},
'{step_type : POLL,	value : 32'd14529,	reg_addr : 32'd279153},
'{step_type : POLL,	value : 32'd738199680,	reg_addr : 32'd279154},
'{step_type : POLL,	value : 32'd14337,	reg_addr : 32'd279155},
'{step_type : POLL,	value : 32'd738201728,	reg_addr : 32'd279156},
'{step_type : POLL,	value : 32'd14401,	reg_addr : 32'd279157},
'{step_type : POLL,	value : 32'd738199680,	reg_addr : 32'd279158},
'{step_type : POLL,	value : 32'd14465,	reg_addr : 32'd279159},
'{step_type : POLL,	value : 32'd738201728,	reg_addr : 32'd279160},
'{step_type : POLL,	value : 32'd14529,	reg_addr : 32'd279161},
'{step_type : POLL,	value : 32'd33555968,	reg_addr : 32'd279162},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd279163},
'{step_type : POLL,	value : 32'd738201792,	reg_addr : 32'd279164},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279165},
'{step_type : POLL,	value : 32'd1476395136,	reg_addr : 32'd279166},
'{step_type : POLL,	value : 32'd15,	reg_addr : 32'd279167},
'{step_type : POLL,	value : 32'd1543504000,	reg_addr : 32'd279168},
'{step_type : POLL,	value : 32'd15,	reg_addr : 32'd279169},
'{step_type : POLL,	value : 32'd1476395136,	reg_addr : 32'd279170},
'{step_type : POLL,	value : 32'd79,	reg_addr : 32'd279171},
'{step_type : POLL,	value : 32'd1543504000,	reg_addr : 32'd279172},
'{step_type : POLL,	value : 32'd79,	reg_addr : 32'd279173},
'{step_type : POLL,	value : 32'd1476395136,	reg_addr : 32'd279174},
'{step_type : POLL,	value : 32'd143,	reg_addr : 32'd279175},
'{step_type : POLL,	value : 32'd1543504000,	reg_addr : 32'd279176},
'{step_type : POLL,	value : 32'd143,	reg_addr : 32'd279177},
'{step_type : POLL,	value : 32'd1476395136,	reg_addr : 32'd279178},
'{step_type : POLL,	value : 32'd207,	reg_addr : 32'd279179},
'{step_type : POLL,	value : 32'd1476395136,	reg_addr : 32'd279180},
'{step_type : POLL,	value : 32'd271,	reg_addr : 32'd279181},
'{step_type : POLL,	value : 32'd1543504000,	reg_addr : 32'd279182},
'{step_type : POLL,	value : 32'd271,	reg_addr : 32'd279183},
'{step_type : POLL,	value : 32'd1476395136,	reg_addr : 32'd279184},
'{step_type : POLL,	value : 32'd335,	reg_addr : 32'd279185},
'{step_type : POLL,	value : 32'd1543504000,	reg_addr : 32'd279186},
'{step_type : POLL,	value : 32'd335,	reg_addr : 32'd279187},
'{step_type : POLL,	value : 32'd536871040,	reg_addr : 32'd279188},
'{step_type : POLL,	value : 32'd11212,	reg_addr : 32'd279189},
'{step_type : POLL,	value : 32'd342321,	reg_addr : 32'd279190},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279191},
'{step_type : POLL,	value : 32'd1073748480,	reg_addr : 32'd279192},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279193},
'{step_type : POLL,	value : 32'd342368,	reg_addr : 32'd279194},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279195},
'{step_type : POLL,	value : 32'd67121312,	reg_addr : 32'd279196},
'{step_type : POLL,	value : 32'd11264,	reg_addr : 32'd279197},
'{step_type : POLL,	value : 32'd2281701504,	reg_addr : 32'd279198},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279199},
'{step_type : POLL,	value : 32'd1545600128,	reg_addr : 32'd279200},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279201},
'{step_type : POLL,	value : 32'd8390144,	reg_addr : 32'd279202},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd279203},
'{step_type : POLL,	value : 32'd3154118912,	reg_addr : 32'd279204},
'{step_type : POLL,	value : 32'd93196,	reg_addr : 32'd279205},
'{step_type : POLL,	value : 32'd67109056,	reg_addr : 32'd279206},
'{step_type : POLL,	value : 32'd9252,	reg_addr : 32'd279207},
'{step_type : POLL,	value : 32'd67141856,	reg_addr : 32'd279208},
'{step_type : POLL,	value : 32'd9252,	reg_addr : 32'd279209},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd279210},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279211},
'{step_type : POLL,	value : 32'd2550144181,	reg_addr : 32'd279212},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279213},
'{step_type : POLL,	value : 32'd2617254069,	reg_addr : 32'd279214},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279215},
'{step_type : POLL,	value : 32'd2550136981,	reg_addr : 32'd279216},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279217},
'{step_type : POLL,	value : 32'd2617245845,	reg_addr : 32'd279218},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279219},
'{step_type : POLL,	value : 32'd1073741973,	reg_addr : 32'd279220},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279221},
'{step_type : POLL,	value : 32'd1541,	reg_addr : 32'd279222},
'{step_type : POLL,	value : 32'd8192,	reg_addr : 32'd279223},
'{step_type : POLL,	value : 32'd1073742021,	reg_addr : 32'd279224},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279225},
'{step_type : POLL,	value : 32'd2147484869,	reg_addr : 32'd279226},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279227},
'{step_type : POLL,	value : 32'd2147483845,	reg_addr : 32'd279228},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279229},
'{step_type : POLL,	value : 32'd67109093,	reg_addr : 32'd279230},
'{step_type : POLL,	value : 32'd11264,	reg_addr : 32'd279231},
'{step_type : POLL,	value : 32'd3154116837,	reg_addr : 32'd279232},
'{step_type : POLL,	value : 32'd93196,	reg_addr : 32'd279233},
'{step_type : POLL,	value : 32'd67108864,	reg_addr : 32'd279234},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279235},
'{step_type : POLL,	value : 32'd2617115877,	reg_addr : 32'd279236},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279237},
'{step_type : POLL,	value : 32'd2684224741,	reg_addr : 32'd279238},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279239},
'{step_type : POLL,	value : 32'd2617114853,	reg_addr : 32'd279240},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279241},
'{step_type : POLL,	value : 32'd2684223717,	reg_addr : 32'd279242},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279243},
'{step_type : POLL,	value : 32'd1073743077,	reg_addr : 32'd279244},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279245},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279246},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279247},
'{step_type : POLL,	value : 32'd3154118821,	reg_addr : 32'd279248},
'{step_type : POLL,	value : 32'd93196,	reg_addr : 32'd279249},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd279250},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279251},
'{step_type : POLL,	value : 32'd3892513920,	reg_addr : 32'd279252},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279253},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279254},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279255},
'{step_type : POLL,	value : 32'd3892314240,	reg_addr : 32'd279256},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279257},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd279258},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279259},
'{step_type : POLL,	value : 32'd2281701504,	reg_addr : 32'd279260},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279261},
'{step_type : POLL,	value : 32'd67111936,	reg_addr : 32'd279262},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279263},
'{step_type : POLL,	value : 32'd52352,	reg_addr : 32'd279264},
'{step_type : POLL,	value : 32'd2056,	reg_addr : 32'd279265},
'{step_type : POLL,	value : 32'd469763200,	reg_addr : 32'd279266},
'{step_type : POLL,	value : 32'd4033,	reg_addr : 32'd279267},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279268},
'{step_type : POLL,	value : 32'd4033,	reg_addr : 32'd279269},
'{step_type : POLL,	value : 32'd469763200,	reg_addr : 32'd279270},
'{step_type : POLL,	value : 32'd1985,	reg_addr : 32'd279271},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279272},
'{step_type : POLL,	value : 32'd1985,	reg_addr : 32'd279273},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd279274},
'{step_type : POLL,	value : 32'd2056,	reg_addr : 32'd279275},
'{step_type : POLL,	value : 32'd1342177408,	reg_addr : 32'd279276},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279277},
'{step_type : POLL,	value : 32'd3087008896,	reg_addr : 32'd279278},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279279},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279280},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279281},
'{step_type : POLL,	value : 32'd263680,	reg_addr : 32'd279282},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd279283},
'{step_type : POLL,	value : 32'd1501561056,	reg_addr : 32'd279284},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd279285},
'{step_type : POLL,	value : 32'd671089792,	reg_addr : 32'd279286},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279287},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279288},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279289},
'{step_type : POLL,	value : 32'd3758096512,	reg_addr : 32'd279290},
'{step_type : POLL,	value : 32'd2051,	reg_addr : 32'd279291},
'{step_type : POLL,	value : 32'd67113984,	reg_addr : 32'd279292},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279293},
'{step_type : POLL,	value : 32'd2281703552,	reg_addr : 32'd279294},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279295},
'{step_type : POLL,	value : 32'd3104,	reg_addr : 32'd279296},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279297},
'{step_type : POLL,	value : 32'd1073759744,	reg_addr : 32'd279298},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279299},
'{step_type : POLL,	value : 32'd396640,	reg_addr : 32'd279300},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279301},
'{step_type : POLL,	value : 32'd469764224,	reg_addr : 32'd279302},
'{step_type : POLL,	value : 32'd4033,	reg_addr : 32'd279303},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279304},
'{step_type : POLL,	value : 32'd4033,	reg_addr : 32'd279305},
'{step_type : POLL,	value : 32'd469764224,	reg_addr : 32'd279306},
'{step_type : POLL,	value : 32'd1985,	reg_addr : 32'd279307},
'{step_type : POLL,	value : 32'd469762176,	reg_addr : 32'd279308},
'{step_type : POLL,	value : 32'd1985,	reg_addr : 32'd279309},
'{step_type : POLL,	value : 32'd67124224,	reg_addr : 32'd279310},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279311},
'{step_type : POLL,	value : 32'd263680,	reg_addr : 32'd279312},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd279313},
'{step_type : POLL,	value : 32'd404800,	reg_addr : 32'd279314},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279315},
'{step_type : POLL,	value : 32'd113088,	reg_addr : 32'd279316},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279317},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279318},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279319},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279320},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279321},
'{step_type : POLL,	value : 32'd2550136960,	reg_addr : 32'd279322},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279323},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279324},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279325},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279326},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279327},
'{step_type : POLL,	value : 32'd2285633664,	reg_addr : 32'd279328},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279329},
'{step_type : POLL,	value : 32'd2147746304,	reg_addr : 32'd279330},
'{step_type : POLL,	value : 32'd16399,	reg_addr : 32'd279331},
'{step_type : POLL,	value : 32'd419136,	reg_addr : 32'd279332},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279333},
'{step_type : POLL,	value : 32'd524800,	reg_addr : 32'd279334},
'{step_type : POLL,	value : 32'd16398,	reg_addr : 32'd279335},
'{step_type : POLL,	value : 32'd419136,	reg_addr : 32'd279336},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279337},
'{step_type : POLL,	value : 32'd3825206400,	reg_addr : 32'd279338},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279339},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279340},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279341},
'{step_type : POLL,	value : 32'd3825205376,	reg_addr : 32'd279342},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279343},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279344},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279345},
'{step_type : POLL,	value : 32'd3892513921,	reg_addr : 32'd279346},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279347},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279348},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279349},
'{step_type : POLL,	value : 32'd3892314241,	reg_addr : 32'd279350},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279351},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279352},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279353},
'{step_type : POLL,	value : 32'd1073748481,	reg_addr : 32'd279354},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279355},
'{step_type : POLL,	value : 32'd430401,	reg_addr : 32'd279356},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279357},
'{step_type : POLL,	value : 32'd2684355713,	reg_addr : 32'd279358},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd279359},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279360},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279361},
'{step_type : POLL,	value : 32'd1073754625,	reg_addr : 32'd279362},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279363},
'{step_type : POLL,	value : 32'd438593,	reg_addr : 32'd279364},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279365},
'{step_type : POLL,	value : 32'd430433,	reg_addr : 32'd279366},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279367},
'{step_type : POLL,	value : 32'd7201,	reg_addr : 32'd279368},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279369},
'{step_type : POLL,	value : 32'd2684354689,	reg_addr : 32'd279370},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd279371},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279372},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279373},
'{step_type : POLL,	value : 32'd132609,	reg_addr : 32'd279374},
'{step_type : POLL,	value : 32'd2,	reg_addr : 32'd279375},
'{step_type : POLL,	value : 32'd3892513985,	reg_addr : 32'd279376},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279377},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279378},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279379},
'{step_type : POLL,	value : 32'd3892314305,	reg_addr : 32'd279380},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279381},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279382},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279383},
'{step_type : POLL,	value : 32'd2684354689,	reg_addr : 32'd279384},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd279385},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279386},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279387},
'{step_type : POLL,	value : 32'd3892513937,	reg_addr : 32'd279388},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279389},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279390},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279391},
'{step_type : POLL,	value : 32'd3892314257,	reg_addr : 32'd279392},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279393},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279394},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279395},
'{step_type : POLL,	value : 32'd2818573440,	reg_addr : 32'd279396},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279397},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279398},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279399},
'{step_type : POLL,	value : 32'd402653313,	reg_addr : 32'd279400},
'{step_type : POLL,	value : 32'd123936,	reg_addr : 32'd279401},
'{step_type : POLL,	value : 32'd1073767953,	reg_addr : 32'd279402},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279403},
'{step_type : POLL,	value : 32'd450897,	reg_addr : 32'd279404},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279405},
'{step_type : POLL,	value : 32'd8657,	reg_addr : 32'd279406},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279407},
'{step_type : POLL,	value : 32'd2684355729,	reg_addr : 32'd279408},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd279409},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279410},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279411},
'{step_type : POLL,	value : 32'd1409294513,	reg_addr : 32'd279412},
'{step_type : POLL,	value : 32'd85952,	reg_addr : 32'd279413},
'{step_type : POLL,	value : 32'd4026541233,	reg_addr : 32'd279414},
'{step_type : POLL,	value : 32'd83905,	reg_addr : 32'd279415},
'{step_type : POLL,	value : 32'd2684354705,	reg_addr : 32'd279416},
'{step_type : POLL,	value : 32'd9248,	reg_addr : 32'd279417},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd279418},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279419},
'{step_type : POLL,	value : 32'd2818572416,	reg_addr : 32'd279420},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279421},
'{step_type : POLL,	value : 32'd2147561600,	reg_addr : 32'd279422},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279423},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279424},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279425},
'{step_type : POLL,	value : 32'd2147562624,	reg_addr : 32'd279426},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279427},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279428},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279429},
'{step_type : POLL,	value : 32'd67116032,	reg_addr : 32'd279430},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279431},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279432},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279433},
'{step_type : POLL,	value : 32'd1056,	reg_addr : 32'd279434},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279435},
'{step_type : POLL,	value : 32'd2818572416,	reg_addr : 32'd279436},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279437},
'{step_type : POLL,	value : 32'd2147563648,	reg_addr : 32'd279438},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279439},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279440},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279441},
'{step_type : POLL,	value : 32'd2147564672,	reg_addr : 32'd279442},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279443},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279444},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279445},
'{step_type : POLL,	value : 32'd67116032,	reg_addr : 32'd279446},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279447},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279448},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279449},
'{step_type : POLL,	value : 32'd1056,	reg_addr : 32'd279450},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279451},
'{step_type : POLL,	value : 32'd2818572416,	reg_addr : 32'd279452},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279453},
'{step_type : POLL,	value : 32'd2147565696,	reg_addr : 32'd279454},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279455},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279456},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279457},
'{step_type : POLL,	value : 32'd2147566720,	reg_addr : 32'd279458},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279459},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279460},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279461},
'{step_type : POLL,	value : 32'd67116032,	reg_addr : 32'd279462},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279463},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279464},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279465},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd279466},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279467},
'{step_type : POLL,	value : 32'd536871046,	reg_addr : 32'd279468},
'{step_type : POLL,	value : 32'd116676,	reg_addr : 32'd279469},
'{step_type : POLL,	value : 32'd2650801280,	reg_addr : 32'd279470},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279471},
'{step_type : POLL,	value : 32'd3288727680,	reg_addr : 32'd279472},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279473},
'{step_type : POLL,	value : 32'd3556770944,	reg_addr : 32'd279474},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279475},
'{step_type : POLL,	value : 32'd3825206400,	reg_addr : 32'd279476},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279477},
'{step_type : POLL,	value : 32'd2617258112,	reg_addr : 32'd279478},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279479},
'{step_type : POLL,	value : 32'd2080374912,	reg_addr : 32'd279480},
'{step_type : POLL,	value : 32'd116673,	reg_addr : 32'd279481},
'{step_type : POLL,	value : 32'd2281704576,	reg_addr : 32'd279482},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279483},
'{step_type : POLL,	value : 32'd1677724800,	reg_addr : 32'd279484},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279485},
'{step_type : POLL,	value : 32'd2415921280,	reg_addr : 32'd279486},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279487},
'{step_type : POLL,	value : 32'd3960470656,	reg_addr : 32'd279488},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279489},
'{step_type : POLL,	value : 32'd3959423104,	reg_addr : 32'd279490},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279491},
'{step_type : POLL,	value : 32'd4160749696,	reg_addr : 32'd279492},
'{step_type : POLL,	value : 32'd2046,	reg_addr : 32'd279493},
'{step_type : POLL,	value : 32'd4160750720,	reg_addr : 32'd279494},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279495},
'{step_type : POLL,	value : 32'd4160750720,	reg_addr : 32'd279496},
'{step_type : POLL,	value : 32'd2002,	reg_addr : 32'd279497},
'{step_type : POLL,	value : 32'd2818576512,	reg_addr : 32'd279498},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279499},
'{step_type : POLL,	value : 32'd2147567744,	reg_addr : 32'd279500},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279501},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279502},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279503},
'{step_type : POLL,	value : 32'd2147568768,	reg_addr : 32'd279504},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279505},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279506},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279507},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd279508},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd279509},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279510},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279511},
'{step_type : POLL,	value : 32'd4160749696,	reg_addr : 32'd279512},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279513},
'{step_type : POLL,	value : 32'd4160749696,	reg_addr : 32'd279514},
'{step_type : POLL,	value : 32'd2002,	reg_addr : 32'd279515},
'{step_type : POLL,	value : 32'd3960470656,	reg_addr : 32'd279516},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279517},
'{step_type : POLL,	value : 32'd3959423104,	reg_addr : 32'd279518},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279519},
'{step_type : POLL,	value : 32'd4160750720,	reg_addr : 32'd279520},
'{step_type : POLL,	value : 32'd1990,	reg_addr : 32'd279521},
'{step_type : POLL,	value : 32'd4160750720,	reg_addr : 32'd279522},
'{step_type : POLL,	value : 32'd2006,	reg_addr : 32'd279523},
'{step_type : POLL,	value : 32'd2818576512,	reg_addr : 32'd279524},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279525},
'{step_type : POLL,	value : 32'd2147569792,	reg_addr : 32'd279526},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279527},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279528},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279529},
'{step_type : POLL,	value : 32'd2147570816,	reg_addr : 32'd279530},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279531},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279532},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279533},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd279534},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd279535},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279536},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279537},
'{step_type : POLL,	value : 32'd4160749696,	reg_addr : 32'd279538},
'{step_type : POLL,	value : 32'd1990,	reg_addr : 32'd279539},
'{step_type : POLL,	value : 32'd4160749696,	reg_addr : 32'd279540},
'{step_type : POLL,	value : 32'd2006,	reg_addr : 32'd279541},
'{step_type : POLL,	value : 32'd1677723776,	reg_addr : 32'd279542},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279543},
'{step_type : POLL,	value : 32'd5152,	reg_addr : 32'd279544},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279545},
'{step_type : POLL,	value : 32'd3288335488,	reg_addr : 32'd279546},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd279547},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279548},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279549},
'{step_type : POLL,	value : 32'd3288334464,	reg_addr : 32'd279550},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd279551},
'{step_type : POLL,	value : 32'd67110400,	reg_addr : 32'd279552},
'{step_type : POLL,	value : 32'd1024,	reg_addr : 32'd279553},
'{step_type : POLL,	value : 32'd617138368,	reg_addr : 32'd279554},
'{step_type : POLL,	value : 32'd83912,	reg_addr : 32'd279555},
'{step_type : POLL,	value : 32'd2147484800,	reg_addr : 32'd279556},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279557},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279558},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279559},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279560},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279561},
'{step_type : POLL,	value : 32'd2415919232,	reg_addr : 32'd279562},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279563},
'{step_type : POLL,	value : 32'd2550140032,	reg_addr : 32'd279564},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279565},
'{step_type : POLL,	value : 32'd2818576512,	reg_addr : 32'd279566},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279567},
'{step_type : POLL,	value : 32'd2147571840,	reg_addr : 32'd279568},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279569},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279570},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279571},
'{step_type : POLL,	value : 32'd2147572864,	reg_addr : 32'd279572},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279573},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279574},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279575},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd279576},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd279577},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279578},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279579},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279580},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279581},
'{step_type : POLL,	value : 32'd2550136960,	reg_addr : 32'd279582},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279583},
'{step_type : POLL,	value : 32'd2281701504,	reg_addr : 32'd279584},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279585},
'{step_type : POLL,	value : 32'd1677721728,	reg_addr : 32'd279586},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279587},
'{step_type : POLL,	value : 32'd2080375936,	reg_addr : 32'd279588},
'{step_type : POLL,	value : 32'd116673,	reg_addr : 32'd279589},
'{step_type : POLL,	value : 32'd3825206400,	reg_addr : 32'd279590},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279591},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279592},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279593},
'{step_type : POLL,	value : 32'd3825205376,	reg_addr : 32'd279594},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279595},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279596},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279597},
'{step_type : POLL,	value : 32'd6176,	reg_addr : 32'd279598},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279599},
'{step_type : POLL,	value : 32'd2415920256,	reg_addr : 32'd279600},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279601},
'{step_type : POLL,	value : 32'd2818576512,	reg_addr : 32'd279602},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279603},
'{step_type : POLL,	value : 32'd2147573888,	reg_addr : 32'd279604},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279605},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279606},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279607},
'{step_type : POLL,	value : 32'd2147574912,	reg_addr : 32'd279608},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279609},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279610},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279611},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd279612},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd279613},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279614},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279615},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279616},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279617},
'{step_type : POLL,	value : 32'd2147484800,	reg_addr : 32'd279618},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279619},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279620},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279621},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279622},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279623},
'{step_type : POLL,	value : 32'd2415919232,	reg_addr : 32'd279624},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279625},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279626},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279627},
'{step_type : POLL,	value : 32'd3825206400,	reg_addr : 32'd279628},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279629},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279630},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279631},
'{step_type : POLL,	value : 32'd3825205376,	reg_addr : 32'd279632},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279633},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279634},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279635},
'{step_type : POLL,	value : 32'd2818572416,	reg_addr : 32'd279636},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279637},
'{step_type : POLL,	value : 32'd1342178432,	reg_addr : 32'd279638},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279639},
'{step_type : POLL,	value : 32'd536872070,	reg_addr : 32'd279640},
'{step_type : POLL,	value : 32'd116676,	reg_addr : 32'd279641},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd279642},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279643},
'{step_type : POLL,	value : 32'd2147517952,	reg_addr : 32'd279644},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279645},
'{step_type : POLL,	value : 32'd581984,	reg_addr : 32'd279646},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279647},
'{step_type : POLL,	value : 32'd2147484800,	reg_addr : 32'd279648},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279649},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279650},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279651},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279652},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279653},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279654},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279655},
'{step_type : POLL,	value : 32'd3825206400,	reg_addr : 32'd279656},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279657},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279658},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279659},
'{step_type : POLL,	value : 32'd3825205376,	reg_addr : 32'd279660},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279661},
'{step_type : POLL,	value : 32'd2818572416,	reg_addr : 32'd279662},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279663},
'{step_type : POLL,	value : 32'd3087007872,	reg_addr : 32'd279664},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279665},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279666},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279667},
'{step_type : POLL,	value : 32'd4224,	reg_addr : 32'd279668},
'{step_type : POLL,	value : 32'd13250,	reg_addr : 32'd279669},
'{step_type : POLL,	value : 32'd1342178432,	reg_addr : 32'd279670},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279671},
'{step_type : POLL,	value : 32'd3019899008,	reg_addr : 32'd279672},
'{step_type : POLL,	value : 32'd9216,	reg_addr : 32'd279673},
'{step_type : POLL,	value : 32'd2281702529,	reg_addr : 32'd279674},
'{step_type : POLL,	value : 32'd3072,	reg_addr : 32'd279675},
'{step_type : POLL,	value : 32'd603980928,	reg_addr : 32'd279676},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279677},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd279678},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279679},
'{step_type : POLL,	value : 32'd1073742976,	reg_addr : 32'd279680},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279681},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd279682},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279683},
'{step_type : POLL,	value : 32'd2348810368,	reg_addr : 32'd279684},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279685},
'{step_type : POLL,	value : 32'd2098688,	reg_addr : 32'd279686},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd279687},
'{step_type : POLL,	value : 32'd2282487936,	reg_addr : 32'd279688},
'{step_type : POLL,	value : 32'd3074,	reg_addr : 32'd279689},
'{step_type : POLL,	value : 32'd2282488000,	reg_addr : 32'd279690},
'{step_type : POLL,	value : 32'd3138,	reg_addr : 32'd279691},
'{step_type : POLL,	value : 32'd612367488,	reg_addr : 32'd279692},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279693},
'{step_type : POLL,	value : 32'd673184896,	reg_addr : 32'd279694},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279695},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279696},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279697},
'{step_type : POLL,	value : 32'd2550137984,	reg_addr : 32'd279698},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279699},
'{step_type : POLL,	value : 32'd671089792,	reg_addr : 32'd279700},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279701},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279702},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279703},
'{step_type : POLL,	value : 32'd2164259968,	reg_addr : 32'd279704},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279705},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279706},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279707},
'{step_type : POLL,	value : 32'd3758097536,	reg_addr : 32'd279708},
'{step_type : POLL,	value : 32'd2051,	reg_addr : 32'd279709},
'{step_type : POLL,	value : 32'd67117056,	reg_addr : 32'd279710},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279711},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279712},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279713},
'{step_type : POLL,	value : 32'd1342177408,	reg_addr : 32'd279714},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279715},
'{step_type : POLL,	value : 32'd1152,	reg_addr : 32'd279716},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279717},
'{step_type : POLL,	value : 32'd201326720,	reg_addr : 32'd279718},
'{step_type : POLL,	value : 32'd6144,	reg_addr : 32'd279719},
'{step_type : POLL,	value : 32'd1543504000,	reg_addr : 32'd279720},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279721},
'{step_type : POLL,	value : 32'd67108992,	reg_addr : 32'd279722},
'{step_type : POLL,	value : 32'd11264,	reg_addr : 32'd279723},
'{step_type : POLL,	value : 32'd33555968,	reg_addr : 32'd279724},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd279725},
'{step_type : POLL,	value : 32'd738201792,	reg_addr : 32'd279726},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279727},
'{step_type : POLL,	value : 32'd738203776,	reg_addr : 32'd279728},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279729},
'{step_type : POLL,	value : 32'd402659456,	reg_addr : 32'd279730},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279731},
'{step_type : POLL,	value : 32'd469768320,	reg_addr : 32'd279732},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279733},
'{step_type : POLL,	value : 32'd536877184,	reg_addr : 32'd279734},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279735},
'{step_type : POLL,	value : 32'd603986048,	reg_addr : 32'd279736},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279737},
'{step_type : POLL,	value : 32'd671094912,	reg_addr : 32'd279738},
'{step_type : POLL,	value : 32'd15297,	reg_addr : 32'd279739},
'{step_type : POLL,	value : 32'd536873088,	reg_addr : 32'd279740},
'{step_type : POLL,	value : 32'd11212,	reg_addr : 32'd279741},
'{step_type : POLL,	value : 32'd67121312,	reg_addr : 32'd279742},
'{step_type : POLL,	value : 32'd11264,	reg_addr : 32'd279743},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279744},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279745},
'{step_type : POLL,	value : 32'd3019900032,	reg_addr : 32'd279746},
'{step_type : POLL,	value : 32'd9216,	reg_addr : 32'd279747},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd279748},
'{step_type : POLL,	value : 32'd16384,	reg_addr : 32'd279749},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd279750},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279751},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd279752},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279753},
'{step_type : POLL,	value : 32'd2281704576,	reg_addr : 32'd279754},
'{step_type : POLL,	value : 32'd3072,	reg_addr : 32'd279755},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279756},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279757},
'{step_type : POLL,	value : 32'd67111936,	reg_addr : 32'd279758},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279759},
'{step_type : POLL,	value : 32'd2281702528,	reg_addr : 32'd279760},
'{step_type : POLL,	value : 32'd2050,	reg_addr : 32'd279761},
'{step_type : POLL,	value : 32'd480,	reg_addr : 32'd279762},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279763},
'{step_type : POLL,	value : 32'd6272,	reg_addr : 32'd279764},
'{step_type : POLL,	value : 32'd13250,	reg_addr : 32'd279765},
'{step_type : POLL,	value : 32'd2497,	reg_addr : 32'd279766},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279767},
'{step_type : POLL,	value : 32'd2617249041,	reg_addr : 32'd279768},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279769},
'{step_type : POLL,	value : 32'd67112977,	reg_addr : 32'd279770},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279771},
'{step_type : POLL,	value : 32'd2617250065,	reg_addr : 32'd279772},
'{step_type : POLL,	value : 32'd7171,	reg_addr : 32'd279773},
'{step_type : POLL,	value : 32'd67112977,	reg_addr : 32'd279774},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279775},
'{step_type : POLL,	value : 32'd2617245841,	reg_addr : 32'd279776},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279777},
'{step_type : POLL,	value : 32'd2617245841,	reg_addr : 32'd279778},
'{step_type : POLL,	value : 32'd7171,	reg_addr : 32'd279779},
'{step_type : POLL,	value : 32'd649505,	reg_addr : 32'd279780},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279781},
'{step_type : POLL,	value : 32'd3087008896,	reg_addr : 32'd279782},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279783},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279784},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279785},
'{step_type : POLL,	value : 32'd2147910144,	reg_addr : 32'd279786},
'{step_type : POLL,	value : 32'd16399,	reg_addr : 32'd279787},
'{step_type : POLL,	value : 32'd647488,	reg_addr : 32'd279788},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279789},
'{step_type : POLL,	value : 32'd36288,	reg_addr : 32'd279790},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279791},
'{step_type : POLL,	value : 32'd97728,	reg_addr : 32'd279792},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279793},
'{step_type : POLL,	value : 32'd172480,	reg_addr : 32'd279794},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279795},
'{step_type : POLL,	value : 32'd224704,	reg_addr : 32'd279796},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279797},
'{step_type : POLL,	value : 32'd234944,	reg_addr : 32'd279798},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279799},
'{step_type : POLL,	value : 32'd241088,	reg_addr : 32'd279800},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279801},
'{step_type : POLL,	value : 32'd375232,	reg_addr : 32'd279802},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279803},
'{step_type : POLL,	value : 32'd1610727552,	reg_addr : 32'd279804},
'{step_type : POLL,	value : 32'd9253,	reg_addr : 32'd279805},
'{step_type : POLL,	value : 32'd524800,	reg_addr : 32'd279806},
'{step_type : POLL,	value : 32'd16398,	reg_addr : 32'd279807},
'{step_type : POLL,	value : 32'd665920,	reg_addr : 32'd279808},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279809},
'{step_type : POLL,	value : 32'd658737,	reg_addr : 32'd279810},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279811},
'{step_type : POLL,	value : 32'd457152,	reg_addr : 32'd279812},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279813},
'{step_type : POLL,	value : 32'd2147517952,	reg_addr : 32'd279814},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279815},
'{step_type : POLL,	value : 32'd665920,	reg_addr : 32'd279816},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279817},
'{step_type : POLL,	value : 32'd481730,	reg_addr : 32'd279818},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279819},
'{step_type : POLL,	value : 32'd2147910144,	reg_addr : 32'd279820},
'{step_type : POLL,	value : 32'd16399,	reg_addr : 32'd279821},
'{step_type : POLL,	value : 32'd3288335552,	reg_addr : 32'd279822},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd279823},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279824},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279825},
'{step_type : POLL,	value : 32'd3288334528,	reg_addr : 32'd279826},
'{step_type : POLL,	value : 32'd1984,	reg_addr : 32'd279827},
'{step_type : POLL,	value : 32'd1073767953,	reg_addr : 32'd279828},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279829},
'{step_type : POLL,	value : 32'd684369,	reg_addr : 32'd279830},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279831},
'{step_type : POLL,	value : 32'd2147910161,	reg_addr : 32'd279832},
'{step_type : POLL,	value : 32'd16399,	reg_addr : 32'd279833},
'{step_type : POLL,	value : 32'd684369,	reg_addr : 32'd279834},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279835},
'{step_type : POLL,	value : 32'd524817,	reg_addr : 32'd279836},
'{step_type : POLL,	value : 32'd16398,	reg_addr : 32'd279837},
'{step_type : POLL,	value : 32'd674129,	reg_addr : 32'd279838},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279839},
'{step_type : POLL,	value : 32'd2147517969,	reg_addr : 32'd279840},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279841},
'{step_type : POLL,	value : 32'd677233,	reg_addr : 32'd279842},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279843},
'{step_type : POLL,	value : 32'd4145,	reg_addr : 32'd279844},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279845},
'{step_type : POLL,	value : 32'd4145,	reg_addr : 32'd279846},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279847},
'{step_type : POLL,	value : 32'd11313,	reg_addr : 32'd279848},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279849},
'{step_type : POLL,	value : 32'd2818572433,	reg_addr : 32'd279850},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279851},
'{step_type : POLL,	value : 32'd2147575953,	reg_addr : 32'd279852},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279853},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279854},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279855},
'{step_type : POLL,	value : 32'd2147576977,	reg_addr : 32'd279856},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279857},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279858},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279859},
'{step_type : POLL,	value : 32'd2129,	reg_addr : 32'd279860},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd279861},
'{step_type : POLL,	value : 32'd2147483793,	reg_addr : 32'd279862},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279863},
'{step_type : POLL,	value : 32'd603979921,	reg_addr : 32'd279864},
'{step_type : POLL,	value : 32'd123936,	reg_addr : 32'd279865},
'{step_type : POLL,	value : 32'd571840,	reg_addr : 32'd279866},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279867},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279868},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279869},
'{step_type : POLL,	value : 32'd590272,	reg_addr : 32'd279870},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279871},
'{step_type : POLL,	value : 32'd603980928,	reg_addr : 32'd279872},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279873},
'{step_type : POLL,	value : 32'd1024,	reg_addr : 32'd279874},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279875},
'{step_type : POLL,	value : 32'd1342177408,	reg_addr : 32'd279876},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279877},
'{step_type : POLL,	value : 32'd2617249024,	reg_addr : 32'd279878},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279879},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279880},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279881},
'{step_type : POLL,	value : 32'd2617250048,	reg_addr : 32'd279882},
'{step_type : POLL,	value : 32'd7171,	reg_addr : 32'd279883},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279884},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279885},
'{step_type : POLL,	value : 32'd2617245824,	reg_addr : 32'd279886},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279887},
'{step_type : POLL,	value : 32'd2617245824,	reg_addr : 32'd279888},
'{step_type : POLL,	value : 32'd7171,	reg_addr : 32'd279889},
'{step_type : POLL,	value : 32'd6272,	reg_addr : 32'd279890},
'{step_type : POLL,	value : 32'd13250,	reg_addr : 32'd279891},
'{step_type : POLL,	value : 32'd3087008896,	reg_addr : 32'd279892},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd279893},
'{step_type : POLL,	value : 32'd67111936,	reg_addr : 32'd279894},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279895},
'{step_type : POLL,	value : 32'd603980945,	reg_addr : 32'd279896},
'{step_type : POLL,	value : 32'd123936,	reg_addr : 32'd279897},
'{step_type : POLL,	value : 32'd2818572416,	reg_addr : 32'd279898},
'{step_type : POLL,	value : 32'd7174,	reg_addr : 32'd279899},
'{step_type : POLL,	value : 32'd2147559552,	reg_addr : 32'd279900},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279901},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279902},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279903},
'{step_type : POLL,	value : 32'd2147560576,	reg_addr : 32'd279904},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279905},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279906},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279907},
'{step_type : POLL,	value : 32'd2112,	reg_addr : 32'd279908},
'{step_type : POLL,	value : 32'd24576,	reg_addr : 32'd279909},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279910},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd279911},
'{step_type : POLL,	value : 32'd738197632,	reg_addr : 32'd279912},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279913},
'{step_type : POLL,	value : 32'd2350907520,	reg_addr : 32'd279914},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279915},
'{step_type : POLL,	value : 32'd2098688,	reg_addr : 32'd279916},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd279917},
'{step_type : POLL,	value : 32'd2285633664,	reg_addr : 32'd279918},
'{step_type : POLL,	value : 32'd3074,	reg_addr : 32'd279919},
'{step_type : POLL,	value : 32'd2285633728,	reg_addr : 32'd279920},
'{step_type : POLL,	value : 32'd3138,	reg_addr : 32'd279921},
'{step_type : POLL,	value : 32'd2550137984,	reg_addr : 32'd279922},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279923},
'{step_type : POLL,	value : 32'd671089792,	reg_addr : 32'd279924},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279925},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279926},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279927},
'{step_type : POLL,	value : 32'd2164259968,	reg_addr : 32'd279928},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279929},
'{step_type : POLL,	value : 32'd612367488,	reg_addr : 32'd279930},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279931},
'{step_type : POLL,	value : 32'd673184896,	reg_addr : 32'd279932},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279933},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd279934},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279935},
'{step_type : POLL,	value : 32'd3758097536,	reg_addr : 32'd279936},
'{step_type : POLL,	value : 32'd2051,	reg_addr : 32'd279937},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279938},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279939},
'{step_type : POLL,	value : 32'd8390144,	reg_addr : 32'd279940},
'{step_type : POLL,	value : 32'd128,	reg_addr : 32'd279941},
'{step_type : POLL,	value : 32'd67109056,	reg_addr : 32'd279942},
'{step_type : POLL,	value : 32'd9252,	reg_addr : 32'd279943},
'{step_type : POLL,	value : 32'd67141856,	reg_addr : 32'd279944},
'{step_type : POLL,	value : 32'd9252,	reg_addr : 32'd279945},
'{step_type : POLL,	value : 32'd1073743074,	reg_addr : 32'd279946},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279947},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279948},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279949},
'{step_type : POLL,	value : 32'd1073742050,	reg_addr : 32'd279950},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279951},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279952},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279953},
'{step_type : POLL,	value : 32'd2147484896,	reg_addr : 32'd279954},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279955},
'{step_type : POLL,	value : 32'd2147483872,	reg_addr : 32'd279956},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279957},
'{step_type : POLL,	value : 32'd1541,	reg_addr : 32'd279958},
'{step_type : POLL,	value : 32'd8192,	reg_addr : 32'd279959},
'{step_type : POLL,	value : 32'd1073743042,	reg_addr : 32'd279960},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279961},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279962},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279963},
'{step_type : POLL,	value : 32'd1073742018,	reg_addr : 32'd279964},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279965},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279966},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279967},
'{step_type : POLL,	value : 32'd2147484864,	reg_addr : 32'd279968},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279969},
'{step_type : POLL,	value : 32'd2147483840,	reg_addr : 32'd279970},
'{step_type : POLL,	value : 32'd11276,	reg_addr : 32'd279971},
'{step_type : POLL,	value : 32'd67111936,	reg_addr : 32'd279972},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279973},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279974},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd279975},
'{step_type : POLL,	value : 32'd268435968,	reg_addr : 32'd279976},
'{step_type : POLL,	value : 32'd20480,	reg_addr : 32'd279977},
'{step_type : POLL,	value : 32'd744768,	reg_addr : 32'd279978},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279979},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd279980},
'{step_type : POLL,	value : 32'd16384,	reg_addr : 32'd279981},
'{step_type : POLL,	value : 32'd671089792,	reg_addr : 32'd279982},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279983},
'{step_type : POLL,	value : 32'd67112960,	reg_addr : 32'd279984},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279985},
'{step_type : POLL,	value : 32'd3758096512,	reg_addr : 32'd279986},
'{step_type : POLL,	value : 32'd2051,	reg_addr : 32'd279987},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd279988},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd279989},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279990},
'{step_type : POLL,	value : 32'd4032,	reg_addr : 32'd279991},
'{step_type : POLL,	value : 32'd2147483776,	reg_addr : 32'd279992},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279993},
'{step_type : POLL,	value : 32'd2550136960,	reg_addr : 32'd279994},
'{step_type : POLL,	value : 32'd4034,	reg_addr : 32'd279995},
'{step_type : POLL,	value : 32'd603979904,	reg_addr : 32'd279996},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279997},
'{step_type : POLL,	value : 32'd671088768,	reg_addr : 32'd279998},
'{step_type : POLL,	value : 32'd1986,	reg_addr : 32'd279999},
'{step_type : POLL,	value : 32'd3825206400,	reg_addr : 32'd280000},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd280001},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd280002},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280003},
'{step_type : POLL,	value : 32'd3825205376,	reg_addr : 32'd280004},
'{step_type : POLL,	value : 32'd2049,	reg_addr : 32'd280005},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd280006},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280007},
'{step_type : POLL,	value : 32'd2818573440,	reg_addr : 32'd280008},
'{step_type : POLL,	value : 32'd7172,	reg_addr : 32'd280009},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd280010},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280011},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd280012},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280013},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd280014},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280015},
'{step_type : POLL,	value : 32'd4128,	reg_addr : 32'd280016},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280017},
'{step_type : POLL,	value : 32'd3892513920,	reg_addr : 32'd280018},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd280019},
'{step_type : POLL,	value : 32'd67110912,	reg_addr : 32'd280020},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280021},
'{step_type : POLL,	value : 32'd3892314240,	reg_addr : 32'd280022},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd280023},
'{step_type : POLL,	value : 32'd67109888,	reg_addr : 32'd280024},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280025},
'{step_type : POLL,	value : 32'd2617248928,	reg_addr : 32'd280026},
'{step_type : POLL,	value : 32'd7169,	reg_addr : 32'd280027},
'{step_type : POLL,	value : 32'd2617249952,	reg_addr : 32'd280028},
'{step_type : POLL,	value : 32'd7171,	reg_addr : 32'd280029},
'{step_type : POLL,	value : 32'd658720,	reg_addr : 32'd280030},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd280031},
'{step_type : POLL,	value : 32'd1024,	reg_addr : 32'd852199},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459146},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd459556},
'{step_type : POLL,	value : 32'd25,	reg_addr : 32'd459557},
'{step_type : POLL,	value : 32'd46,	reg_addr : 32'd459558},
'{step_type : POLL,	value : 32'd67,	reg_addr : 32'd459559},
'{step_type : POLL,	value : 32'd91,	reg_addr : 32'd459560},
'{step_type : POLL,	value : 32'd112,	reg_addr : 32'd459561},
'{step_type : POLL,	value : 32'd133,	reg_addr : 32'd459562},
'{step_type : POLL,	value : 32'd157,	reg_addr : 32'd459563},
'{step_type : POLL,	value : 32'd178,	reg_addr : 32'd459564},
'{step_type : POLL,	value : 32'd199,	reg_addr : 32'd459565},
'{step_type : POLL,	value : 32'd223,	reg_addr : 32'd459566},
'{step_type : POLL,	value : 32'd244,	reg_addr : 32'd459567},
'{step_type : POLL,	value : 32'd265,	reg_addr : 32'd459568},
'{step_type : POLL,	value : 32'd275,	reg_addr : 32'd459569},
'{step_type : POLL,	value : 32'd277,	reg_addr : 32'd459570},
'{step_type : POLL,	value : 32'd281,	reg_addr : 32'd459571},
'{step_type : POLL,	value : 32'd283,	reg_addr : 32'd459572},
'{step_type : POLL,	value : 32'd287,	reg_addr : 32'd459573},
'{step_type : POLL,	value : 32'd289,	reg_addr : 32'd459574},
'{step_type : POLL,	value : 32'd290,	reg_addr : 32'd459575},
'{step_type : POLL,	value : 32'd291,	reg_addr : 32'd459577},
'{step_type : POLL,	value : 32'd293,	reg_addr : 32'd459578},
'{step_type : POLL,	value : 32'd295,	reg_addr : 32'd459579},
'{step_type : POLL,	value : 32'd296,	reg_addr : 32'd459580},
'{step_type : POLL,	value : 32'd321,	reg_addr : 32'd459581},
'{step_type : POLL,	value : 32'd331,	reg_addr : 32'd459582},
'{step_type : POLL,	value : 32'd355,	reg_addr : 32'd459583},
'{step_type : POLL,	value : 32'd371,	reg_addr : 32'd459600},
'{step_type : POLL,	value : 32'd395,	reg_addr : 32'd459601},
'{step_type : POLL,	value : 32'd404,	reg_addr : 32'd459602},
'{step_type : POLL,	value : 32'd422,	reg_addr : 32'd459603},
'{step_type : POLL,	value : 32'd24,	reg_addr : 32'd459659},
'{step_type : POLL,	value : 32'd45,	reg_addr : 32'd459660},
'{step_type : POLL,	value : 32'd66,	reg_addr : 32'd459661},
'{step_type : POLL,	value : 32'd90,	reg_addr : 32'd459662},
'{step_type : POLL,	value : 32'd111,	reg_addr : 32'd459663},
'{step_type : POLL,	value : 32'd132,	reg_addr : 32'd459664},
'{step_type : POLL,	value : 32'd156,	reg_addr : 32'd459665},
'{step_type : POLL,	value : 32'd177,	reg_addr : 32'd459666},
'{step_type : POLL,	value : 32'd198,	reg_addr : 32'd459667},
'{step_type : POLL,	value : 32'd222,	reg_addr : 32'd459668},
'{step_type : POLL,	value : 32'd243,	reg_addr : 32'd459669},
'{step_type : POLL,	value : 32'd264,	reg_addr : 32'd459670},
'{step_type : POLL,	value : 32'd274,	reg_addr : 32'd459671},
'{step_type : POLL,	value : 32'd276,	reg_addr : 32'd459672},
'{step_type : POLL,	value : 32'd280,	reg_addr : 32'd459673},
'{step_type : POLL,	value : 32'd282,	reg_addr : 32'd459674},
'{step_type : POLL,	value : 32'd286,	reg_addr : 32'd459675},
'{step_type : POLL,	value : 32'd288,	reg_addr : 32'd459676},
'{step_type : POLL,	value : 32'd289,	reg_addr : 32'd459677},
'{step_type : POLL,	value : 32'd290,	reg_addr : 32'd459678},
'{step_type : POLL,	value : 32'd292,	reg_addr : 32'd459680},
'{step_type : POLL,	value : 32'd294,	reg_addr : 32'd459681},
'{step_type : POLL,	value : 32'd295,	reg_addr : 32'd459682},
'{step_type : POLL,	value : 32'd320,	reg_addr : 32'd459683},
'{step_type : POLL,	value : 32'd330,	reg_addr : 32'd459684},
'{step_type : POLL,	value : 32'd354,	reg_addr : 32'd459685},
'{step_type : POLL,	value : 32'd370,	reg_addr : 32'd459686},
'{step_type : POLL,	value : 32'd394,	reg_addr : 32'd459703},
'{step_type : POLL,	value : 32'd403,	reg_addr : 32'd459704},
'{step_type : POLL,	value : 32'd421,	reg_addr : 32'd459705},
'{step_type : POLL,	value : 32'd438,	reg_addr : 32'd459706},
'{step_type : POLL,	value : 32'd1038,	reg_addr : 32'd459264},
'{step_type : POLL,	value : 32'd1103,	reg_addr : 32'd459266},
'{step_type : POLL,	value : 32'd192,	reg_addr : 32'd459268},
'{step_type : POLL,	value : 32'd582,	reg_addr : 32'd459269},
'{step_type : POLL,	value : 32'd257,	reg_addr : 32'd459270},
'{step_type : POLL,	value : 32'd647,	reg_addr : 32'd459271},
'{step_type : POLL,	value : 32'd322,	reg_addr : 32'd459272},
'{step_type : POLL,	value : 32'd712,	reg_addr : 32'd459273},
'{step_type : POLL,	value : 32'd18,	reg_addr : 32'd459274},
'{step_type : POLL,	value : 32'd844,	reg_addr : 32'd459275},
'{step_type : POLL,	value : 32'd21,	reg_addr : 32'd459276},
'{step_type : POLL,	value : 32'd22,	reg_addr : 32'd459278},
'{step_type : POLL,	value : 32'd23,	reg_addr : 32'd459280},
'{step_type : POLL,	value : 32'd44,	reg_addr : 32'd459282},
'{step_type : POLL,	value : 32'd24,	reg_addr : 32'd459283},
'{step_type : POLL,	value : 32'd45,	reg_addr : 32'd459284},
'{step_type : POLL,	value : 32'd25,	reg_addr : 32'd459285},
'{step_type : POLL,	value : 32'd46,	reg_addr : 32'd459286},
'{step_type : POLL,	value : 32'd26,	reg_addr : 32'd459287},
'{step_type : POLL,	value : 32'd47,	reg_addr : 32'd459288},
'{step_type : POLL,	value : 32'd27,	reg_addr : 32'd459289},
'{step_type : POLL,	value : 32'd19,	reg_addr : 32'd459290},
'{step_type : POLL,	value : 32'd618,	reg_addr : 32'd589852},
'{step_type : POLL,	value : 32'd618,	reg_addr : 32'd589853},
'{step_type : POLL,	value : 32'd618,	reg_addr : 32'd589854},
'{step_type : POLL,	value : 32'd618,	reg_addr : 32'd589855},
'{step_type : POLL,	value : 32'd674,	reg_addr : 32'd589856},
'{step_type : POLL,	value : 32'd618,	reg_addr : 32'd589857},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd589858},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd589859},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd589860},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd589861},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd589862},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd589863},
'{step_type : POLL,	value : 32'd671,	reg_addr : 32'd589867},
'{step_type : POLL,	value : 32'd2,	reg_addr : 32'd459077},
'{step_type : POLL,	value : 32'd51672,	reg_addr : 32'd266244},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266245},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266246},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266247},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266248},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266249},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266250},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266251},
'{step_type : POLL,	value : 32'd51544,	reg_addr : 32'd266252},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266253},
'{step_type : POLL,	value : 32'd53000,	reg_addr : 32'd266254},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266255},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266256},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266257},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266258},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266259},
'{step_type : POLL,	value : 32'd49368,	reg_addr : 32'd266260},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266261},
'{step_type : POLL,	value : 32'd55368,	reg_addr : 32'd266262},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266263},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266264},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266265},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266266},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266267},
'{step_type : POLL,	value : 32'd49496,	reg_addr : 32'd266268},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266269},
'{step_type : POLL,	value : 32'd56776,	reg_addr : 32'd266270},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266271},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266272},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266273},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266274},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266275},
'{step_type : POLL,	value : 32'd49624,	reg_addr : 32'd266276},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266277},
'{step_type : POLL,	value : 32'd49928,	reg_addr : 32'd266278},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266279},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266280},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266281},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266282},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266283},
'{step_type : POLL,	value : 32'd50520,	reg_addr : 32'd266284},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266285},
'{step_type : POLL,	value : 32'd60424,	reg_addr : 32'd266286},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266287},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266288},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266289},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266290},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266291},
'{step_type : POLL,	value : 32'd50648,	reg_addr : 32'd266292},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266293},
'{step_type : POLL,	value : 32'd55944,	reg_addr : 32'd266294},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266295},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266296},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266297},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266298},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266299},
'{step_type : POLL,	value : 32'd18648,	reg_addr : 32'd266300},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266301},
'{step_type : POLL,	value : 32'd23816,	reg_addr : 32'd266302},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266303},
'{step_type : POLL,	value : 32'd35032,	reg_addr : 32'd266304},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266305},
'{step_type : POLL,	value : 32'd40200,	reg_addr : 32'd266306},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266307},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266308},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266309},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266310},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266311},
'{step_type : POLL,	value : 32'd51800,	reg_addr : 32'd266312},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266313},
'{step_type : POLL,	value : 32'd49416,	reg_addr : 32'd266314},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266315},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266316},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266317},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266318},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266319},
'{step_type : POLL,	value : 32'd52056,	reg_addr : 32'd266320},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266321},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266322},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266323},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266324},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266325},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266326},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266327},
'{step_type : POLL,	value : 32'd54488,	reg_addr : 32'd266328},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266329},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266330},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266331},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266332},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266333},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266334},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266335},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266336},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266337},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266338},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266339},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266340},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266341},
'{step_type : POLL,	value : 32'd22408,	reg_addr : 32'd266342},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266343},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266344},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266345},
'{step_type : POLL,	value : 32'd38792,	reg_addr : 32'd266346},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266347},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266348},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266349},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266350},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266351},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266352},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266353},
'{step_type : POLL,	value : 32'd22472,	reg_addr : 32'd266354},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266355},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266356},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266357},
'{step_type : POLL,	value : 32'd38792,	reg_addr : 32'd266358},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266359},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266360},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266361},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266362},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266363},
'{step_type : POLL,	value : 32'd18264,	reg_addr : 32'd266364},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266365},
'{step_type : POLL,	value : 32'd18824,	reg_addr : 32'd266366},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266367},
'{step_type : POLL,	value : 32'd34648,	reg_addr : 32'd266368},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266369},
'{step_type : POLL,	value : 32'd35208,	reg_addr : 32'd266370},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266371},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266372},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266373},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266374},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266375},
'{step_type : POLL,	value : 32'd18392,	reg_addr : 32'd266376},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266377},
'{step_type : POLL,	value : 32'd26376,	reg_addr : 32'd266378},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266379},
'{step_type : POLL,	value : 32'd34776,	reg_addr : 32'd266380},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266381},
'{step_type : POLL,	value : 32'd42760,	reg_addr : 32'd266382},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266383},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266384},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266385},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266386},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266387},
'{step_type : POLL,	value : 32'd19544,	reg_addr : 32'd266388},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266389},
'{step_type : POLL,	value : 32'd18760,	reg_addr : 32'd266390},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266391},
'{step_type : POLL,	value : 32'd35928,	reg_addr : 32'd266392},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266393},
'{step_type : POLL,	value : 32'd35144,	reg_addr : 32'd266394},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266395},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266396},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266397},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266398},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266399},
'{step_type : POLL,	value : 32'd20312,	reg_addr : 32'd266400},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266401},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd266402},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266403},
'{step_type : POLL,	value : 32'd36696,	reg_addr : 32'd266404},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266405},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd266406},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266407},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266408},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266409},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266410},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266411},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266412},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266413},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266414},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266415},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266416},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266417},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266418},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266419},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266420},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266421},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266422},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266423},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266424},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266425},
'{step_type : POLL,	value : 32'd22408,	reg_addr : 32'd266426},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266427},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266428},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266429},
'{step_type : POLL,	value : 32'd38792,	reg_addr : 32'd266430},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266431},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266432},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266433},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266434},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266435},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266436},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266437},
'{step_type : POLL,	value : 32'd22408,	reg_addr : 32'd266438},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266439},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266440},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266441},
'{step_type : POLL,	value : 32'd38792,	reg_addr : 32'd266442},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266443},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266444},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266445},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266446},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266447},
'{step_type : POLL,	value : 32'd18264,	reg_addr : 32'd266448},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266449},
'{step_type : POLL,	value : 32'd18824,	reg_addr : 32'd266450},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266451},
'{step_type : POLL,	value : 32'd34648,	reg_addr : 32'd266452},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266453},
'{step_type : POLL,	value : 32'd35208,	reg_addr : 32'd266454},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266455},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266456},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266457},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266458},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266459},
'{step_type : POLL,	value : 32'd18392,	reg_addr : 32'd266460},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266461},
'{step_type : POLL,	value : 32'd26376,	reg_addr : 32'd266462},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266463},
'{step_type : POLL,	value : 32'd34776,	reg_addr : 32'd266464},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266465},
'{step_type : POLL,	value : 32'd42760,	reg_addr : 32'd266466},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266467},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266468},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266469},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266470},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266471},
'{step_type : POLL,	value : 32'd19544,	reg_addr : 32'd266472},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266473},
'{step_type : POLL,	value : 32'd18760,	reg_addr : 32'd266474},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266475},
'{step_type : POLL,	value : 32'd35928,	reg_addr : 32'd266476},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266477},
'{step_type : POLL,	value : 32'd35144,	reg_addr : 32'd266478},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266479},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266480},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266481},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266482},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266483},
'{step_type : POLL,	value : 32'd20312,	reg_addr : 32'd266484},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266485},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd266486},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266487},
'{step_type : POLL,	value : 32'd36696,	reg_addr : 32'd266488},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266489},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd266490},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266491},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266492},
'{step_type : POLL,	value : 32'd1258291200,	reg_addr : 32'd266493},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266494},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266495},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266496},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266497},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266498},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266499},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266500},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266501},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266502},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266503},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266504},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266505},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266506},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266507},
'{step_type : POLL,	value : 32'd51672,	reg_addr : 32'd266508},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266509},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266510},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266511},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266512},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266513},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266514},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266515},
'{step_type : POLL,	value : 32'd51544,	reg_addr : 32'd266516},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266517},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266518},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266519},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266520},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266521},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266522},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266523},
'{step_type : POLL,	value : 32'd49368,	reg_addr : 32'd266524},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266525},
'{step_type : POLL,	value : 32'd59400,	reg_addr : 32'd266526},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266527},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266528},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266529},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266530},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266531},
'{step_type : POLL,	value : 32'd49496,	reg_addr : 32'd266532},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266533},
'{step_type : POLL,	value : 32'd60040,	reg_addr : 32'd266534},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266535},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266536},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266537},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266538},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266539},
'{step_type : POLL,	value : 32'd49624,	reg_addr : 32'd266540},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266541},
'{step_type : POLL,	value : 32'd50952,	reg_addr : 32'd266542},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266543},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266544},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266545},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266546},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266547},
'{step_type : POLL,	value : 32'd50520,	reg_addr : 32'd266548},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266549},
'{step_type : POLL,	value : 32'd59912,	reg_addr : 32'd266550},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266551},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266552},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266553},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266554},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266555},
'{step_type : POLL,	value : 32'd50648,	reg_addr : 32'd266556},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266557},
'{step_type : POLL,	value : 32'd57864,	reg_addr : 32'd266558},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266559},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266560},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266561},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266562},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266563},
'{step_type : POLL,	value : 32'd18648,	reg_addr : 32'd266564},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266565},
'{step_type : POLL,	value : 32'd16968,	reg_addr : 32'd266566},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266567},
'{step_type : POLL,	value : 32'd35032,	reg_addr : 32'd266568},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266569},
'{step_type : POLL,	value : 32'd38472,	reg_addr : 32'd266570},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266571},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266572},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266573},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266574},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266575},
'{step_type : POLL,	value : 32'd51800,	reg_addr : 32'd266576},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266577},
'{step_type : POLL,	value : 32'd49416,	reg_addr : 32'd266578},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266579},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266580},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266581},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266582},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266583},
'{step_type : POLL,	value : 32'd52056,	reg_addr : 32'd266584},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266585},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266586},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266587},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266588},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266589},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266590},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266591},
'{step_type : POLL,	value : 32'd54488,	reg_addr : 32'd266592},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266593},
'{step_type : POLL,	value : 32'd61448,	reg_addr : 32'd266594},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266595},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266596},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266597},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266598},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266599},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266600},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266601},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266602},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266603},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266604},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266605},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266606},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266607},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266608},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266609},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266610},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266611},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266612},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266613},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266614},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266615},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266616},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266617},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266618},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266619},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266620},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266621},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266622},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266623},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266624},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266625},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266626},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266627},
'{step_type : POLL,	value : 32'd18264,	reg_addr : 32'd266628},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266629},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266630},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266631},
'{step_type : POLL,	value : 32'd34648,	reg_addr : 32'd266632},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266633},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266634},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266635},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266636},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266637},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266638},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266639},
'{step_type : POLL,	value : 32'd18392,	reg_addr : 32'd266640},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266641},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266642},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266643},
'{step_type : POLL,	value : 32'd34776,	reg_addr : 32'd266644},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266645},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266646},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266647},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266648},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266649},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266650},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266651},
'{step_type : POLL,	value : 32'd19544,	reg_addr : 32'd266652},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266653},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd266654},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266655},
'{step_type : POLL,	value : 32'd35928,	reg_addr : 32'd266656},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266657},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd266658},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266659},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266660},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266661},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266662},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266663},
'{step_type : POLL,	value : 32'd20312,	reg_addr : 32'd266664},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266665},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd266666},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266667},
'{step_type : POLL,	value : 32'd36696,	reg_addr : 32'd266668},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266669},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd266670},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266671},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266672},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266673},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266674},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266675},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266676},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266677},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266678},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266679},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266680},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266681},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266682},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266683},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266684},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266685},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266686},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266687},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266688},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266689},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266690},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266691},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266692},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266693},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266694},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266695},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266696},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266697},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266698},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266699},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266700},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266701},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266702},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266703},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266704},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266705},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266706},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266707},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266708},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266709},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266710},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266711},
'{step_type : POLL,	value : 32'd18264,	reg_addr : 32'd266712},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266713},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266714},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266715},
'{step_type : POLL,	value : 32'd34648,	reg_addr : 32'd266716},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266717},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266718},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266719},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266720},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266721},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266722},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266723},
'{step_type : POLL,	value : 32'd18392,	reg_addr : 32'd266724},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266725},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266726},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266727},
'{step_type : POLL,	value : 32'd34776,	reg_addr : 32'd266728},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266729},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266730},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266731},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266732},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266733},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266734},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266735},
'{step_type : POLL,	value : 32'd19544,	reg_addr : 32'd266736},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266737},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd266738},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266739},
'{step_type : POLL,	value : 32'd35928,	reg_addr : 32'd266740},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266741},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd266742},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266743},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266744},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266745},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266746},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266747},
'{step_type : POLL,	value : 32'd20312,	reg_addr : 32'd266748},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266749},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd266750},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266751},
'{step_type : POLL,	value : 32'd36696,	reg_addr : 32'd266752},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266753},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd266754},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266755},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266756},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266757},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266758},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266759},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266760},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266761},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266762},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266763},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266764},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266765},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266766},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266767},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266768},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266769},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266770},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266771},
'{step_type : POLL,	value : 32'd51672,	reg_addr : 32'd266772},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266773},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266774},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266775},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266776},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266777},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266778},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266779},
'{step_type : POLL,	value : 32'd51544,	reg_addr : 32'd266780},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266781},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266782},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266783},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266784},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266785},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266786},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266787},
'{step_type : POLL,	value : 32'd49368,	reg_addr : 32'd266788},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266789},
'{step_type : POLL,	value : 32'd59400,	reg_addr : 32'd266790},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266791},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266792},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266793},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266794},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266795},
'{step_type : POLL,	value : 32'd49496,	reg_addr : 32'd266796},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266797},
'{step_type : POLL,	value : 32'd60040,	reg_addr : 32'd266798},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266799},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266800},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266801},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266802},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266803},
'{step_type : POLL,	value : 32'd49624,	reg_addr : 32'd266804},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266805},
'{step_type : POLL,	value : 32'd50952,	reg_addr : 32'd266806},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266807},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266808},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266809},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266810},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266811},
'{step_type : POLL,	value : 32'd50520,	reg_addr : 32'd266812},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266813},
'{step_type : POLL,	value : 32'd59912,	reg_addr : 32'd266814},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266815},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266816},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266817},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266818},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266819},
'{step_type : POLL,	value : 32'd50648,	reg_addr : 32'd266820},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266821},
'{step_type : POLL,	value : 32'd57864,	reg_addr : 32'd266822},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266823},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266824},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266825},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266826},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266827},
'{step_type : POLL,	value : 32'd18648,	reg_addr : 32'd266828},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266829},
'{step_type : POLL,	value : 32'd16968,	reg_addr : 32'd266830},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266831},
'{step_type : POLL,	value : 32'd35032,	reg_addr : 32'd266832},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266833},
'{step_type : POLL,	value : 32'd38472,	reg_addr : 32'd266834},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266835},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266836},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266837},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266838},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266839},
'{step_type : POLL,	value : 32'd51800,	reg_addr : 32'd266840},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266841},
'{step_type : POLL,	value : 32'd49416,	reg_addr : 32'd266842},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266843},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266844},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266845},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266846},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266847},
'{step_type : POLL,	value : 32'd52056,	reg_addr : 32'd266848},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266849},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd266850},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266851},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266852},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266853},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266854},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266855},
'{step_type : POLL,	value : 32'd54488,	reg_addr : 32'd266856},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266857},
'{step_type : POLL,	value : 32'd61448,	reg_addr : 32'd266858},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266859},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266860},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266861},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266862},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266863},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266864},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266865},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266866},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266867},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266868},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266869},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266870},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266871},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266872},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266873},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266874},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266875},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266876},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266877},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266878},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266879},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266880},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266881},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266882},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266883},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266884},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266885},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266886},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266887},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266888},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266889},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266890},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266891},
'{step_type : POLL,	value : 32'd18264,	reg_addr : 32'd266892},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266893},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266894},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266895},
'{step_type : POLL,	value : 32'd34648,	reg_addr : 32'd266896},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266897},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266898},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266899},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266900},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266901},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266902},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266903},
'{step_type : POLL,	value : 32'd18392,	reg_addr : 32'd266904},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266905},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266906},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266907},
'{step_type : POLL,	value : 32'd34776,	reg_addr : 32'd266908},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266909},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266910},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266911},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266912},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266913},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266914},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266915},
'{step_type : POLL,	value : 32'd19544,	reg_addr : 32'd266916},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266917},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd266918},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266919},
'{step_type : POLL,	value : 32'd35928,	reg_addr : 32'd266920},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266921},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd266922},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266923},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266924},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266925},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266926},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266927},
'{step_type : POLL,	value : 32'd20312,	reg_addr : 32'd266928},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266929},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd266930},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266931},
'{step_type : POLL,	value : 32'd36696,	reg_addr : 32'd266932},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266933},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd266934},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266935},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266936},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266937},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266938},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266939},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266940},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266941},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266942},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266943},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266944},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266945},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266946},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266947},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266948},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266949},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266950},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266951},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266952},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266953},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266954},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266955},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266956},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266957},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266958},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266959},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266960},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266961},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266962},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266963},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd266964},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266965},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266966},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266967},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd266968},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266969},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266970},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266971},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266972},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266973},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266974},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266975},
'{step_type : POLL,	value : 32'd18264,	reg_addr : 32'd266976},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266977},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266978},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266979},
'{step_type : POLL,	value : 32'd34648,	reg_addr : 32'd266980},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266981},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266982},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266983},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266984},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266985},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266986},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266987},
'{step_type : POLL,	value : 32'd18392,	reg_addr : 32'd266988},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266989},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd266990},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266991},
'{step_type : POLL,	value : 32'd34776,	reg_addr : 32'd266992},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266993},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd266994},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266995},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266996},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd266997},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266998},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd266999},
'{step_type : POLL,	value : 32'd19544,	reg_addr : 32'd267000},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267001},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd267002},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267003},
'{step_type : POLL,	value : 32'd35928,	reg_addr : 32'd267004},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267005},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd267006},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267007},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267008},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267009},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267010},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267011},
'{step_type : POLL,	value : 32'd20312,	reg_addr : 32'd267012},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267013},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd267014},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267015},
'{step_type : POLL,	value : 32'd36696,	reg_addr : 32'd267016},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267017},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd267018},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267019},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267020},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267021},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267022},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267023},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267024},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267025},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267026},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267027},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267028},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267029},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267030},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267031},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267032},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267033},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267034},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267035},
'{step_type : POLL,	value : 32'd51672,	reg_addr : 32'd267036},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267037},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267038},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267039},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267040},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267041},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267042},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267043},
'{step_type : POLL,	value : 32'd51544,	reg_addr : 32'd267044},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267045},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267046},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267047},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267048},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267049},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267050},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267051},
'{step_type : POLL,	value : 32'd49368,	reg_addr : 32'd267052},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267053},
'{step_type : POLL,	value : 32'd59400,	reg_addr : 32'd267054},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267055},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267056},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267057},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267058},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267059},
'{step_type : POLL,	value : 32'd49496,	reg_addr : 32'd267060},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267061},
'{step_type : POLL,	value : 32'd60040,	reg_addr : 32'd267062},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267063},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267064},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267065},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267066},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267067},
'{step_type : POLL,	value : 32'd49624,	reg_addr : 32'd267068},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267069},
'{step_type : POLL,	value : 32'd50952,	reg_addr : 32'd267070},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267071},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267072},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267073},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267074},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267075},
'{step_type : POLL,	value : 32'd50520,	reg_addr : 32'd267076},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267077},
'{step_type : POLL,	value : 32'd59912,	reg_addr : 32'd267078},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267079},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267080},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267081},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267082},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267083},
'{step_type : POLL,	value : 32'd50648,	reg_addr : 32'd267084},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267085},
'{step_type : POLL,	value : 32'd57864,	reg_addr : 32'd267086},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267087},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267088},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267089},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267090},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267091},
'{step_type : POLL,	value : 32'd18648,	reg_addr : 32'd267092},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267093},
'{step_type : POLL,	value : 32'd16968,	reg_addr : 32'd267094},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267095},
'{step_type : POLL,	value : 32'd35032,	reg_addr : 32'd267096},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267097},
'{step_type : POLL,	value : 32'd38472,	reg_addr : 32'd267098},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267099},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267100},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267101},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267102},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267103},
'{step_type : POLL,	value : 32'd51800,	reg_addr : 32'd267104},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267105},
'{step_type : POLL,	value : 32'd49416,	reg_addr : 32'd267106},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267107},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267108},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267109},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267110},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267111},
'{step_type : POLL,	value : 32'd52056,	reg_addr : 32'd267112},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267113},
'{step_type : POLL,	value : 32'd49160,	reg_addr : 32'd267114},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267115},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267116},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267117},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267118},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267119},
'{step_type : POLL,	value : 32'd54488,	reg_addr : 32'd267120},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267121},
'{step_type : POLL,	value : 32'd61448,	reg_addr : 32'd267122},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267123},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267124},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267125},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267126},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267127},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267128},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267129},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267130},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267131},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd267132},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267133},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd267134},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267135},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd267136},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267137},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd267138},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267139},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267140},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267141},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267142},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267143},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd267144},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267145},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd267146},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267147},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd267148},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267149},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd267150},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267151},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267152},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267153},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267154},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267155},
'{step_type : POLL,	value : 32'd18264,	reg_addr : 32'd267156},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267157},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd267158},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267159},
'{step_type : POLL,	value : 32'd34648,	reg_addr : 32'd267160},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267161},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd267162},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267163},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267164},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267165},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267166},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267167},
'{step_type : POLL,	value : 32'd18392,	reg_addr : 32'd267168},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267169},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd267170},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267171},
'{step_type : POLL,	value : 32'd34776,	reg_addr : 32'd267172},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267173},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd267174},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267175},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267176},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267177},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267178},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267179},
'{step_type : POLL,	value : 32'd19544,	reg_addr : 32'd267180},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267181},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd267182},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267183},
'{step_type : POLL,	value : 32'd35928,	reg_addr : 32'd267184},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267185},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd267186},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267187},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267188},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267189},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267190},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267191},
'{step_type : POLL,	value : 32'd20312,	reg_addr : 32'd267192},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267193},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd267194},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267195},
'{step_type : POLL,	value : 32'd36696,	reg_addr : 32'd267196},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267197},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd267198},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267199},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267200},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267201},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267202},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267203},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267204},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267205},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267206},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267207},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267208},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267209},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267210},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267211},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267212},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267213},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267214},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267215},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd267216},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267217},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd267218},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267219},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd267220},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267221},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd267222},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267223},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267224},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267225},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267226},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267227},
'{step_type : POLL,	value : 32'd18008,	reg_addr : 32'd267228},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267229},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd267230},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267231},
'{step_type : POLL,	value : 32'd34392,	reg_addr : 32'd267232},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267233},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd267234},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267235},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267236},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267237},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267238},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267239},
'{step_type : POLL,	value : 32'd18264,	reg_addr : 32'd267240},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267241},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd267242},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267243},
'{step_type : POLL,	value : 32'd34648,	reg_addr : 32'd267244},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267245},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd267246},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267247},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267248},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267249},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267250},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267251},
'{step_type : POLL,	value : 32'd18392,	reg_addr : 32'd267252},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267253},
'{step_type : POLL,	value : 32'd26632,	reg_addr : 32'd267254},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267255},
'{step_type : POLL,	value : 32'd34776,	reg_addr : 32'd267256},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267257},
'{step_type : POLL,	value : 32'd43016,	reg_addr : 32'd267258},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267259},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267260},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267261},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267262},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267263},
'{step_type : POLL,	value : 32'd19544,	reg_addr : 32'd267264},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267265},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd267266},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267267},
'{step_type : POLL,	value : 32'd35928,	reg_addr : 32'd267268},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267269},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd267270},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267271},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267272},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267273},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267274},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267275},
'{step_type : POLL,	value : 32'd20312,	reg_addr : 32'd267276},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267277},
'{step_type : POLL,	value : 32'd16392,	reg_addr : 32'd267278},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267279},
'{step_type : POLL,	value : 32'd36696,	reg_addr : 32'd267280},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267281},
'{step_type : POLL,	value : 32'd32776,	reg_addr : 32'd267282},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267283},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267284},
'{step_type : POLL,	value : 32'd721420288,	reg_addr : 32'd267285},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267286},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267287},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267288},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267289},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267290},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267291},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267292},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267293},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267294},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267295},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267296},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267297},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267298},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd267299},
'{step_type : POLL,	value : 32'd22561,	reg_addr : 32'd786433},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591628},
'{step_type : POLL,	value : 32'd254,	reg_addr : 32'd591629},
'{step_type : POLL,	value : 32'd65535,	reg_addr : 32'd591630},
'{step_type : POLL,	value : 32'd61504,	reg_addr : 32'd591631},
'{step_type : POLL,	value : 32'd61504,	reg_addr : 32'd591632},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591633},
'{step_type : POLL,	value : 32'd65535,	reg_addr : 32'd591634},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591635},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591636},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591637},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591638},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591639},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591640},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591641},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591642},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd591643},
'{step_type : POLL,	value : 32'd2925,	reg_addr : 32'd458992},
'{step_type : POLL,	value : 32'd195,	reg_addr : 32'd458878},
'{step_type : POLL,	value : 32'd32767,	reg_addr : 32'd459247},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd196774},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd200870},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459176},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459048},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459057},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459058},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459059},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459060},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459074},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd459076},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd721683},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd852017},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd786483},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd786484},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd786486},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65726},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65982},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd66238},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd66494},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd66750},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd67006},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd67262},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd67518},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd67774},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65712},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65664},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd65665},
'{step_type : POLL,	value : 32'd2,	reg_addr : 32'd65666},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd65667},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd65668},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd65669},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd65670},
'{step_type : POLL,	value : 32'd7,	reg_addr : 32'd65671},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd65672},
'{step_type : POLL,	value : 32'd156,	reg_addr : 32'd65753},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd65585},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69822},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd70078},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd70334},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd70590},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd70846},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd71102},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd71358},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd71614},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd71870},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69808},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69760},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd69761},
'{step_type : POLL,	value : 32'd2,	reg_addr : 32'd69762},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd69763},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd69764},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd69765},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd69766},
'{step_type : POLL,	value : 32'd7,	reg_addr : 32'd69767},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd69768},
'{step_type : POLL,	value : 32'd156,	reg_addr : 32'd69849},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd69681},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73918},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd74174},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd74430},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd74686},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd74942},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd75198},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd75454},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd75710},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd75966},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73904},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73856},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd73857},
'{step_type : POLL,	value : 32'd2,	reg_addr : 32'd73858},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd73859},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd73860},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd73861},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd73862},
'{step_type : POLL,	value : 32'd7,	reg_addr : 32'd73863},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd73864},
'{step_type : POLL,	value : 32'd156,	reg_addr : 32'd73945},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd73777},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78014},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78270},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78526},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78782},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd79038},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd79294},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd79550},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd79806},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd80062},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78000},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd77952},
'{step_type : POLL,	value : 32'd1,	reg_addr : 32'd77953},
'{step_type : POLL,	value : 32'd2,	reg_addr : 32'd77954},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd77955},
'{step_type : POLL,	value : 32'd4,	reg_addr : 32'd77956},
'{step_type : POLL,	value : 32'd5,	reg_addr : 32'd77957},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd77958},
'{step_type : POLL,	value : 32'd7,	reg_addr : 32'd77959},
'{step_type : POLL,	value : 32'd8,	reg_addr : 32'd77960},
'{step_type : POLL,	value : 32'd156,	reg_addr : 32'd78041},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd77873},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917516},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921612},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917542},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921638},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917543},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921639},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917544},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921640},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917545},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921641},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921642},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925708},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929804},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925734},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929830},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925735},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929831},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925736},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929832},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925737},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929833},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929834},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933900},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd937996},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933926},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938022},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933927},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938023},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933928},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938024},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd933929},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938025},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938026},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942092},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946188},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942118},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946214},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942119},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946215},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942120},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946216},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942121},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946217},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946218},
'{step_type : POLL,	value : 32'd102,	reg_addr : 32'd131185},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd196825},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd196824},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd197080},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd197336},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd197592},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd197848},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd198104},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd198360},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd198616},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd198872},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd199128},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd200921},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd200920},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd201176},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd201432},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd201688},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd201944},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd202200},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd202456},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd202712},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd202968},
'{step_type : POLL,	value : 32'd64,	reg_addr : 32'd203224},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1632},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1633},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1376},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1377},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd5728},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd5729},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd5472},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd5473},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd9824},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd9825},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd9568},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd9569},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd13920},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd13921},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd13664},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd13665},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd18016},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd18017},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd17760},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd17761},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd30304},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd30305},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd30048},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd30049},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd34400},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd34401},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd34144},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd34145},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd38496},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd38497},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd38240},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd38241},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd42592},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd42593},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd42336},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd42337},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd46688},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd46689},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd46432},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd46433},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd65536},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd66221},
'{step_type : POLL,	value : 32'd76,	reg_addr : 32'd66223},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd66208},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd66209},
'{step_type : POLL,	value : 32'd10,	reg_addr : 32'd66210},
'{step_type : POLL,	value : 32'd62,	reg_addr : 32'd66211},
'{step_type : POLL,	value : 32'd114,	reg_addr : 32'd66212},
'{step_type : POLL,	value : 32'd793,	reg_addr : 32'd65568},
'{step_type : POLL,	value : 32'd793,	reg_addr : 32'd65569},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd65576},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd65577},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd65578},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd65579},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd65656},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd65657},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd65658},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd65659},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd65552},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd65553},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd65554},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd65555},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd65736},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65640},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65641},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65642},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65643},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65644},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65645},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65646},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65647},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65632},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65633},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65635},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65636},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd65912},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd65913},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd65914},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd65915},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd65808},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd65809},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd65810},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd65811},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd65992},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65896},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65897},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65898},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65899},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65900},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65901},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65902},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65903},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65888},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65889},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65891},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65892},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd66168},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd66169},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd66170},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd66171},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66064},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66065},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66066},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66067},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd66248},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66152},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66153},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66154},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66155},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66156},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66157},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66158},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66159},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66144},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66145},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66147},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66148},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd66424},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd66425},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd66426},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd66427},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66320},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66321},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66322},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66323},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd66504},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66408},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66409},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66410},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66411},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66412},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66413},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66414},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66415},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66400},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66401},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66403},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66404},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd66680},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd66681},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd66682},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd66683},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66576},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66577},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66578},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66579},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd66760},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66664},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66665},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66666},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66667},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66668},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66669},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66670},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66671},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66656},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66657},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66659},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66660},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd66936},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd66937},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd66938},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd66939},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66832},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66833},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66834},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd66835},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd67016},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66920},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66921},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66922},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66923},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66924},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66925},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66926},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66927},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66912},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66913},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66915},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd66916},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd67192},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd67193},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd67194},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd67195},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67088},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67089},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67090},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67091},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd67272},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67176},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67177},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67178},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67179},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67180},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67181},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67182},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67183},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67168},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67169},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67171},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67172},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd67448},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd67449},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd67450},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd67451},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67344},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67345},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67346},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67347},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd67528},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67432},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67433},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67434},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67435},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67436},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67437},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67438},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67439},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67424},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67425},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67427},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67428},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd67704},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd67705},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd67706},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd67707},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67600},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67601},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67602},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd67603},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd67784},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67688},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67689},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67690},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67691},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67692},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67693},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67694},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67695},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67680},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67681},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67683},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd67684},
'{step_type : POLL,	value : 32'd204,	reg_addr : 32'd65548},
'{step_type : POLL,	value : 32'd204,	reg_addr : 32'd65549},
'{step_type : POLL,	value : 32'd408,	reg_addr : 32'd65556},
'{step_type : POLL,	value : 32'd408,	reg_addr : 32'd65557},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65561},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65563},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65570},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd65571},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd65887},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd69632},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd70317},
'{step_type : POLL,	value : 32'd76,	reg_addr : 32'd70319},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd70304},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd70305},
'{step_type : POLL,	value : 32'd10,	reg_addr : 32'd70306},
'{step_type : POLL,	value : 32'd62,	reg_addr : 32'd70307},
'{step_type : POLL,	value : 32'd114,	reg_addr : 32'd70308},
'{step_type : POLL,	value : 32'd793,	reg_addr : 32'd69664},
'{step_type : POLL,	value : 32'd793,	reg_addr : 32'd69665},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd69672},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd69673},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd69674},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd69675},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd69752},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd69753},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd69754},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd69755},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd69648},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd69649},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd69650},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd69651},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd69832},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69736},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69737},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69738},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69739},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69740},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69741},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69742},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69743},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69728},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69729},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69731},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69732},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd70008},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd70009},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd70010},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd70011},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd69904},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd69905},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd69906},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd69907},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd70088},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69992},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69993},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69994},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69995},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69996},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69997},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69998},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69999},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69984},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69985},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69987},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69988},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd70264},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd70265},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd70266},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd70267},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70160},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70161},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70162},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70163},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd70344},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70248},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70249},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70250},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70251},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70252},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70253},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70254},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70255},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70240},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70241},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70243},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70244},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd70520},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd70521},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd70522},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd70523},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70416},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70417},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70418},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70419},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd70600},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70504},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70505},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70506},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70507},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70508},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70509},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70510},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70511},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70496},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70497},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70499},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70500},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd70776},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd70777},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd70778},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd70779},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70672},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70673},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70674},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70675},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd70856},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70760},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70761},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70762},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70763},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70764},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70765},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70766},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70767},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70752},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70753},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70755},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd70756},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd71032},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd71033},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd71034},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd71035},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70928},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70929},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70930},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd70931},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd71112},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71016},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71017},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71018},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71019},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71020},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71021},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71022},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71023},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71008},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71009},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71011},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71012},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd71288},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd71289},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd71290},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd71291},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71184},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71185},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71186},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71187},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd71368},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71272},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71273},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71274},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71275},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71276},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71277},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71278},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71279},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71264},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71265},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71267},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71268},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd71544},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd71545},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd71546},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd71547},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71440},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71441},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71442},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71443},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd71624},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71528},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71529},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71530},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71531},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71532},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71533},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71534},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71535},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71520},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71521},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71523},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71524},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd71800},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd71801},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd71802},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd71803},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71696},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71697},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71698},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd71699},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd71880},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71784},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71785},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71786},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71787},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71788},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71789},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71790},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71791},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71776},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71777},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71779},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd71780},
'{step_type : POLL,	value : 32'd204,	reg_addr : 32'd69644},
'{step_type : POLL,	value : 32'd204,	reg_addr : 32'd69645},
'{step_type : POLL,	value : 32'd408,	reg_addr : 32'd69652},
'{step_type : POLL,	value : 32'd408,	reg_addr : 32'd69653},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69657},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69659},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69666},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd69667},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd69983},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd73728},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd74413},
'{step_type : POLL,	value : 32'd76,	reg_addr : 32'd74415},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd74400},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd74401},
'{step_type : POLL,	value : 32'd10,	reg_addr : 32'd74402},
'{step_type : POLL,	value : 32'd62,	reg_addr : 32'd74403},
'{step_type : POLL,	value : 32'd114,	reg_addr : 32'd74404},
'{step_type : POLL,	value : 32'd793,	reg_addr : 32'd73760},
'{step_type : POLL,	value : 32'd793,	reg_addr : 32'd73761},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd73768},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd73769},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd73770},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd73771},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd73848},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd73849},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd73850},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd73851},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd73744},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd73745},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd73746},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd73747},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd73928},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73832},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73833},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73834},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73835},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73836},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73837},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73838},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73839},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73824},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73825},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73827},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73828},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd74104},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd74105},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd74106},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd74107},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74000},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74001},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74002},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74003},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd74184},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74088},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74089},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74090},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74091},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74092},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74093},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74094},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74095},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74080},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74081},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74083},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74084},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd74360},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd74361},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd74362},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd74363},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74256},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74257},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74258},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74259},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd74440},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74344},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74345},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74346},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74347},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74348},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74349},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74350},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74351},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74336},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74337},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74339},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74340},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd74616},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd74617},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd74618},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd74619},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74512},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74513},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74514},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74515},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd74696},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74600},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74601},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74602},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74603},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74604},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74605},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74606},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74607},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74592},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74593},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74595},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74596},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd74872},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd74873},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd74874},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd74875},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74768},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74769},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74770},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd74771},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd74952},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74856},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74857},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74858},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74859},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74860},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74861},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74862},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74863},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74848},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74849},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74851},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd74852},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd75128},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd75129},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd75130},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd75131},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75024},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75025},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75026},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75027},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd75208},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75112},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75113},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75114},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75115},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75116},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75117},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75118},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75119},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75104},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75105},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75107},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75108},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd75384},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd75385},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd75386},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd75387},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75280},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75281},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75282},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75283},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd75464},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75368},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75369},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75370},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75371},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75372},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75373},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75374},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75375},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75360},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75361},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75363},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75364},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd75640},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd75641},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd75642},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd75643},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75536},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75537},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75538},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75539},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd75720},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75624},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75625},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75626},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75627},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75628},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75629},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75630},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75631},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75616},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75617},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75619},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75620},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd75896},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd75897},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd75898},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd75899},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75792},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75793},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75794},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd75795},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd75976},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75880},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75881},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75882},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75883},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75884},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75885},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75886},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75887},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75872},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75873},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75875},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd75876},
'{step_type : POLL,	value : 32'd204,	reg_addr : 32'd73740},
'{step_type : POLL,	value : 32'd204,	reg_addr : 32'd73741},
'{step_type : POLL,	value : 32'd408,	reg_addr : 32'd73748},
'{step_type : POLL,	value : 32'd408,	reg_addr : 32'd73749},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73753},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73755},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73762},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd73763},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd74079},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd77824},
'{step_type : POLL,	value : 32'd3,	reg_addr : 32'd78509},
'{step_type : POLL,	value : 32'd76,	reg_addr : 32'd78511},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78496},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd78497},
'{step_type : POLL,	value : 32'd10,	reg_addr : 32'd78498},
'{step_type : POLL,	value : 32'd62,	reg_addr : 32'd78499},
'{step_type : POLL,	value : 32'd114,	reg_addr : 32'd78500},
'{step_type : POLL,	value : 32'd793,	reg_addr : 32'd77856},
'{step_type : POLL,	value : 32'd793,	reg_addr : 32'd77857},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd77864},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd77865},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd77866},
'{step_type : POLL,	value : 32'd512,	reg_addr : 32'd77867},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd77944},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd77945},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd77946},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd77947},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd77840},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd77841},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd77842},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd77843},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd78024},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77928},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77929},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77930},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77931},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77932},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77933},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77934},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77935},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77920},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77921},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77923},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77924},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd78200},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd78201},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd78202},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd78203},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78096},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78097},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78098},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78099},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd78280},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78184},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78185},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78186},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78187},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78188},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78189},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78190},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78191},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78176},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78177},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78179},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78180},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd78456},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd78457},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd78458},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd78459},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78352},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78353},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78354},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78355},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd78536},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78440},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78441},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78442},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78443},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78444},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78445},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78446},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78447},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78432},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78433},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78435},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78436},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd78712},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd78713},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd78714},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd78715},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78608},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78609},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78610},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78611},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd78792},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78696},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78697},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78698},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78699},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78700},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78701},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78702},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78703},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78688},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78689},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78691},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78692},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd78968},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd78969},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd78970},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd78971},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78864},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78865},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78866},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd78867},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd79048},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78952},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78953},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78954},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78955},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78956},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78957},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78958},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78959},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78944},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78945},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78947},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd78948},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd79224},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd79225},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd79226},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd79227},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79120},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79121},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79122},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79123},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd79304},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79208},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79209},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79210},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79211},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79212},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79213},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79214},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79215},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79200},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79201},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79203},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79204},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd79480},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd79481},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd79482},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd79483},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79376},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79377},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79378},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79379},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd79560},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79464},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79465},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79466},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79467},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79468},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79469},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79470},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79471},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79456},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79457},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79459},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79460},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd79736},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd79737},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd79738},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd79739},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79632},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79633},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79634},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79635},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd79816},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79720},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79721},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79722},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79723},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79724},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79725},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79726},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79727},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79712},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79713},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79715},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79716},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd79992},
'{step_type : POLL,	value : 32'd953,	reg_addr : 32'd79993},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd79994},
'{step_type : POLL,	value : 32'd237,	reg_addr : 32'd79995},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79888},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79889},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79890},
'{step_type : POLL,	value : 32'd299,	reg_addr : 32'd79891},
'{step_type : POLL,	value : 32'd255,	reg_addr : 32'd80072},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79976},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79977},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79978},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79979},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79980},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79981},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79982},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79983},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79968},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79969},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79971},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd79972},
'{step_type : POLL,	value : 32'd204,	reg_addr : 32'd77836},
'{step_type : POLL,	value : 32'd204,	reg_addr : 32'd77837},
'{step_type : POLL,	value : 32'd408,	reg_addr : 32'd77844},
'{step_type : POLL,	value : 32'd408,	reg_addr : 32'd77845},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77849},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77851},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77858},
'{step_type : POLL,	value : 32'd31,	reg_addr : 32'd77859},
'{step_type : POLL,	value : 32'd98,	reg_addr : 32'd78175},
'{step_type : POLL,	value : 32'd16,	reg_addr : 32'd393225},
'{step_type : POLL,	value : 32'd6,	reg_addr : 32'd458765},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917616},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921712},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917617},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921713},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917618},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921714},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917619},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921715},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921716},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917621},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921717},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917622},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921718},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917623},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921719},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917624},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921720},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921721},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917744},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921840},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917745},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921841},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917746},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921842},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917747},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921843},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921844},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917749},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921845},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd918016},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd922112},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd918017},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd922113},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd918018},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd922114},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd918019},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd922115},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd922116},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd918021},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd922117},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917664},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921760},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917680},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921776},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917696},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921792},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917712},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921808},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921824},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917665},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921761},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917681},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921777},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917697},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921793},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917713},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921809},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921825},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917668},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921764},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917684},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921780},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917700},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921796},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917716},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921812},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921828},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917669},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921765},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917685},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921781},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917701},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921797},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd917717},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921813},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd921829},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd918864},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd922960},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd918865},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd918880},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd922976},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd918881},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd922977},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd918896},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd922992},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd918897},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd922993},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd918912},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd923008},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd918913},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd923009},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925808},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929904},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925809},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929905},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925810},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929906},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925811},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929907},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929908},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925813},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929909},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925814},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929910},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925815},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929911},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925816},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929912},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929913},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925936},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930032},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925937},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930033},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925938},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930034},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925939},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930035},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930036},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925941},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930037},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd926208},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930304},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd926209},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930305},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd926210},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930306},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd926211},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930307},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930308},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd926213},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930309},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925856},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929952},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925872},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929968},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925888},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929984},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925904},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930000},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930016},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925857},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929953},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925873},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929969},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925889},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929985},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925905},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930001},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930017},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925860},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929956},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925876},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929972},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925892},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929988},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925908},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930004},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930020},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925861},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929957},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925877},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929973},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925893},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd929989},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd925909},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930005},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd930021},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd927056},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd931152},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd927057},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd927072},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd931168},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd927073},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd931169},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd927088},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd931184},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd927089},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd931185},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd927104},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd931200},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd927105},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd931201},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934000},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938096},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934001},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938097},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934002},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938098},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934003},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938099},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938100},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934005},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938101},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934006},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938102},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934007},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938103},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934008},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938104},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938105},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934128},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938224},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934129},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938225},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934130},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938226},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934131},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938227},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938228},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934133},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938229},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934400},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938496},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934401},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938497},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934402},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938498},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934403},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938499},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938500},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934405},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938501},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934048},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938144},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934064},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938160},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934080},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938176},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934096},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938192},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938208},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934049},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938145},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934065},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938161},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934081},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938177},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934097},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938193},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938209},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934052},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938148},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934068},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938164},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934084},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938180},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934100},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938196},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938212},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934053},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938149},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934069},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938165},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934085},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938181},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd934101},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938197},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd938213},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd935248},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd939344},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd935249},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd935264},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd939360},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd935265},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd939361},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd935280},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd939376},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd935281},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd939377},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd935296},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd939392},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd935297},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd939393},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942192},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946288},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942193},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946289},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942194},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946290},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942195},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946291},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946292},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942197},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946293},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942198},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946294},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942199},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946295},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942200},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946296},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946297},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942320},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946416},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942321},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946417},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942322},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946418},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942323},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946419},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946420},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942325},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946421},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942592},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946688},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942593},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946689},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942594},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946690},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942595},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946691},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946692},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942597},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946693},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942240},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946336},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942256},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946352},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942272},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946368},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942288},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946384},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946400},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942241},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946337},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942257},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946353},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942273},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946369},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942289},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946385},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946401},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942244},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946340},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942260},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946356},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942276},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946372},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942292},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946388},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946404},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942245},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946341},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942261},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946357},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942277},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946373},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd942293},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946389},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd946405},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd943440},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd947536},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd943441},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd943456},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd947552},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd943457},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd947553},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd943472},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd947568},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd943473},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd947569},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd943488},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd947584},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd943489},
'{step_type : POLL,	value : 32'd870,	reg_addr : 32'd947585},
'{step_type : POLL,	value : 32'd38657,	reg_addr : 32'd591879},
'{step_type : POLL,	value : 32'd46721,	reg_addr : 32'd591880},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd458871},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd131079},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd720897},
'{step_type : REG_WRITE,	value : 32'd4,	reg_addr : 32'd786560},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd851968},
'{step_type : REG_WRITE,	value : 32'd0,	reg_addr : 32'd851968},
'{step_type : REG_WRITE,	value : 32'd6,	reg_addr : 32'd131077},
'{step_type : REG_WRITE,	value : 32'd9,	reg_addr : 32'd458855},
'{step_type : REG_WRITE,	value : 32'd9,	reg_addr : 32'd458983},
'{step_type : POLL,	value : 32'd91,	reg_addr : 32'd458816},
'{step_type : REG_WRITE,	value : 32'd94,	reg_addr : 32'd458816},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1507392},
'{step_type : REG_WRITE,	value : 32'd14,	reg_addr : 32'd1507392},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd2555968},
'{step_type : REG_WRITE,	value : 32'd14,	reg_addr : 32'd2555968},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd3604544},
'{step_type : REG_WRITE,	value : 32'd14,	reg_addr : 32'd3604544},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd458854},
'{step_type : REG_WRITE,	value : 32'd2848,	reg_addr : 32'd458854},
'{step_type : POLL,	value : 32'd32,	reg_addr : 32'd458982},
'{step_type : REG_WRITE,	value : 32'd2848,	reg_addr : 32'd458982},
'{step_type : POLL,	value : 32'd546,	reg_addr : 32'd458859},
'{step_type : REG_WRITE,	value : 32'd2850,	reg_addr : 32'd458859},
'{step_type : POLL,	value : 32'd546,	reg_addr : 32'd458987},
'{step_type : REG_WRITE,	value : 32'd2850,	reg_addr : 32'd458987},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1507430},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd1507430},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1507558},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd1507558},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1507435},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd1507435},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd1507563},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd1507563},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd2556006},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd2556006},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd2556134},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd2556134},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd2556011},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd2556011},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd2556139},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd2556139},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd3604582},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd3604582},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd3604710},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd3604710},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd3604587},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd3604587},
'{step_type : POLL,	value : 32'd0,	reg_addr : 32'd3604715},
'{step_type : REG_WRITE,	value : 32'd2816,	reg_addr : 32'd3604715},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd458767},
'{step_type : REG_WRITE,	value : 32'd1,	reg_addr : 32'd851968}

}};
