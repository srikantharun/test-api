// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_v_center
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_v_center_p (
  output logic [41:0] o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld,
  input logic [7:0] i_sdma_0_init_tok_ocpl_s_maddr,
  input logic i_sdma_0_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_sdma_0_init_tok_ocpl_s_mdata,
  output logic  o_sdma_0_init_tok_ocpl_s_scmdaccept,
  output logic  o_sdma_0_pwr_tok_idle_val,
  output logic  o_sdma_0_pwr_tok_idle_ack,
  input logic  i_sdma_0_pwr_tok_idle_req,
  output logic [7:0] o_sdma_0_targ_tok_ocpl_m_maddr,
  output logic o_sdma_0_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_sdma_0_targ_tok_ocpl_m_mdata,
  input logic  i_sdma_0_targ_tok_ocpl_m_scmdaccept,
  input logic [7:0] i_sdma_1_init_tok_ocpl_s_maddr,
  input logic i_sdma_1_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_sdma_1_init_tok_ocpl_s_mdata,
  output logic  o_sdma_1_init_tok_ocpl_s_scmdaccept,
  output logic  o_sdma_1_pwr_tok_idle_val,
  output logic  o_sdma_1_pwr_tok_idle_ack,
  input logic  i_sdma_1_pwr_tok_idle_req,
  output logic [7:0] o_sdma_1_targ_tok_ocpl_m_maddr,
  output logic o_sdma_1_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_sdma_1_targ_tok_ocpl_m_mdata,
  input logic  i_sdma_1_targ_tok_ocpl_m_scmdaccept,

    output logic [686:0]                      o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld,
    output logic [182:0]                      o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld,
    input  logic [182:0]                      i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld,
    output logic [182:0]                      o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld,
    input  logic [182:0]                      i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld,
    output logic [182:0]                      o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld,
    input  logic [182:0]                      i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld,
    input  logic [182:0]                      i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld,
    output logic [182:0]                      o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld,
    input  logic [182:0]                      i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data,
    input  logic                              i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head,
    output logic                              o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy,
    input  logic                              i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail,
    input  logic                              i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld,
    output logic [182:0]                      o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data,
    output logic                              o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head,
    input  logic                              i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail,
    output logic                              o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld,
    input  logic [182:0]                      i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld,
    output logic [182:0]                      o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld,
    input  logic [182:0]                      i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld,
    output logic [182:0]                      o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld,
    input  logic                              i_l2_addr_mode_port_b0,
    input  logic                              i_l2_addr_mode_port_b1,
    input  logic                              i_l2_intr_mode_port_b0,
    input  logic                              i_l2_intr_mode_port_b1,
    input  logic                              i_lpddr_graph_addr_mode_port_b0,
    input  logic                              i_lpddr_graph_addr_mode_port_b1,
    input  logic                              i_lpddr_graph_intr_mode_port_b0,
    input  logic                              i_lpddr_graph_intr_mode_port_b1,
    input  logic                              i_lpddr_ppp_addr_mode_port_b0,
    input  logic                              i_lpddr_ppp_addr_mode_port_b1,
    input  logic                              i_lpddr_ppp_intr_mode_port_b0,
    input  logic                              i_lpddr_ppp_intr_mode_port_b1,
    input  wire                               i_noc_clk,
    input  wire                               i_noc_rst_n,
    input  wire                               i_sdma_0_aon_clk,
    input  wire                               i_sdma_0_aon_rst_n,
    input  wire                               i_sdma_0_clk,
    input  wire                               i_sdma_0_clken,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_ht_0_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_ht_0_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_ht_0_axi_s_arcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_0_init_ht_0_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_ht_0_axi_s_arlen,
    input  logic                              i_sdma_0_init_ht_0_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_ht_0_axi_s_arprot,
    output logic                              o_sdma_0_init_ht_0_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_ht_0_axi_s_arsize,
    input  logic                              i_sdma_0_init_ht_0_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t       o_sdma_0_init_ht_0_axi_s_rdata,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_0_init_ht_0_axi_s_rid,
    output logic                              o_sdma_0_init_ht_0_axi_s_rlast,
    input  logic                              i_sdma_0_init_ht_0_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_ht_0_axi_s_rresp,
    output logic                              o_sdma_0_init_ht_0_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_ht_0_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_ht_0_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_ht_0_axi_s_awcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_0_init_ht_0_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_ht_0_axi_s_awlen,
    input  logic                              i_sdma_0_init_ht_0_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_ht_0_axi_s_awprot,
    output logic                              o_sdma_0_init_ht_0_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_ht_0_axi_s_awsize,
    input  logic                              i_sdma_0_init_ht_0_axi_s_awvalid,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_0_init_ht_0_axi_s_bid,
    input  logic                              i_sdma_0_init_ht_0_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_ht_0_axi_s_bresp,
    output logic                              o_sdma_0_init_ht_0_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t       i_sdma_0_init_ht_0_axi_s_wdata,
    input  logic                              i_sdma_0_init_ht_0_axi_s_wlast,
    output logic                              o_sdma_0_init_ht_0_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t      i_sdma_0_init_ht_0_axi_s_wstrb,
    input  logic                              i_sdma_0_init_ht_0_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_ht_1_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_ht_1_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_ht_1_axi_s_arcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_0_init_ht_1_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_ht_1_axi_s_arlen,
    input  logic                              i_sdma_0_init_ht_1_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_ht_1_axi_s_arprot,
    output logic                              o_sdma_0_init_ht_1_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_ht_1_axi_s_arsize,
    input  logic                              i_sdma_0_init_ht_1_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t       o_sdma_0_init_ht_1_axi_s_rdata,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_0_init_ht_1_axi_s_rid,
    output logic                              o_sdma_0_init_ht_1_axi_s_rlast,
    input  logic                              i_sdma_0_init_ht_1_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_ht_1_axi_s_rresp,
    output logic                              o_sdma_0_init_ht_1_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_ht_1_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_ht_1_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_ht_1_axi_s_awcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_0_init_ht_1_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_ht_1_axi_s_awlen,
    input  logic                              i_sdma_0_init_ht_1_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_ht_1_axi_s_awprot,
    output logic                              o_sdma_0_init_ht_1_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_ht_1_axi_s_awsize,
    input  logic                              i_sdma_0_init_ht_1_axi_s_awvalid,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_0_init_ht_1_axi_s_bid,
    input  logic                              i_sdma_0_init_ht_1_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_ht_1_axi_s_bresp,
    output logic                              o_sdma_0_init_ht_1_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t       i_sdma_0_init_ht_1_axi_s_wdata,
    input  logic                              i_sdma_0_init_ht_1_axi_s_wlast,
    output logic                              o_sdma_0_init_ht_1_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t      i_sdma_0_init_ht_1_axi_s_wstrb,
    input  logic                              i_sdma_0_init_ht_1_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_lt_axi_s_arcache,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_0_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_lt_axi_s_arlen,
    input  logic                              i_sdma_0_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                 i_sdma_0_init_lt_axi_s_arqos,
    output logic                              o_sdma_0_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_lt_axi_s_arsize,
    input  logic                              i_sdma_0_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_lt_axi_s_awcache,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_0_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_lt_axi_s_awlen,
    input  logic                              i_sdma_0_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                 i_sdma_0_init_lt_axi_s_awqos,
    output logic                              o_sdma_0_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_lt_axi_s_awsize,
    input  logic                              i_sdma_0_init_lt_axi_s_awvalid,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_0_init_lt_axi_s_bid,
    input  logic                              i_sdma_0_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_lt_axi_s_bresp,
    output logic                              o_sdma_0_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t       o_sdma_0_init_lt_axi_s_rdata,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_0_init_lt_axi_s_rid,
    output logic                              o_sdma_0_init_lt_axi_s_rlast,
    input  logic                              i_sdma_0_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_lt_axi_s_rresp,
    output logic                              o_sdma_0_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t       i_sdma_0_init_lt_axi_s_wdata,
    input  logic                              i_sdma_0_init_lt_axi_s_wlast,
    output logic                              o_sdma_0_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t      i_sdma_0_init_lt_axi_s_wstrb,
    input  logic                              i_sdma_0_init_lt_axi_s_wvalid,
    output logic                              o_sdma_0_pwr_idle_val,
    output logic                              o_sdma_0_pwr_idle_ack,
    input  logic                              i_sdma_0_pwr_idle_req,
    input  wire                               i_sdma_0_rst_n,
    output chip_pkg::chip_axi_addr_t          o_sdma_0_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t               o_sdma_0_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t               o_sdma_0_targ_lt_axi_m_arcache,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_0_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                 o_sdma_0_targ_lt_axi_m_arlen,
    output logic                              o_sdma_0_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                o_sdma_0_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                 o_sdma_0_targ_lt_axi_m_arqos,
    input  logic                              i_sdma_0_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                o_sdma_0_targ_lt_axi_m_arsize,
    output logic                              o_sdma_0_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t          o_sdma_0_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t               o_sdma_0_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t               o_sdma_0_targ_lt_axi_m_awcache,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_0_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                 o_sdma_0_targ_lt_axi_m_awlen,
    output logic                              o_sdma_0_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                o_sdma_0_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                 o_sdma_0_targ_lt_axi_m_awqos,
    input  logic                              i_sdma_0_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                o_sdma_0_targ_lt_axi_m_awsize,
    output logic                              o_sdma_0_targ_lt_axi_m_awvalid,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_0_targ_lt_axi_m_bid,
    output logic                              o_sdma_0_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                i_sdma_0_targ_lt_axi_m_bresp,
    input  logic                              i_sdma_0_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t       i_sdma_0_targ_lt_axi_m_rdata,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_0_targ_lt_axi_m_rid,
    input  logic                              i_sdma_0_targ_lt_axi_m_rlast,
    output logic                              o_sdma_0_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                i_sdma_0_targ_lt_axi_m_rresp,
    input  logic                              i_sdma_0_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t       o_sdma_0_targ_lt_axi_m_wdata,
    output logic                              o_sdma_0_targ_lt_axi_m_wlast,
    input  logic                              i_sdma_0_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t      o_sdma_0_targ_lt_axi_m_wstrb,
    output logic                              o_sdma_0_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t       o_sdma_0_targ_syscfg_apb_m_paddr,
    output logic                              o_sdma_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t            o_sdma_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t   i_sdma_0_targ_syscfg_apb_m_prdata,
    input  logic                              i_sdma_0_targ_syscfg_apb_m_pready,
    output logic                              o_sdma_0_targ_syscfg_apb_m_psel,
    input  logic                              i_sdma_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t   o_sdma_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t   o_sdma_0_targ_syscfg_apb_m_pwdata,
    output logic                              o_sdma_0_targ_syscfg_apb_m_pwrite,
    input  wire                               i_sdma_1_aon_clk,
    input  wire                               i_sdma_1_aon_rst_n,
    input  wire                               i_sdma_1_clk,
    input  wire                               i_sdma_1_clken,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_ht_0_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_ht_0_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_ht_0_axi_s_arcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_1_init_ht_0_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_ht_0_axi_s_arlen,
    input  logic                              i_sdma_1_init_ht_0_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_ht_0_axi_s_arprot,
    output logic                              o_sdma_1_init_ht_0_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_ht_0_axi_s_arsize,
    input  logic                              i_sdma_1_init_ht_0_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t       o_sdma_1_init_ht_0_axi_s_rdata,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_1_init_ht_0_axi_s_rid,
    output logic                              o_sdma_1_init_ht_0_axi_s_rlast,
    input  logic                              i_sdma_1_init_ht_0_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_ht_0_axi_s_rresp,
    output logic                              o_sdma_1_init_ht_0_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_ht_0_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_ht_0_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_ht_0_axi_s_awcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_1_init_ht_0_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_ht_0_axi_s_awlen,
    input  logic                              i_sdma_1_init_ht_0_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_ht_0_axi_s_awprot,
    output logic                              o_sdma_1_init_ht_0_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_ht_0_axi_s_awsize,
    input  logic                              i_sdma_1_init_ht_0_axi_s_awvalid,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_1_init_ht_0_axi_s_bid,
    input  logic                              i_sdma_1_init_ht_0_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_ht_0_axi_s_bresp,
    output logic                              o_sdma_1_init_ht_0_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t       i_sdma_1_init_ht_0_axi_s_wdata,
    input  logic                              i_sdma_1_init_ht_0_axi_s_wlast,
    output logic                              o_sdma_1_init_ht_0_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t      i_sdma_1_init_ht_0_axi_s_wstrb,
    input  logic                              i_sdma_1_init_ht_0_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_ht_1_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_ht_1_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_ht_1_axi_s_arcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_1_init_ht_1_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_ht_1_axi_s_arlen,
    input  logic                              i_sdma_1_init_ht_1_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_ht_1_axi_s_arprot,
    output logic                              o_sdma_1_init_ht_1_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_ht_1_axi_s_arsize,
    input  logic                              i_sdma_1_init_ht_1_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t       o_sdma_1_init_ht_1_axi_s_rdata,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_1_init_ht_1_axi_s_rid,
    output logic                              o_sdma_1_init_ht_1_axi_s_rlast,
    input  logic                              i_sdma_1_init_ht_1_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_ht_1_axi_s_rresp,
    output logic                              o_sdma_1_init_ht_1_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_ht_1_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_ht_1_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_ht_1_axi_s_awcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_1_init_ht_1_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_ht_1_axi_s_awlen,
    input  logic                              i_sdma_1_init_ht_1_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_ht_1_axi_s_awprot,
    output logic                              o_sdma_1_init_ht_1_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_ht_1_axi_s_awsize,
    input  logic                              i_sdma_1_init_ht_1_axi_s_awvalid,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_1_init_ht_1_axi_s_bid,
    input  logic                              i_sdma_1_init_ht_1_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_ht_1_axi_s_bresp,
    output logic                              o_sdma_1_init_ht_1_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t       i_sdma_1_init_ht_1_axi_s_wdata,
    input  logic                              i_sdma_1_init_ht_1_axi_s_wlast,
    output logic                              o_sdma_1_init_ht_1_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t      i_sdma_1_init_ht_1_axi_s_wstrb,
    input  logic                              i_sdma_1_init_ht_1_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_lt_axi_s_arcache,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_1_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_lt_axi_s_arlen,
    input  logic                              i_sdma_1_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                 i_sdma_1_init_lt_axi_s_arqos,
    output logic                              o_sdma_1_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_lt_axi_s_arsize,
    input  logic                              i_sdma_1_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_lt_axi_s_awcache,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_1_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_lt_axi_s_awlen,
    input  logic                              i_sdma_1_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                 i_sdma_1_init_lt_axi_s_awqos,
    output logic                              o_sdma_1_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_lt_axi_s_awsize,
    input  logic                              i_sdma_1_init_lt_axi_s_awvalid,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_1_init_lt_axi_s_bid,
    input  logic                              i_sdma_1_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_lt_axi_s_bresp,
    output logic                              o_sdma_1_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t       o_sdma_1_init_lt_axi_s_rdata,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_1_init_lt_axi_s_rid,
    output logic                              o_sdma_1_init_lt_axi_s_rlast,
    input  logic                              i_sdma_1_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_lt_axi_s_rresp,
    output logic                              o_sdma_1_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t       i_sdma_1_init_lt_axi_s_wdata,
    input  logic                              i_sdma_1_init_lt_axi_s_wlast,
    output logic                              o_sdma_1_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t      i_sdma_1_init_lt_axi_s_wstrb,
    input  logic                              i_sdma_1_init_lt_axi_s_wvalid,
    output logic                              o_sdma_1_pwr_idle_val,
    output logic                              o_sdma_1_pwr_idle_ack,
    input  logic                              i_sdma_1_pwr_idle_req,
    input  wire                               i_sdma_1_rst_n,
    output chip_pkg::chip_axi_addr_t          o_sdma_1_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t               o_sdma_1_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t               o_sdma_1_targ_lt_axi_m_arcache,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_1_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                 o_sdma_1_targ_lt_axi_m_arlen,
    output logic                              o_sdma_1_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                o_sdma_1_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                 o_sdma_1_targ_lt_axi_m_arqos,
    input  logic                              i_sdma_1_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                o_sdma_1_targ_lt_axi_m_arsize,
    output logic                              o_sdma_1_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t          o_sdma_1_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t               o_sdma_1_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t               o_sdma_1_targ_lt_axi_m_awcache,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_1_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                 o_sdma_1_targ_lt_axi_m_awlen,
    output logic                              o_sdma_1_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                o_sdma_1_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                 o_sdma_1_targ_lt_axi_m_awqos,
    input  logic                              i_sdma_1_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                o_sdma_1_targ_lt_axi_m_awsize,
    output logic                              o_sdma_1_targ_lt_axi_m_awvalid,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_1_targ_lt_axi_m_bid,
    output logic                              o_sdma_1_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                i_sdma_1_targ_lt_axi_m_bresp,
    input  logic                              i_sdma_1_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t       i_sdma_1_targ_lt_axi_m_rdata,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_1_targ_lt_axi_m_rid,
    input  logic                              i_sdma_1_targ_lt_axi_m_rlast,
    output logic                              o_sdma_1_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                i_sdma_1_targ_lt_axi_m_rresp,
    input  logic                              i_sdma_1_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t       o_sdma_1_targ_lt_axi_m_wdata,
    output logic                              o_sdma_1_targ_lt_axi_m_wlast,
    input  logic                              i_sdma_1_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t      o_sdma_1_targ_lt_axi_m_wstrb,
    output logic                              o_sdma_1_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t       o_sdma_1_targ_syscfg_apb_m_paddr,
    output logic                              o_sdma_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t            o_sdma_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t   i_sdma_1_targ_syscfg_apb_m_prdata,
    input  logic                              i_sdma_1_targ_syscfg_apb_m_pready,
    output logic                              o_sdma_1_targ_syscfg_apb_m_psel,
    input  logic                              i_sdma_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t   o_sdma_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t   o_sdma_1_targ_syscfg_apb_m_pwdata,
    output logic                              o_sdma_1_targ_syscfg_apb_m_pwrite,
    // DFT Interface
    input  wire           tck,
    input  wire           trst,
    input  logic          tms,
    input  logic          tdi,
    output logic          tdo_en,
    output logic          tdo,
    input  wire           test_clk,
    input  logic          test_mode,
    input  logic          edt_update,
    input  logic          scan_en,
    input  logic [12-1:0] scan_in,
    output logic [12-1:0] scan_out
);

logic [2:0] sdma_0_targ_tok_ocpl_m_mcmd_ext;
assign o_sdma_0_targ_tok_ocpl_m_mcmd = sdma_0_targ_tok_ocpl_m_mcmd_ext[0];
logic [2:0] sdma_1_targ_tok_ocpl_m_mcmd_ext;
assign o_sdma_1_targ_tok_ocpl_m_mcmd = sdma_1_targ_tok_ocpl_m_mcmd_ext[0];


    // -- Automatically-generated Reset Synchronizers -- //
    wire sdma_0_aon_rst_n_synced;
    wire sdma_1_aon_rst_n_synced;

    // SDMA 0 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_sdma_0_aon_rst_n_sync (
        .i_clk          (i_sdma_0_aon_clk),
        .i_rst_n        (i_sdma_0_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (sdma_0_aon_rst_n_synced)
    );

    // SDMA 1 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_sdma_1_aon_rst_n_sync (
        .i_clk          (i_sdma_1_aon_clk),
        .i_rst_n        (i_sdma_1_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (sdma_1_aon_rst_n_synced)
    );

    noc_v_center u_noc_v_center (
    .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data),
    .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head),
    .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy),
    .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail),
    .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld),
    .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data),
    .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head),
    .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail),
    .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data),
    .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head),
    .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy),
    .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail),
    .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld),
    .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data),
    .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head),
    .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail),
    .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data),
    .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head),
    .i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy(i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail),
    .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld),
    .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data),
    .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head),
    .i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy(i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy),
    .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail),
    .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld),
    .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data),
    .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head),
    .o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy(o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data),
    .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head),
    .i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy(i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy),
    .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail),
    .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld),
    .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data),
    .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head),
    .o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy(o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy),
    .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail),
    .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld),
    .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data),
    .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head),
    .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy),
    .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail),
    .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld),
    .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data),
    .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head),
    .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy),
    .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail),
    .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld),
    .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data),
    .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head),
    .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy),
    .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail),
    .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld),
    .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data),
    .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head),
    .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy),
    .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail),
    .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld),
    .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data),
    .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head),
    .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy),
    .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail),
    .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld),
    .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data),
    .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head),
    .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy),
    .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail),
    .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld),
    .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data),
    .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head),
    .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy),
    .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail),
    .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld),
    .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data),
    .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head),
    .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy),
    .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail),
    .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld),
    .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data),
    .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head),
    .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy),
    .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail),
    .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld),
    .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data),
    .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head),
    .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy),
    .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail),
    .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld),
    .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data),
    .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head),
    .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy),
    .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail),
    .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld),
    .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data),
    .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head),
    .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data),
    .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head),
    .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy),
    .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail),
    .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld),
    .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data),
    .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head),
    .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data),
    .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head),
    .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy),
    .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail),
    .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld),
    .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data),
    .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head),
    .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy),
    .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail),
    .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data),
    .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head),
    .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail),
    .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld),
    .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data),
    .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head),
    .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail),
    .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld),
    .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data),
    .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head),
    .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail),
    .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld),
    .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data),
    .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head),
    .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail),
    .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld),
    .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data),
    .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head),
    .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail),
    .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld),
    .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data),
    .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head),
    .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail),
    .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld),
    .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data),
    .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head),
    .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail),
    .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld),
    .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data),
    .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head),
    .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail),
    .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld),
    .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data),
    .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head),
    .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail),
    .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld),
    .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data),
    .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head),
    .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail),
    .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld),
    .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data),
    .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head),
    .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail),
    .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld),
    .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data),
    .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head),
    .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy),
    .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail),
    .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld),
    .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data),
    .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head),
    .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data),
    .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head),
    .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy),
    .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail),
    .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld),
    .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data),
    .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head),
    .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy),
    .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail),
    .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data),
    .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head),
    .o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy(o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail),
    .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld),
    .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data),
    .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head),
    .o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy(o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail),
    .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld),
    .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data),
    .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head),
    .o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy(o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail),
    .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld),
    .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data),
    .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head),
    .o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy(o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail),
    .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld),
    .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data),
    .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head),
    .o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy(o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail),
    .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld),
    .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data),
    .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head),
    .o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy(o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail),
    .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld),
    .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data),
    .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head),
    .o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy(o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail),
    .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld),
    .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data),
    .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head),
    .o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy(o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail),
    .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld),
    .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data),
    .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head),
    .o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy(o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail),
    .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld),
    .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data),
    .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head),
    .o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy(o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail),
    .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld),
    .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data),
    .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head),
    .o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy(o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail),
    .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld),
    .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data),
    .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head),
    .o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy(o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy),
    .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail),
    .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld),
    .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data),
    .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head),
    .i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy(i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data),
    .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head),
    .o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy(o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy),
    .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail),
    .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld),
    .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data),
    .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head),
    .i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy(i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy),
    .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail),
    .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld),
    .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .i_noc_clk(i_noc_clk),
    .i_noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en),
    .i_sdma_0_aon_clk(i_sdma_0_aon_clk),
    .i_sdma_0_aon_rst_n(sdma_0_aon_rst_n_synced),
    .i_sdma_0_clk(i_sdma_0_clk),
    .i_sdma_0_clken(i_sdma_0_clken),
    .i_sdma_0_init_ht_0_axi_s_araddr(i_sdma_0_init_ht_0_axi_s_araddr),
    .i_sdma_0_init_ht_0_axi_s_arburst(i_sdma_0_init_ht_0_axi_s_arburst),
    .i_sdma_0_init_ht_0_axi_s_arcache(i_sdma_0_init_ht_0_axi_s_arcache),
    .i_sdma_0_init_ht_0_axi_s_arid(i_sdma_0_init_ht_0_axi_s_arid),
    .i_sdma_0_init_ht_0_axi_s_arlen(i_sdma_0_init_ht_0_axi_s_arlen),
    .i_sdma_0_init_ht_0_axi_s_arlock(i_sdma_0_init_ht_0_axi_s_arlock),
    .i_sdma_0_init_ht_0_axi_s_arprot(i_sdma_0_init_ht_0_axi_s_arprot),
    .o_sdma_0_init_ht_0_axi_s_arready(o_sdma_0_init_ht_0_axi_s_arready),
    .i_sdma_0_init_ht_0_axi_s_arsize(i_sdma_0_init_ht_0_axi_s_arsize),
    .i_sdma_0_init_ht_0_axi_s_arvalid(i_sdma_0_init_ht_0_axi_s_arvalid),
    .o_sdma_0_init_ht_0_axi_s_rdata(o_sdma_0_init_ht_0_axi_s_rdata),
    .o_sdma_0_init_ht_0_axi_s_rid(o_sdma_0_init_ht_0_axi_s_rid),
    .o_sdma_0_init_ht_0_axi_s_rlast(o_sdma_0_init_ht_0_axi_s_rlast),
    .i_sdma_0_init_ht_0_axi_s_rready(i_sdma_0_init_ht_0_axi_s_rready),
    .o_sdma_0_init_ht_0_axi_s_rresp(o_sdma_0_init_ht_0_axi_s_rresp),
    .o_sdma_0_init_ht_0_axi_s_rvalid(o_sdma_0_init_ht_0_axi_s_rvalid),
    .i_sdma_0_init_ht_0_axi_s_awaddr(i_sdma_0_init_ht_0_axi_s_awaddr),
    .i_sdma_0_init_ht_0_axi_s_awburst(i_sdma_0_init_ht_0_axi_s_awburst),
    .i_sdma_0_init_ht_0_axi_s_awcache(i_sdma_0_init_ht_0_axi_s_awcache),
    .i_sdma_0_init_ht_0_axi_s_awid(i_sdma_0_init_ht_0_axi_s_awid),
    .i_sdma_0_init_ht_0_axi_s_awlen(i_sdma_0_init_ht_0_axi_s_awlen),
    .i_sdma_0_init_ht_0_axi_s_awlock(i_sdma_0_init_ht_0_axi_s_awlock),
    .i_sdma_0_init_ht_0_axi_s_awprot(i_sdma_0_init_ht_0_axi_s_awprot),
    .o_sdma_0_init_ht_0_axi_s_awready(o_sdma_0_init_ht_0_axi_s_awready),
    .i_sdma_0_init_ht_0_axi_s_awsize(i_sdma_0_init_ht_0_axi_s_awsize),
    .i_sdma_0_init_ht_0_axi_s_awvalid(i_sdma_0_init_ht_0_axi_s_awvalid),
    .o_sdma_0_init_ht_0_axi_s_bid(o_sdma_0_init_ht_0_axi_s_bid),
    .i_sdma_0_init_ht_0_axi_s_bready(i_sdma_0_init_ht_0_axi_s_bready),
    .o_sdma_0_init_ht_0_axi_s_bresp(o_sdma_0_init_ht_0_axi_s_bresp),
    .o_sdma_0_init_ht_0_axi_s_bvalid(o_sdma_0_init_ht_0_axi_s_bvalid),
    .i_sdma_0_init_ht_0_axi_s_wdata(i_sdma_0_init_ht_0_axi_s_wdata),
    .i_sdma_0_init_ht_0_axi_s_wlast(i_sdma_0_init_ht_0_axi_s_wlast),
    .o_sdma_0_init_ht_0_axi_s_wready(o_sdma_0_init_ht_0_axi_s_wready),
    .i_sdma_0_init_ht_0_axi_s_wstrb(i_sdma_0_init_ht_0_axi_s_wstrb),
    .i_sdma_0_init_ht_0_axi_s_wvalid(i_sdma_0_init_ht_0_axi_s_wvalid),
    .i_sdma_0_init_ht_1_axi_s_araddr(i_sdma_0_init_ht_1_axi_s_araddr),
    .i_sdma_0_init_ht_1_axi_s_arburst(i_sdma_0_init_ht_1_axi_s_arburst),
    .i_sdma_0_init_ht_1_axi_s_arcache(i_sdma_0_init_ht_1_axi_s_arcache),
    .i_sdma_0_init_ht_1_axi_s_arid(i_sdma_0_init_ht_1_axi_s_arid),
    .i_sdma_0_init_ht_1_axi_s_arlen(i_sdma_0_init_ht_1_axi_s_arlen),
    .i_sdma_0_init_ht_1_axi_s_arlock(i_sdma_0_init_ht_1_axi_s_arlock),
    .i_sdma_0_init_ht_1_axi_s_arprot(i_sdma_0_init_ht_1_axi_s_arprot),
    .o_sdma_0_init_ht_1_axi_s_arready(o_sdma_0_init_ht_1_axi_s_arready),
    .i_sdma_0_init_ht_1_axi_s_arsize(i_sdma_0_init_ht_1_axi_s_arsize),
    .i_sdma_0_init_ht_1_axi_s_arvalid(i_sdma_0_init_ht_1_axi_s_arvalid),
    .o_sdma_0_init_ht_1_axi_s_rdata(o_sdma_0_init_ht_1_axi_s_rdata),
    .o_sdma_0_init_ht_1_axi_s_rid(o_sdma_0_init_ht_1_axi_s_rid),
    .o_sdma_0_init_ht_1_axi_s_rlast(o_sdma_0_init_ht_1_axi_s_rlast),
    .i_sdma_0_init_ht_1_axi_s_rready(i_sdma_0_init_ht_1_axi_s_rready),
    .o_sdma_0_init_ht_1_axi_s_rresp(o_sdma_0_init_ht_1_axi_s_rresp),
    .o_sdma_0_init_ht_1_axi_s_rvalid(o_sdma_0_init_ht_1_axi_s_rvalid),
    .i_sdma_0_init_ht_1_axi_s_awaddr(i_sdma_0_init_ht_1_axi_s_awaddr),
    .i_sdma_0_init_ht_1_axi_s_awburst(i_sdma_0_init_ht_1_axi_s_awburst),
    .i_sdma_0_init_ht_1_axi_s_awcache(i_sdma_0_init_ht_1_axi_s_awcache),
    .i_sdma_0_init_ht_1_axi_s_awid(i_sdma_0_init_ht_1_axi_s_awid),
    .i_sdma_0_init_ht_1_axi_s_awlen(i_sdma_0_init_ht_1_axi_s_awlen),
    .i_sdma_0_init_ht_1_axi_s_awlock(i_sdma_0_init_ht_1_axi_s_awlock),
    .i_sdma_0_init_ht_1_axi_s_awprot(i_sdma_0_init_ht_1_axi_s_awprot),
    .o_sdma_0_init_ht_1_axi_s_awready(o_sdma_0_init_ht_1_axi_s_awready),
    .i_sdma_0_init_ht_1_axi_s_awsize(i_sdma_0_init_ht_1_axi_s_awsize),
    .i_sdma_0_init_ht_1_axi_s_awvalid(i_sdma_0_init_ht_1_axi_s_awvalid),
    .o_sdma_0_init_ht_1_axi_s_bid(o_sdma_0_init_ht_1_axi_s_bid),
    .i_sdma_0_init_ht_1_axi_s_bready(i_sdma_0_init_ht_1_axi_s_bready),
    .o_sdma_0_init_ht_1_axi_s_bresp(o_sdma_0_init_ht_1_axi_s_bresp),
    .o_sdma_0_init_ht_1_axi_s_bvalid(o_sdma_0_init_ht_1_axi_s_bvalid),
    .i_sdma_0_init_ht_1_axi_s_wdata(i_sdma_0_init_ht_1_axi_s_wdata),
    .i_sdma_0_init_ht_1_axi_s_wlast(i_sdma_0_init_ht_1_axi_s_wlast),
    .o_sdma_0_init_ht_1_axi_s_wready(o_sdma_0_init_ht_1_axi_s_wready),
    .i_sdma_0_init_ht_1_axi_s_wstrb(i_sdma_0_init_ht_1_axi_s_wstrb),
    .i_sdma_0_init_ht_1_axi_s_wvalid(i_sdma_0_init_ht_1_axi_s_wvalid),
    .i_sdma_0_init_lt_axi_s_araddr(i_sdma_0_init_lt_axi_s_araddr),
    .i_sdma_0_init_lt_axi_s_arburst(i_sdma_0_init_lt_axi_s_arburst),
    .i_sdma_0_init_lt_axi_s_arcache(i_sdma_0_init_lt_axi_s_arcache),
    .i_sdma_0_init_lt_axi_s_arid(i_sdma_0_init_lt_axi_s_arid),
    .i_sdma_0_init_lt_axi_s_arlen(i_sdma_0_init_lt_axi_s_arlen),
    .i_sdma_0_init_lt_axi_s_arlock(i_sdma_0_init_lt_axi_s_arlock),
    .i_sdma_0_init_lt_axi_s_arprot(i_sdma_0_init_lt_axi_s_arprot),
    .i_sdma_0_init_lt_axi_s_arqos(i_sdma_0_init_lt_axi_s_arqos),
    .o_sdma_0_init_lt_axi_s_arready(o_sdma_0_init_lt_axi_s_arready),
    .i_sdma_0_init_lt_axi_s_arsize(i_sdma_0_init_lt_axi_s_arsize),
    .i_sdma_0_init_lt_axi_s_arvalid(i_sdma_0_init_lt_axi_s_arvalid),
    .i_sdma_0_init_lt_axi_s_awaddr(i_sdma_0_init_lt_axi_s_awaddr),
    .i_sdma_0_init_lt_axi_s_awburst(i_sdma_0_init_lt_axi_s_awburst),
    .i_sdma_0_init_lt_axi_s_awcache(i_sdma_0_init_lt_axi_s_awcache),
    .i_sdma_0_init_lt_axi_s_awid(i_sdma_0_init_lt_axi_s_awid),
    .i_sdma_0_init_lt_axi_s_awlen(i_sdma_0_init_lt_axi_s_awlen),
    .i_sdma_0_init_lt_axi_s_awlock(i_sdma_0_init_lt_axi_s_awlock),
    .i_sdma_0_init_lt_axi_s_awprot(i_sdma_0_init_lt_axi_s_awprot),
    .i_sdma_0_init_lt_axi_s_awqos(i_sdma_0_init_lt_axi_s_awqos),
    .o_sdma_0_init_lt_axi_s_awready(o_sdma_0_init_lt_axi_s_awready),
    .i_sdma_0_init_lt_axi_s_awsize(i_sdma_0_init_lt_axi_s_awsize),
    .i_sdma_0_init_lt_axi_s_awvalid(i_sdma_0_init_lt_axi_s_awvalid),
    .o_sdma_0_init_lt_axi_s_bid(o_sdma_0_init_lt_axi_s_bid),
    .i_sdma_0_init_lt_axi_s_bready(i_sdma_0_init_lt_axi_s_bready),
    .o_sdma_0_init_lt_axi_s_bresp(o_sdma_0_init_lt_axi_s_bresp),
    .o_sdma_0_init_lt_axi_s_bvalid(o_sdma_0_init_lt_axi_s_bvalid),
    .o_sdma_0_init_lt_axi_s_rdata(o_sdma_0_init_lt_axi_s_rdata),
    .o_sdma_0_init_lt_axi_s_rid(o_sdma_0_init_lt_axi_s_rid),
    .o_sdma_0_init_lt_axi_s_rlast(o_sdma_0_init_lt_axi_s_rlast),
    .i_sdma_0_init_lt_axi_s_rready(i_sdma_0_init_lt_axi_s_rready),
    .o_sdma_0_init_lt_axi_s_rresp(o_sdma_0_init_lt_axi_s_rresp),
    .o_sdma_0_init_lt_axi_s_rvalid(o_sdma_0_init_lt_axi_s_rvalid),
    .i_sdma_0_init_lt_axi_s_wdata(i_sdma_0_init_lt_axi_s_wdata),
    .i_sdma_0_init_lt_axi_s_wlast(i_sdma_0_init_lt_axi_s_wlast),
    .o_sdma_0_init_lt_axi_s_wready(o_sdma_0_init_lt_axi_s_wready),
    .i_sdma_0_init_lt_axi_s_wstrb(i_sdma_0_init_lt_axi_s_wstrb),
    .i_sdma_0_init_lt_axi_s_wvalid(i_sdma_0_init_lt_axi_s_wvalid),
    .o_sdma_0_pwr_idle_val(o_sdma_0_pwr_idle_val),
    .o_sdma_0_pwr_idle_ack(o_sdma_0_pwr_idle_ack),
    .i_sdma_0_pwr_idle_req(i_sdma_0_pwr_idle_req),
    .i_sdma_0_rst_n(i_sdma_0_rst_n),
    .o_sdma_0_targ_lt_axi_m_araddr(o_sdma_0_targ_lt_axi_m_araddr),
    .o_sdma_0_targ_lt_axi_m_arburst(o_sdma_0_targ_lt_axi_m_arburst),
    .o_sdma_0_targ_lt_axi_m_arcache(o_sdma_0_targ_lt_axi_m_arcache),
    .o_sdma_0_targ_lt_axi_m_arid(o_sdma_0_targ_lt_axi_m_arid),
    .o_sdma_0_targ_lt_axi_m_arlen(o_sdma_0_targ_lt_axi_m_arlen),
    .o_sdma_0_targ_lt_axi_m_arlock(o_sdma_0_targ_lt_axi_m_arlock),
    .o_sdma_0_targ_lt_axi_m_arprot(o_sdma_0_targ_lt_axi_m_arprot),
    .o_sdma_0_targ_lt_axi_m_arqos(o_sdma_0_targ_lt_axi_m_arqos),
    .i_sdma_0_targ_lt_axi_m_arready(i_sdma_0_targ_lt_axi_m_arready),
    .o_sdma_0_targ_lt_axi_m_arsize(o_sdma_0_targ_lt_axi_m_arsize),
    .o_sdma_0_targ_lt_axi_m_arvalid(o_sdma_0_targ_lt_axi_m_arvalid),
    .o_sdma_0_targ_lt_axi_m_awaddr(o_sdma_0_targ_lt_axi_m_awaddr),
    .o_sdma_0_targ_lt_axi_m_awburst(o_sdma_0_targ_lt_axi_m_awburst),
    .o_sdma_0_targ_lt_axi_m_awcache(o_sdma_0_targ_lt_axi_m_awcache),
    .o_sdma_0_targ_lt_axi_m_awid(o_sdma_0_targ_lt_axi_m_awid),
    .o_sdma_0_targ_lt_axi_m_awlen(o_sdma_0_targ_lt_axi_m_awlen),
    .o_sdma_0_targ_lt_axi_m_awlock(o_sdma_0_targ_lt_axi_m_awlock),
    .o_sdma_0_targ_lt_axi_m_awprot(o_sdma_0_targ_lt_axi_m_awprot),
    .o_sdma_0_targ_lt_axi_m_awqos(o_sdma_0_targ_lt_axi_m_awqos),
    .i_sdma_0_targ_lt_axi_m_awready(i_sdma_0_targ_lt_axi_m_awready),
    .o_sdma_0_targ_lt_axi_m_awsize(o_sdma_0_targ_lt_axi_m_awsize),
    .o_sdma_0_targ_lt_axi_m_awvalid(o_sdma_0_targ_lt_axi_m_awvalid),
    .i_sdma_0_targ_lt_axi_m_bid(i_sdma_0_targ_lt_axi_m_bid),
    .o_sdma_0_targ_lt_axi_m_bready(o_sdma_0_targ_lt_axi_m_bready),
    .i_sdma_0_targ_lt_axi_m_bresp(i_sdma_0_targ_lt_axi_m_bresp),
    .i_sdma_0_targ_lt_axi_m_bvalid(i_sdma_0_targ_lt_axi_m_bvalid),
    .i_sdma_0_targ_lt_axi_m_rdata(i_sdma_0_targ_lt_axi_m_rdata),
    .i_sdma_0_targ_lt_axi_m_rid(i_sdma_0_targ_lt_axi_m_rid),
    .i_sdma_0_targ_lt_axi_m_rlast(i_sdma_0_targ_lt_axi_m_rlast),
    .o_sdma_0_targ_lt_axi_m_rready(o_sdma_0_targ_lt_axi_m_rready),
    .i_sdma_0_targ_lt_axi_m_rresp(i_sdma_0_targ_lt_axi_m_rresp),
    .i_sdma_0_targ_lt_axi_m_rvalid(i_sdma_0_targ_lt_axi_m_rvalid),
    .o_sdma_0_targ_lt_axi_m_wdata(o_sdma_0_targ_lt_axi_m_wdata),
    .o_sdma_0_targ_lt_axi_m_wlast(o_sdma_0_targ_lt_axi_m_wlast),
    .i_sdma_0_targ_lt_axi_m_wready(i_sdma_0_targ_lt_axi_m_wready),
    .o_sdma_0_targ_lt_axi_m_wstrb(o_sdma_0_targ_lt_axi_m_wstrb),
    .o_sdma_0_targ_lt_axi_m_wvalid(o_sdma_0_targ_lt_axi_m_wvalid),
    .o_sdma_0_targ_syscfg_apb_m_paddr(o_sdma_0_targ_syscfg_apb_m_paddr),
    .o_sdma_0_targ_syscfg_apb_m_penable(o_sdma_0_targ_syscfg_apb_m_penable),
    .o_sdma_0_targ_syscfg_apb_m_pprot(o_sdma_0_targ_syscfg_apb_m_pprot),
    .i_sdma_0_targ_syscfg_apb_m_prdata(i_sdma_0_targ_syscfg_apb_m_prdata),
    .i_sdma_0_targ_syscfg_apb_m_pready(i_sdma_0_targ_syscfg_apb_m_pready),
    .o_sdma_0_targ_syscfg_apb_m_psel(o_sdma_0_targ_syscfg_apb_m_psel),
    .i_sdma_0_targ_syscfg_apb_m_pslverr(i_sdma_0_targ_syscfg_apb_m_pslverr),
    .o_sdma_0_targ_syscfg_apb_m_pstrb(o_sdma_0_targ_syscfg_apb_m_pstrb),
    .o_sdma_0_targ_syscfg_apb_m_pwdata(o_sdma_0_targ_syscfg_apb_m_pwdata),
    .o_sdma_0_targ_syscfg_apb_m_pwrite(o_sdma_0_targ_syscfg_apb_m_pwrite),
    .i_sdma_1_aon_clk(i_sdma_1_aon_clk),
    .i_sdma_1_aon_rst_n(sdma_1_aon_rst_n_synced),
    .i_sdma_1_clk(i_sdma_1_clk),
    .i_sdma_1_clken(i_sdma_1_clken),
    .i_sdma_1_init_ht_0_axi_s_araddr(i_sdma_1_init_ht_0_axi_s_araddr),
    .i_sdma_1_init_ht_0_axi_s_arburst(i_sdma_1_init_ht_0_axi_s_arburst),
    .i_sdma_1_init_ht_0_axi_s_arcache(i_sdma_1_init_ht_0_axi_s_arcache),
    .i_sdma_1_init_ht_0_axi_s_arid(i_sdma_1_init_ht_0_axi_s_arid),
    .i_sdma_1_init_ht_0_axi_s_arlen(i_sdma_1_init_ht_0_axi_s_arlen),
    .i_sdma_1_init_ht_0_axi_s_arlock(i_sdma_1_init_ht_0_axi_s_arlock),
    .i_sdma_1_init_ht_0_axi_s_arprot(i_sdma_1_init_ht_0_axi_s_arprot),
    .o_sdma_1_init_ht_0_axi_s_arready(o_sdma_1_init_ht_0_axi_s_arready),
    .i_sdma_1_init_ht_0_axi_s_arsize(i_sdma_1_init_ht_0_axi_s_arsize),
    .i_sdma_1_init_ht_0_axi_s_arvalid(i_sdma_1_init_ht_0_axi_s_arvalid),
    .o_sdma_1_init_ht_0_axi_s_rdata(o_sdma_1_init_ht_0_axi_s_rdata),
    .o_sdma_1_init_ht_0_axi_s_rid(o_sdma_1_init_ht_0_axi_s_rid),
    .o_sdma_1_init_ht_0_axi_s_rlast(o_sdma_1_init_ht_0_axi_s_rlast),
    .i_sdma_1_init_ht_0_axi_s_rready(i_sdma_1_init_ht_0_axi_s_rready),
    .o_sdma_1_init_ht_0_axi_s_rresp(o_sdma_1_init_ht_0_axi_s_rresp),
    .o_sdma_1_init_ht_0_axi_s_rvalid(o_sdma_1_init_ht_0_axi_s_rvalid),
    .i_sdma_1_init_ht_0_axi_s_awaddr(i_sdma_1_init_ht_0_axi_s_awaddr),
    .i_sdma_1_init_ht_0_axi_s_awburst(i_sdma_1_init_ht_0_axi_s_awburst),
    .i_sdma_1_init_ht_0_axi_s_awcache(i_sdma_1_init_ht_0_axi_s_awcache),
    .i_sdma_1_init_ht_0_axi_s_awid(i_sdma_1_init_ht_0_axi_s_awid),
    .i_sdma_1_init_ht_0_axi_s_awlen(i_sdma_1_init_ht_0_axi_s_awlen),
    .i_sdma_1_init_ht_0_axi_s_awlock(i_sdma_1_init_ht_0_axi_s_awlock),
    .i_sdma_1_init_ht_0_axi_s_awprot(i_sdma_1_init_ht_0_axi_s_awprot),
    .o_sdma_1_init_ht_0_axi_s_awready(o_sdma_1_init_ht_0_axi_s_awready),
    .i_sdma_1_init_ht_0_axi_s_awsize(i_sdma_1_init_ht_0_axi_s_awsize),
    .i_sdma_1_init_ht_0_axi_s_awvalid(i_sdma_1_init_ht_0_axi_s_awvalid),
    .o_sdma_1_init_ht_0_axi_s_bid(o_sdma_1_init_ht_0_axi_s_bid),
    .i_sdma_1_init_ht_0_axi_s_bready(i_sdma_1_init_ht_0_axi_s_bready),
    .o_sdma_1_init_ht_0_axi_s_bresp(o_sdma_1_init_ht_0_axi_s_bresp),
    .o_sdma_1_init_ht_0_axi_s_bvalid(o_sdma_1_init_ht_0_axi_s_bvalid),
    .i_sdma_1_init_ht_0_axi_s_wdata(i_sdma_1_init_ht_0_axi_s_wdata),
    .i_sdma_1_init_ht_0_axi_s_wlast(i_sdma_1_init_ht_0_axi_s_wlast),
    .o_sdma_1_init_ht_0_axi_s_wready(o_sdma_1_init_ht_0_axi_s_wready),
    .i_sdma_1_init_ht_0_axi_s_wstrb(i_sdma_1_init_ht_0_axi_s_wstrb),
    .i_sdma_1_init_ht_0_axi_s_wvalid(i_sdma_1_init_ht_0_axi_s_wvalid),
    .i_sdma_1_init_ht_1_axi_s_araddr(i_sdma_1_init_ht_1_axi_s_araddr),
    .i_sdma_1_init_ht_1_axi_s_arburst(i_sdma_1_init_ht_1_axi_s_arburst),
    .i_sdma_1_init_ht_1_axi_s_arcache(i_sdma_1_init_ht_1_axi_s_arcache),
    .i_sdma_1_init_ht_1_axi_s_arid(i_sdma_1_init_ht_1_axi_s_arid),
    .i_sdma_1_init_ht_1_axi_s_arlen(i_sdma_1_init_ht_1_axi_s_arlen),
    .i_sdma_1_init_ht_1_axi_s_arlock(i_sdma_1_init_ht_1_axi_s_arlock),
    .i_sdma_1_init_ht_1_axi_s_arprot(i_sdma_1_init_ht_1_axi_s_arprot),
    .o_sdma_1_init_ht_1_axi_s_arready(o_sdma_1_init_ht_1_axi_s_arready),
    .i_sdma_1_init_ht_1_axi_s_arsize(i_sdma_1_init_ht_1_axi_s_arsize),
    .i_sdma_1_init_ht_1_axi_s_arvalid(i_sdma_1_init_ht_1_axi_s_arvalid),
    .o_sdma_1_init_ht_1_axi_s_rdata(o_sdma_1_init_ht_1_axi_s_rdata),
    .o_sdma_1_init_ht_1_axi_s_rid(o_sdma_1_init_ht_1_axi_s_rid),
    .o_sdma_1_init_ht_1_axi_s_rlast(o_sdma_1_init_ht_1_axi_s_rlast),
    .i_sdma_1_init_ht_1_axi_s_rready(i_sdma_1_init_ht_1_axi_s_rready),
    .o_sdma_1_init_ht_1_axi_s_rresp(o_sdma_1_init_ht_1_axi_s_rresp),
    .o_sdma_1_init_ht_1_axi_s_rvalid(o_sdma_1_init_ht_1_axi_s_rvalid),
    .i_sdma_1_init_ht_1_axi_s_awaddr(i_sdma_1_init_ht_1_axi_s_awaddr),
    .i_sdma_1_init_ht_1_axi_s_awburst(i_sdma_1_init_ht_1_axi_s_awburst),
    .i_sdma_1_init_ht_1_axi_s_awcache(i_sdma_1_init_ht_1_axi_s_awcache),
    .i_sdma_1_init_ht_1_axi_s_awid(i_sdma_1_init_ht_1_axi_s_awid),
    .i_sdma_1_init_ht_1_axi_s_awlen(i_sdma_1_init_ht_1_axi_s_awlen),
    .i_sdma_1_init_ht_1_axi_s_awlock(i_sdma_1_init_ht_1_axi_s_awlock),
    .i_sdma_1_init_ht_1_axi_s_awprot(i_sdma_1_init_ht_1_axi_s_awprot),
    .o_sdma_1_init_ht_1_axi_s_awready(o_sdma_1_init_ht_1_axi_s_awready),
    .i_sdma_1_init_ht_1_axi_s_awsize(i_sdma_1_init_ht_1_axi_s_awsize),
    .i_sdma_1_init_ht_1_axi_s_awvalid(i_sdma_1_init_ht_1_axi_s_awvalid),
    .o_sdma_1_init_ht_1_axi_s_bid(o_sdma_1_init_ht_1_axi_s_bid),
    .i_sdma_1_init_ht_1_axi_s_bready(i_sdma_1_init_ht_1_axi_s_bready),
    .o_sdma_1_init_ht_1_axi_s_bresp(o_sdma_1_init_ht_1_axi_s_bresp),
    .o_sdma_1_init_ht_1_axi_s_bvalid(o_sdma_1_init_ht_1_axi_s_bvalid),
    .i_sdma_1_init_ht_1_axi_s_wdata(i_sdma_1_init_ht_1_axi_s_wdata),
    .i_sdma_1_init_ht_1_axi_s_wlast(i_sdma_1_init_ht_1_axi_s_wlast),
    .o_sdma_1_init_ht_1_axi_s_wready(o_sdma_1_init_ht_1_axi_s_wready),
    .i_sdma_1_init_ht_1_axi_s_wstrb(i_sdma_1_init_ht_1_axi_s_wstrb),
    .i_sdma_1_init_ht_1_axi_s_wvalid(i_sdma_1_init_ht_1_axi_s_wvalid),
    .i_sdma_1_init_lt_axi_s_araddr(i_sdma_1_init_lt_axi_s_araddr),
    .i_sdma_1_init_lt_axi_s_arburst(i_sdma_1_init_lt_axi_s_arburst),
    .i_sdma_1_init_lt_axi_s_arcache(i_sdma_1_init_lt_axi_s_arcache),
    .i_sdma_1_init_lt_axi_s_arid(i_sdma_1_init_lt_axi_s_arid),
    .i_sdma_1_init_lt_axi_s_arlen(i_sdma_1_init_lt_axi_s_arlen),
    .i_sdma_1_init_lt_axi_s_arlock(i_sdma_1_init_lt_axi_s_arlock),
    .i_sdma_1_init_lt_axi_s_arprot(i_sdma_1_init_lt_axi_s_arprot),
    .i_sdma_1_init_lt_axi_s_arqos(i_sdma_1_init_lt_axi_s_arqos),
    .o_sdma_1_init_lt_axi_s_arready(o_sdma_1_init_lt_axi_s_arready),
    .i_sdma_1_init_lt_axi_s_arsize(i_sdma_1_init_lt_axi_s_arsize),
    .i_sdma_1_init_lt_axi_s_arvalid(i_sdma_1_init_lt_axi_s_arvalid),
    .i_sdma_1_init_lt_axi_s_awaddr(i_sdma_1_init_lt_axi_s_awaddr),
    .i_sdma_1_init_lt_axi_s_awburst(i_sdma_1_init_lt_axi_s_awburst),
    .i_sdma_1_init_lt_axi_s_awcache(i_sdma_1_init_lt_axi_s_awcache),
    .i_sdma_1_init_lt_axi_s_awid(i_sdma_1_init_lt_axi_s_awid),
    .i_sdma_1_init_lt_axi_s_awlen(i_sdma_1_init_lt_axi_s_awlen),
    .i_sdma_1_init_lt_axi_s_awlock(i_sdma_1_init_lt_axi_s_awlock),
    .i_sdma_1_init_lt_axi_s_awprot(i_sdma_1_init_lt_axi_s_awprot),
    .i_sdma_1_init_lt_axi_s_awqos(i_sdma_1_init_lt_axi_s_awqos),
    .o_sdma_1_init_lt_axi_s_awready(o_sdma_1_init_lt_axi_s_awready),
    .i_sdma_1_init_lt_axi_s_awsize(i_sdma_1_init_lt_axi_s_awsize),
    .i_sdma_1_init_lt_axi_s_awvalid(i_sdma_1_init_lt_axi_s_awvalid),
    .o_sdma_1_init_lt_axi_s_bid(o_sdma_1_init_lt_axi_s_bid),
    .i_sdma_1_init_lt_axi_s_bready(i_sdma_1_init_lt_axi_s_bready),
    .o_sdma_1_init_lt_axi_s_bresp(o_sdma_1_init_lt_axi_s_bresp),
    .o_sdma_1_init_lt_axi_s_bvalid(o_sdma_1_init_lt_axi_s_bvalid),
    .o_sdma_1_init_lt_axi_s_rdata(o_sdma_1_init_lt_axi_s_rdata),
    .o_sdma_1_init_lt_axi_s_rid(o_sdma_1_init_lt_axi_s_rid),
    .o_sdma_1_init_lt_axi_s_rlast(o_sdma_1_init_lt_axi_s_rlast),
    .i_sdma_1_init_lt_axi_s_rready(i_sdma_1_init_lt_axi_s_rready),
    .o_sdma_1_init_lt_axi_s_rresp(o_sdma_1_init_lt_axi_s_rresp),
    .o_sdma_1_init_lt_axi_s_rvalid(o_sdma_1_init_lt_axi_s_rvalid),
    .i_sdma_1_init_lt_axi_s_wdata(i_sdma_1_init_lt_axi_s_wdata),
    .i_sdma_1_init_lt_axi_s_wlast(i_sdma_1_init_lt_axi_s_wlast),
    .o_sdma_1_init_lt_axi_s_wready(o_sdma_1_init_lt_axi_s_wready),
    .i_sdma_1_init_lt_axi_s_wstrb(i_sdma_1_init_lt_axi_s_wstrb),
    .i_sdma_1_init_lt_axi_s_wvalid(i_sdma_1_init_lt_axi_s_wvalid),
    .o_sdma_1_pwr_idle_val(o_sdma_1_pwr_idle_val),
    .o_sdma_1_pwr_idle_ack(o_sdma_1_pwr_idle_ack),
    .i_sdma_1_pwr_idle_req(i_sdma_1_pwr_idle_req),
    .i_sdma_1_rst_n(i_sdma_1_rst_n),
    .o_sdma_1_targ_lt_axi_m_araddr(o_sdma_1_targ_lt_axi_m_araddr),
    .o_sdma_1_targ_lt_axi_m_arburst(o_sdma_1_targ_lt_axi_m_arburst),
    .o_sdma_1_targ_lt_axi_m_arcache(o_sdma_1_targ_lt_axi_m_arcache),
    .o_sdma_1_targ_lt_axi_m_arid(o_sdma_1_targ_lt_axi_m_arid),
    .o_sdma_1_targ_lt_axi_m_arlen(o_sdma_1_targ_lt_axi_m_arlen),
    .o_sdma_1_targ_lt_axi_m_arlock(o_sdma_1_targ_lt_axi_m_arlock),
    .o_sdma_1_targ_lt_axi_m_arprot(o_sdma_1_targ_lt_axi_m_arprot),
    .o_sdma_1_targ_lt_axi_m_arqos(o_sdma_1_targ_lt_axi_m_arqos),
    .i_sdma_1_targ_lt_axi_m_arready(i_sdma_1_targ_lt_axi_m_arready),
    .o_sdma_1_targ_lt_axi_m_arsize(o_sdma_1_targ_lt_axi_m_arsize),
    .o_sdma_1_targ_lt_axi_m_arvalid(o_sdma_1_targ_lt_axi_m_arvalid),
    .o_sdma_1_targ_lt_axi_m_awaddr(o_sdma_1_targ_lt_axi_m_awaddr),
    .o_sdma_1_targ_lt_axi_m_awburst(o_sdma_1_targ_lt_axi_m_awburst),
    .o_sdma_1_targ_lt_axi_m_awcache(o_sdma_1_targ_lt_axi_m_awcache),
    .o_sdma_1_targ_lt_axi_m_awid(o_sdma_1_targ_lt_axi_m_awid),
    .o_sdma_1_targ_lt_axi_m_awlen(o_sdma_1_targ_lt_axi_m_awlen),
    .o_sdma_1_targ_lt_axi_m_awlock(o_sdma_1_targ_lt_axi_m_awlock),
    .o_sdma_1_targ_lt_axi_m_awprot(o_sdma_1_targ_lt_axi_m_awprot),
    .o_sdma_1_targ_lt_axi_m_awqos(o_sdma_1_targ_lt_axi_m_awqos),
    .i_sdma_1_targ_lt_axi_m_awready(i_sdma_1_targ_lt_axi_m_awready),
    .o_sdma_1_targ_lt_axi_m_awsize(o_sdma_1_targ_lt_axi_m_awsize),
    .o_sdma_1_targ_lt_axi_m_awvalid(o_sdma_1_targ_lt_axi_m_awvalid),
    .i_sdma_1_targ_lt_axi_m_bid(i_sdma_1_targ_lt_axi_m_bid),
    .o_sdma_1_targ_lt_axi_m_bready(o_sdma_1_targ_lt_axi_m_bready),
    .i_sdma_1_targ_lt_axi_m_bresp(i_sdma_1_targ_lt_axi_m_bresp),
    .i_sdma_1_targ_lt_axi_m_bvalid(i_sdma_1_targ_lt_axi_m_bvalid),
    .i_sdma_1_targ_lt_axi_m_rdata(i_sdma_1_targ_lt_axi_m_rdata),
    .i_sdma_1_targ_lt_axi_m_rid(i_sdma_1_targ_lt_axi_m_rid),
    .i_sdma_1_targ_lt_axi_m_rlast(i_sdma_1_targ_lt_axi_m_rlast),
    .o_sdma_1_targ_lt_axi_m_rready(o_sdma_1_targ_lt_axi_m_rready),
    .i_sdma_1_targ_lt_axi_m_rresp(i_sdma_1_targ_lt_axi_m_rresp),
    .i_sdma_1_targ_lt_axi_m_rvalid(i_sdma_1_targ_lt_axi_m_rvalid),
    .o_sdma_1_targ_lt_axi_m_wdata(o_sdma_1_targ_lt_axi_m_wdata),
    .o_sdma_1_targ_lt_axi_m_wlast(o_sdma_1_targ_lt_axi_m_wlast),
    .i_sdma_1_targ_lt_axi_m_wready(i_sdma_1_targ_lt_axi_m_wready),
    .o_sdma_1_targ_lt_axi_m_wstrb(o_sdma_1_targ_lt_axi_m_wstrb),
    .o_sdma_1_targ_lt_axi_m_wvalid(o_sdma_1_targ_lt_axi_m_wvalid),
    .o_sdma_1_targ_syscfg_apb_m_paddr(o_sdma_1_targ_syscfg_apb_m_paddr),
    .o_sdma_1_targ_syscfg_apb_m_penable(o_sdma_1_targ_syscfg_apb_m_penable),
    .o_sdma_1_targ_syscfg_apb_m_pprot(o_sdma_1_targ_syscfg_apb_m_pprot),
    .i_sdma_1_targ_syscfg_apb_m_prdata(i_sdma_1_targ_syscfg_apb_m_prdata),
    .i_sdma_1_targ_syscfg_apb_m_pready(i_sdma_1_targ_syscfg_apb_m_pready),
    .o_sdma_1_targ_syscfg_apb_m_psel(o_sdma_1_targ_syscfg_apb_m_psel),
    .i_sdma_1_targ_syscfg_apb_m_pslverr(i_sdma_1_targ_syscfg_apb_m_pslverr),
    .o_sdma_1_targ_syscfg_apb_m_pstrb(o_sdma_1_targ_syscfg_apb_m_pstrb),
    .o_sdma_1_targ_syscfg_apb_m_pwdata(o_sdma_1_targ_syscfg_apb_m_pwdata),
    .o_sdma_1_targ_syscfg_apb_m_pwrite(o_sdma_1_targ_syscfg_apb_m_pwrite)
);

noc_tok_v_center u_noc_tok_v_center (
  .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data),
  .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head),
  .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy),
  .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail),
  .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld),
  .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data),
  .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head),
  .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy),
  .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail),
  .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld),
  .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data),
  .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head),
  .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy),
  .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail),
  .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld),
  .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data),
  .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head),
  .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy),
  .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail),
  .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld),
  .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data),
  .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head),
  .i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy(i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy),
  .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail),
  .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld),
  .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data),
  .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head),
  .i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy(i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy),
  .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail),
  .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld),
  .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data),
  .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head),
  .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy),
  .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail),
  .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld),
  .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data),
  .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head),
  .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy),
  .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail),
  .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld),
  .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data),
  .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head),
  .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy),
  .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail),
  .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld),
  .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data),
  .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head),
  .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy),
  .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail),
  .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld),
  .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data),
  .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head),
  .o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy(o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy),
  .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail),
  .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld),
  .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data),
  .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head),
  .o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy(o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy),
  .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail),
  .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld),
  .i_noc_clk(i_noc_clk),
  .i_noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en),
  .i_sdma_0_clk(i_sdma_0_clk),
  .i_sdma_0_clken(i_sdma_0_clken),
  .i_sdma_0_init_tok_ocpl_s_maddr(i_sdma_0_init_tok_ocpl_s_maddr),
  .i_sdma_0_init_tok_ocpl_s_mcmd({{ 2'b0, i_sdma_0_init_tok_ocpl_s_mcmd }}),
  .i_sdma_0_init_tok_ocpl_s_mdata(i_sdma_0_init_tok_ocpl_s_mdata),
  .o_sdma_0_init_tok_ocpl_s_scmdaccept(o_sdma_0_init_tok_ocpl_s_scmdaccept),
  .o_sdma_0_pwr_tok_idle_val(o_sdma_0_pwr_tok_idle_val),
  .o_sdma_0_pwr_tok_idle_ack(o_sdma_0_pwr_tok_idle_ack),
  .i_sdma_0_pwr_tok_idle_req(i_sdma_0_pwr_tok_idle_req),
  .i_sdma_0_rst_n(i_sdma_0_rst_n),
  .o_sdma_0_targ_tok_ocpl_m_maddr(o_sdma_0_targ_tok_ocpl_m_maddr),
  .o_sdma_0_targ_tok_ocpl_m_mcmd(sdma_0_targ_tok_ocpl_m_mcmd_ext),
  .o_sdma_0_targ_tok_ocpl_m_mdata(o_sdma_0_targ_tok_ocpl_m_mdata),
  .i_sdma_0_targ_tok_ocpl_m_scmdaccept(i_sdma_0_targ_tok_ocpl_m_scmdaccept),
  .i_sdma_1_clk(i_sdma_1_clk),
  .i_sdma_1_clken(i_sdma_1_clken),
  .i_sdma_1_init_tok_ocpl_s_maddr(i_sdma_1_init_tok_ocpl_s_maddr),
  .i_sdma_1_init_tok_ocpl_s_mcmd({{ 2'b0, i_sdma_1_init_tok_ocpl_s_mcmd }}),
  .i_sdma_1_init_tok_ocpl_s_mdata(i_sdma_1_init_tok_ocpl_s_mdata),
  .o_sdma_1_init_tok_ocpl_s_scmdaccept(o_sdma_1_init_tok_ocpl_s_scmdaccept),
  .o_sdma_1_pwr_tok_idle_val(o_sdma_1_pwr_tok_idle_val),
  .o_sdma_1_pwr_tok_idle_ack(o_sdma_1_pwr_tok_idle_ack),
  .i_sdma_1_pwr_tok_idle_req(i_sdma_1_pwr_tok_idle_req),
  .i_sdma_1_rst_n(i_sdma_1_rst_n),
  .o_sdma_1_targ_tok_ocpl_m_maddr(o_sdma_1_targ_tok_ocpl_m_maddr),
  .o_sdma_1_targ_tok_ocpl_m_mcmd(sdma_1_targ_tok_ocpl_m_mcmd_ext),
  .o_sdma_1_targ_tok_ocpl_m_mdata(o_sdma_1_targ_tok_ocpl_m_mdata),
  .i_sdma_1_targ_tok_ocpl_m_scmdaccept(i_sdma_1_targ_tok_ocpl_m_scmdaccept)
);
endmodule
