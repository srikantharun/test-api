// *** (C) Copyright Axelera AI 2021        *** //
// *** All Rights Reserved                  *** //
// *** Axelera AI Confidential              *** //
// *** Owner : srinivas.prakash@axelera.ai  *** //

`ifndef GUARD_ENOC_TB_INTF_SV
`define GUARD_ENOC_TB_INTF_SV
// User defined interface to control the power    //
// domain fences and other misc signals from test //
interface enoc_tb_intf();

  logic enoc_clk                          ;
  logic enoc_rst_n                        ;
  logic noc_slow_clk                      ;
  logic noc_slow_rst_n                    ;
  logic interleave_mode_select_port       ;
  logic address_scheme_select_port        ;
  logic noc_irq_0                         ;
  bit o_aic_0_pwr_tok_idle_val            ;
  bit o_aic_0_pwr_tok_idle_ack            ;
  bit i_aic_0_pwr_tok_idle_req            ;
  bit o_aic_1_pwr_tok_idle_val            ;
  bit o_aic_1_pwr_tok_idle_ack            ;
  bit i_aic_1_pwr_tok_idle_req            ;
  bit o_aic_2_pwr_tok_idle_val            ;
  bit o_aic_2_pwr_tok_idle_ack            ;
  bit i_aic_2_pwr_tok_idle_req            ;
  bit o_aic_3_pwr_tok_idle_val            ;
  bit o_aic_3_pwr_tok_idle_ack            ;
  bit i_aic_3_pwr_tok_idle_req            ;
  bit o_aic_4_pwr_tok_idle_val            ;
  bit o_aic_4_pwr_tok_idle_ack            ;
  bit i_aic_4_pwr_tok_idle_req            ;
  bit o_aic_5_pwr_tok_idle_val            ;
  bit o_aic_5_pwr_tok_idle_ack            ;
  bit i_aic_5_pwr_tok_idle_req            ;
  bit o_aic_6_pwr_tok_idle_val            ;
  bit o_aic_6_pwr_tok_idle_ack            ;
  bit i_aic_6_pwr_tok_idle_req            ;
  bit o_aic_7_pwr_tok_idle_val            ;
  bit o_aic_7_pwr_tok_idle_ack            ;
  bit i_aic_7_pwr_tok_idle_req            ;
  bit o_apu_pwr_tok_idle_val              ;
  bit o_apu_pwr_tok_idle_ack              ;
  bit i_apu_pwr_tok_idle_req              ;
  bit i_aic_0_pwr_idle_req                ;
  bit i_aic_1_pwr_idle_req                ;
  bit i_aic_2_pwr_idle_req                ;
  bit i_aic_3_pwr_idle_req                ;
  bit i_aic_4_pwr_idle_req                ;
  bit i_aic_5_pwr_idle_req                ;
  bit i_aic_6_pwr_idle_req                ;
  bit i_aic_7_pwr_idle_req                ;
  bit i_apu_pwr_idle_req                  ;
  bit i_dcd_mcu_pwr_idle_req              ;
  bit i_dcd_pwr_idle_req                  ;
  bit i_l2_0_pwr_idle_req                 ;
  bit i_l2_1_pwr_idle_req                 ;
  bit i_l2_2_pwr_idle_req                 ;
  bit i_l2_3_pwr_idle_req                 ;
  bit i_l2_4_pwr_idle_req                 ;
  bit i_l2_5_pwr_idle_req                 ;
  bit i_l2_6_pwr_idle_req                 ;
  bit i_l2_7_pwr_idle_req                 ;
  bit[1:0] i_lpddr_graph_0_pwr_idle_vec_req        ;
  bit[1:0] i_lpddr_graph_1_pwr_idle_vec_req        ;
  bit[1:0] i_lpddr_graph_2_pwr_idle_vec_req        ;
  bit[1:0] i_lpddr_graph_3_pwr_idle_vec_req        ;
  bit[1:0] i_lpddr_ppp_0_pwr_idle_vec_req          ;
  bit[1:0] i_lpddr_ppp_1_pwr_idle_vec_req          ;
  bit[1:0] i_lpddr_ppp_2_pwr_idle_vec_req          ;
  bit[1:0] i_lpddr_ppp_3_pwr_idle_vec_req          ;
  bit i_pcie_init_mt_pwr_idle_req                 ;
  bit i_pcie_targ_mt_pwr_idle_req                 ;
  bit i_pcie_targ_cfg_pwr_idle_req                 ;
  bit i_pcie_targ_cfg_dbi_pwr_idle_req                 ;
  bit i_pve_0_pwr_idle_req                ;
  bit i_pve_1_pwr_idle_req                ;
  bit i_soc_mgmt_pwr_idle_req             ;
  bit i_soc_periph_pwr_idle_req           ;
  bit i_sys_spm_pwr_idle_req              ;
  bit o_aic_0_pwr_idle_val                ;
  bit o_aic_1_pwr_idle_val                ;
  bit o_aic_2_pwr_idle_val                ;
  bit o_aic_3_pwr_idle_val                ;
  bit o_aic_4_pwr_idle_val                ;
  bit o_aic_5_pwr_idle_val                ;
  bit o_aic_6_pwr_idle_val                ;
  bit o_aic_7_pwr_idle_val                ;
  bit o_apu_pwr_idle_val                  ;
  bit o_dcd_mcu_pwr_idle_val              ;
  bit o_dcd_pwr_idle_val                  ;
  bit o_l2_0_pwr_idle_val                 ;
  bit o_l2_1_pwr_idle_val                 ;
  bit o_l2_2_pwr_idle_val                 ;
  bit o_l2_3_pwr_idle_val                 ;
  bit o_l2_4_pwr_idle_val                 ;
  bit o_l2_5_pwr_idle_val                 ;
  bit o_l2_6_pwr_idle_val                 ;
  bit o_l2_7_pwr_idle_val                 ;
  bit[1:0] o_lpddr_graph_0_pwr_idle_vec_val        ;
  bit[1:0] o_lpddr_graph_1_pwr_idle_vec_val        ;
  bit[1:0] o_lpddr_graph_2_pwr_idle_vec_val        ;
  bit[1:0] o_lpddr_graph_3_pwr_idle_vec_val        ;
  bit[1:0] o_lpddr_ppp_0_pwr_idle_vec_val          ;
  bit[1:0] o_lpddr_ppp_1_pwr_idle_vec_val          ;
  bit[1:0] o_lpddr_ppp_2_pwr_idle_vec_val          ;
  bit[1:0] o_lpddr_ppp_3_pwr_idle_vec_val          ;
  bit o_pcie_init_mt_pwr_idle_val                 ;
  bit o_pcie_targ_mt_pwr_idle_val                 ;
  bit o_pcie_targ_cfg_pwr_idle_val                 ;
  bit o_pcie_targ_cfg_dbi_pwr_idle_val                 ;
  bit o_pve_0_pwr_idle_val                ;
  bit o_pve_1_pwr_idle_val                ;
  bit o_soc_mgmt_pwr_idle_val             ;
  bit o_soc_periph_pwr_idle_val           ;
  bit o_sys_spm_pwr_idle_val              ;
  bit o_aic_0_pwr_idle_ack                ;
  bit o_aic_1_pwr_idle_ack                ;
  bit o_aic_2_pwr_idle_ack                ;
  bit o_aic_3_pwr_idle_ack                ;
  bit o_aic_4_pwr_idle_ack                ;
  bit o_aic_5_pwr_idle_ack                ;
  bit o_aic_6_pwr_idle_ack                ;
  bit o_aic_7_pwr_idle_ack                ;
  bit o_apu_pwr_idle_ack                  ;
  bit o_dcd_mcu_pwr_idle_ack              ;
  bit o_dcd_pwr_idle_ack                  ;
  bit o_l2_0_pwr_idle_ack                 ;
  bit o_l2_1_pwr_idle_ack                 ;
  bit o_l2_2_pwr_idle_ack                 ;
  bit o_l2_3_pwr_idle_ack                 ;
  bit o_l2_4_pwr_idle_ack                 ;
  bit o_l2_5_pwr_idle_ack                 ;
  bit o_l2_6_pwr_idle_ack                 ;
  bit o_l2_7_pwr_idle_ack                 ;
  bit[1:0] o_lpddr_graph_0_pwr_idle_vec_ack        ;
  bit[1:0] o_lpddr_graph_1_pwr_idle_vec_ack        ;
  bit[1:0] o_lpddr_graph_2_pwr_idle_vec_ack        ;
  bit[1:0] o_lpddr_graph_3_pwr_idle_vec_ack        ;
  bit[1:0] o_lpddr_ppp_0_pwr_idle_vec_ack          ;
  bit[1:0] o_lpddr_ppp_1_pwr_idle_vec_ack          ;
  bit[1:0] o_lpddr_ppp_2_pwr_idle_vec_ack          ;
  bit[1:0] o_lpddr_ppp_3_pwr_idle_vec_ack          ;
  bit o_pcie_init_mt_pwr_idle_ack                 ;
  bit o_pcie_targ_mt_pwr_idle_ack                 ;
  bit o_pcie_targ_cfg_pwr_idle_ack                 ;
  bit o_pcie_targ_cfg_dbi_pwr_idle_ack                 ;
  bit o_pve_0_pwr_idle_ack                ;
  bit o_pve_1_pwr_idle_ack                ;
  bit o_soc_mgmt_pwr_idle_ack           ;
  bit o_soc_periph_pwr_idle_ack           ;
  bit o_sys_spm_pwr_idle_ack              ;
  bit[7:0] i_aic_0_init_tok_ocpl_s_maddr  ;
  bit i_aic_0_init_tok_ocpl_s_mcmd        ;
  bit[7:0] i_aic_0_init_tok_ocpl_s_mdata  ;
  bit o_aic_0_init_tok_ocpl_s_scmdaccept  ;
  bit[7:0] o_aic_0_targ_tok_ocpl_m_maddr  ;
  bit o_aic_0_targ_tok_ocpl_m_mcmd        ;
  bit[7:0] o_aic_0_targ_tok_ocpl_m_mdata  ;
  bit i_aic_0_targ_tok_ocpl_m_scmdaccept  ;
  bit[7:0] i_aic_1_init_tok_ocpl_s_maddr  ;
  bit i_aic_1_init_tok_ocpl_s_mcmd        ;
  bit[7:0] i_aic_1_init_tok_ocpl_s_mdata  ;
  bit o_aic_1_init_tok_ocpl_s_scmdaccept  ;
  bit[7:0] o_aic_1_targ_tok_ocpl_m_maddr  ;
  bit o_aic_1_targ_tok_ocpl_m_mcmd        ;
  bit[7:0] o_aic_1_targ_tok_ocpl_m_mdata  ;
  bit i_aic_1_targ_tok_ocpl_m_scmdaccept  ;
  bit[7:0] i_aic_2_init_tok_ocpl_s_maddr  ;
  bit i_aic_2_init_tok_ocpl_s_mcmd        ;
  bit[7:0] i_aic_2_init_tok_ocpl_s_mdata  ;
  bit o_aic_2_init_tok_ocpl_s_scmdaccept  ;
  bit[7:0] o_aic_2_targ_tok_ocpl_m_maddr  ;
  bit o_aic_2_targ_tok_ocpl_m_mcmd        ;
  bit[7:0] o_aic_2_targ_tok_ocpl_m_mdata  ;
  bit i_aic_2_targ_tok_ocpl_m_scmdaccept  ;
  bit[7:0] i_aic_3_init_tok_ocpl_s_maddr  ;
  bit i_aic_3_init_tok_ocpl_s_mcmd        ;
  bit[7:0] i_aic_3_init_tok_ocpl_s_mdata  ;
  bit o_aic_3_init_tok_ocpl_s_scmdaccept  ;
  bit[7:0] o_aic_3_targ_tok_ocpl_m_maddr  ;
  bit o_aic_3_targ_tok_ocpl_m_mcmd        ;
  bit[7:0] o_aic_3_targ_tok_ocpl_m_mdata  ;
  bit i_aic_3_targ_tok_ocpl_m_scmdaccept  ;
  bit[7:0] i_aic_4_init_tok_ocpl_s_maddr  ;
  bit i_aic_4_init_tok_ocpl_s_mcmd        ;
  bit[7:0] i_aic_4_init_tok_ocpl_s_mdata  ;
  bit o_aic_4_init_tok_ocpl_s_scmdaccept  ;
  bit[7:0] o_aic_4_targ_tok_ocpl_m_maddr  ;
  bit o_aic_4_targ_tok_ocpl_m_mcmd        ;
  bit[7:0] o_aic_4_targ_tok_ocpl_m_mdata  ;
  bit i_aic_4_targ_tok_ocpl_m_scmdaccept  ;
  bit[7:0] i_aic_5_init_tok_ocpl_s_maddr  ;
  bit i_aic_5_init_tok_ocpl_s_mcmd        ;
  bit[7:0] i_aic_5_init_tok_ocpl_s_mdata  ;
  bit o_aic_5_init_tok_ocpl_s_scmdaccept  ;
  bit[7:0] o_aic_5_targ_tok_ocpl_m_maddr  ;
  bit o_aic_5_targ_tok_ocpl_m_mcmd        ;
  bit[7:0] o_aic_5_targ_tok_ocpl_m_mdata  ;
  bit i_aic_5_targ_tok_ocpl_m_scmdaccept  ;
  bit[7:0] i_aic_6_init_tok_ocpl_s_maddr  ;
  bit i_aic_6_init_tok_ocpl_s_mcmd        ;
  bit[7:0] i_aic_6_init_tok_ocpl_s_mdata  ;
  bit o_aic_6_init_tok_ocpl_s_scmdaccept  ;
  bit[7:0] o_aic_6_targ_tok_ocpl_m_maddr  ;
  bit o_aic_6_targ_tok_ocpl_m_mcmd        ;
  bit[7:0] o_aic_6_targ_tok_ocpl_m_mdata  ;
  bit i_aic_6_targ_tok_ocpl_m_scmdaccept  ;
  bit[7:0] i_aic_7_init_tok_ocpl_s_maddr  ;
  bit i_aic_7_init_tok_ocpl_s_mcmd        ;
  bit[7:0] i_aic_7_init_tok_ocpl_s_mdata  ;
  bit o_aic_7_init_tok_ocpl_s_scmdaccept  ;
  bit[7:0] o_aic_7_targ_tok_ocpl_m_maddr  ;
  bit o_aic_7_targ_tok_ocpl_m_mcmd        ;
  bit[7:0] o_aic_7_targ_tok_ocpl_m_mdata  ;
  bit i_aic_7_targ_tok_ocpl_m_scmdaccept  ;
  bit[7:0] i_apu_init_tok_ocpl_s_maddr    ;
  bit i_apu_init_tok_ocpl_s_mcmd          ;
  bit[7:0] i_apu_init_tok_ocpl_s_mdata    ;
  bit o_apu_init_tok_ocpl_s_scmdaccept    ;
  bit[7:0] o_apu_targ_tok_ocpl_m_maddr    ;
  bit o_apu_targ_tok_ocpl_m_mcmd          ;
  bit[7:0] o_apu_targ_tok_ocpl_m_mdata    ;
  bit i_apu_targ_tok_ocpl_m_scmdaccept    ;
endinterface : enoc_tb_intf
`endif // GUARD_ENOC_TB_INTF_SV
