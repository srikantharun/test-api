//noc_init_hp_ai_core_3

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (9),
				.WID_WIDTH  (9),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_hp_I_ai_core_0
				(
				.ACLK(aic_0_clk),
				.ARESETn(aic_0_rst_n),
				.ARVALID(ai_core_0_init_hp_I_axi_m_arvalid),
				.ARADDR(ai_core_0_init_hp_I_axi_m_araddr ),
				.ARLEN(ai_core_0_init_hp_I_axi_m_arlen),
				.ARSIZE( ai_core_0_init_hp_I_axi_m_arsize),
				.ARBURST( ai_core_0_init_hp_I_axi_m_arburst ),
				.ARLOCK( ai_core_0_init_hp_I_axi_m_arlock),
				.ARCACHE( ai_core_0_init_hp_I_axi_m_arcache ),
				.ARPROT( ai_core_0_init_hp_I_axi_m_arprot ),
				.ARID( ai_core_0_init_hp_I_axi_m_arid ),
				.ARREADY( ai_core_0_init_hp_I_axi_m_arready ),
				.RREADY( ai_core_0_init_hp_I_axi_m_rready ),
				.RVALID( ai_core_0_init_hp_I_axi_m_rvalid ),
				.RLAST( ai_core_0_init_hp_I_axi_m_rlast ),
				.RDATA({ ai_core_0_init_hp_I_axi_m_rdata } ),
				.RRESP( ai_core_0_init_hp_I_axi_m_rresp ),
				.RID( ai_core_0_init_hp_I_axi_m_rid ),
				.AWVALID( ai_core_0_init_hp_I_axi_m_awvalid ),
				.AWADDR( ai_core_0_init_hp_I_axi_m_awaddr ),
				.AWLEN( ai_core_0_init_hp_I_axi_m_awlen),
				.AWSIZE( ai_core_0_init_hp_I_axi_m_awsize ),
				.AWBURST( ai_core_0_init_hp_I_axi_m_awburst ),
				.AWLOCK( ai_core_0_init_hp_I_axi_m_awlock ),
				.AWCACHE( ai_core_0_init_hp_I_axi_m_awcache ),
				.AWPROT( ai_core_0_init_hp_I_axi_m_awprot ),
				.AWID( ai_core_0_init_hp_I_axi_m_awid ),
				.AWREADY( ai_core_0_init_hp_I_axi_m_awready ),
				.WVALID( ai_core_0_init_hp_I_axi_m_wvalid ),
				.WLAST( ai_core_0_init_hp_I_axi_m_wlast ),
				.WDATA(  ai_core_0_init_hp_I_axi_m_wdata ),
				.WSTRB( ai_core_0_init_hp_I_axi_m_wstrb ),
				.WREADY( ai_core_0_init_hp_I_axi_m_wready),
				.BREADY( ai_core_0_init_hp_I_axi_m_bready ),
				.BVALID( ai_core_0_init_hp_I_axi_m_bvalid ),
				.BRESP( ai_core_0_init_hp_I_axi_m_bresp ),
				.BID( ai_core_0_init_hp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

//noc_init_lp_ai_core_0
bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (9),
				.WID_WIDTH  (9),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_lp_I_ai_core_0
				(
				.ACLK(aic_0_clk),
				.ARESETn(aic_0_rst_n),
				.ARVALID(ai_core_0_init_lp_I_axi_m_arvalid),
				.ARADDR(ai_core_0_init_lp_I_axi_m_araddr ),
				.ARLEN(ai_core_0_init_lp_I_axi_m_arlen),
				.ARSIZE( ai_core_0_init_lp_I_axi_m_arsize),
				.ARBURST( ai_core_0_init_lp_I_axi_m_arburst ),
				.ARLOCK( ai_core_0_init_lp_I_axi_m_arlock),
				.ARCACHE( ai_core_0_init_lp_I_axi_m_arcache ),
				.ARPROT( ai_core_0_init_lp_I_axi_m_arprot ),
				.ARID( ai_core_0_init_lp_I_axi_m_arid ),
				.ARREADY( ai_core_0_init_lp_I_axi_m_arready ),
				.RREADY( ai_core_0_init_lp_I_axi_m_rready ),
				.RVALID( ai_core_0_init_lp_I_axi_m_rvalid ),
				.RLAST( ai_core_0_init_lp_I_axi_m_rlast ),
				.RDATA( ai_core_0_init_lp_I_axi_m_rdata ),
				.RRESP( ai_core_0_init_lp_I_axi_m_rresp ),
				.RID( ai_core_0_init_lp_I_axi_m_rid ),
				.AWVALID( ai_core_0_init_lp_I_axi_m_awvalid ),
				.AWADDR( ai_core_0_init_lp_I_axi_m_awaddr ),
				.AWLEN( ai_core_0_init_lp_I_axi_m_awlen),
				.AWSIZE( ai_core_0_init_lp_I_axi_m_awsize ),
				.AWBURST( ai_core_0_init_lp_I_axi_m_awburst ),
				.AWLOCK( ai_core_0_init_lp_I_axi_m_awlock ),
				.AWCACHE( ai_core_0_init_lp_I_axi_m_awcache ),
				.AWPROT( ai_core_0_init_lp_I_axi_m_awprot ),
				.AWID( ai_core_0_init_lp_I_axi_m_awid ),
				.AWREADY( ai_core_0_init_lp_I_axi_m_awready ),
				.WVALID( ai_core_0_init_lp_I_axi_m_wvalid ),
				.WLAST( ai_core_0_init_lp_I_axi_m_wlast ),
				.WDATA(  ai_core_0_init_lp_I_axi_m_wdata ),
				.WSTRB( ai_core_0_init_lp_I_axi_m_wstrb ),
				.WREADY( ai_core_0_init_lp_I_axi_m_wready),
				.BREADY( ai_core_0_init_lp_I_axi_m_bready ),
				.BVALID( ai_core_0_init_lp_I_axi_m_bvalid ),
				.BRESP( ai_core_0_init_lp_I_axi_m_bresp ),
				.BID( ai_core_0_init_lp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//// noc_Targ_lp_ai_core_0

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_targ_lp_I_ai_core_0
				(
				.ACLK(aic_0_clk),
				.ARESETn(aic_0_rst_n),
				.ARVALID(ai_core_0_targ_lp_T_axi_s_arvalid),
				.ARADDR(ai_core_0_targ_lp_T_axi_s_araddr ),
				.ARLEN(ai_core_0_targ_lp_T_axi_s_arlen),
				.ARSIZE( ai_core_0_targ_lp_T_axi_s_arsize),
				.ARBURST( ai_core_0_targ_lp_T_axi_s_arburst ),
				.ARLOCK( ai_core_0_targ_lp_T_axi_s_arlock),
				.ARCACHE( ai_core_0_targ_lp_T_axi_s_arcache ),
				.ARPROT( ai_core_0_targ_lp_T_axi_s_arprot ),
				.ARID( ai_core_0_targ_lp_T_axi_s_arid ),
				.ARREADY( ai_core_0_targ_lp_T_axi_s_arready ),
				.RREADY( ai_core_0_targ_lp_T_axi_s_rready ),
				.RVALID( ai_core_0_targ_lp_T_axi_s_rvalid ),
				.RLAST( ai_core_0_targ_lp_T_axi_s_rlast ),
				.RDATA(  ai_core_0_targ_lp_T_axi_s_rdata ),
				.RRESP( ai_core_0_targ_lp_T_axi_s_rresp ),
				.RID( ai_core_0_targ_lp_T_axi_s_rid ),
				.AWVALID( ai_core_0_targ_lp_T_axi_s_awvalid ),
				.AWADDR( ai_core_0_targ_lp_T_axi_s_awaddr ),
				.AWLEN( ai_core_0_targ_lp_T_axi_s_awlen),
				.AWSIZE( ai_core_0_targ_lp_T_axi_s_awsize ),
				.AWBURST( ai_core_0_targ_lp_T_axi_s_awburst ),
				.AWLOCK( ai_core_0_targ_lp_T_axi_s_awlock ),
				.AWCACHE( ai_core_0_targ_lp_T_axi_s_awcache ),
				.AWPROT( ai_core_0_targ_lp_T_axi_s_awprot ),
				.AWID( ai_core_0_targ_lp_T_axi_s_awid ),
				.AWREADY( ai_core_0_targ_lp_T_axi_s_awready ),
				.WVALID( ai_core_0_targ_lp_T_axi_s_wvalid ),
				.WLAST( ai_core_0_targ_lp_T_axi_s_wlast ),
				.WDATA(  ai_core_0_targ_lp_T_axi_s_wdata ),
				.WSTRB( ai_core_0_targ_lp_T_axi_s_wstrb ),
				.WREADY( ai_core_0_targ_lp_T_axi_s_wready),
				.BREADY( ai_core_0_targ_lp_T_axi_s_bready ),
				.BVALID( ai_core_0_targ_lp_T_axi_s_bvalid ),
				.BRESP( ai_core_0_targ_lp_T_axi_s_bresp ),
				.BID( ai_core_0_targ_lp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//noc_triton_ai_hp_core_1
bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (9),
				.WID_WIDTH  (9),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_hp_I_ai_core_1
				(
				.ACLK(aic_1_clk),
				.ARESETn(aic_1_rst_n),
				.ARVALID(ai_core_1_init_hp_I_axi_m_arvalid),
				.ARADDR(ai_core_1_init_hp_I_axi_m_araddr ),
				.ARLEN(ai_core_1_init_hp_I_axi_m_arlen),
				.ARSIZE( ai_core_1_init_hp_I_axi_m_arsize),
				.ARBURST( ai_core_1_init_hp_I_axi_m_arburst ),
				.ARLOCK( ai_core_1_init_hp_I_axi_m_arlock),
				.ARCACHE( ai_core_1_init_hp_I_axi_m_arcache ),
				.ARPROT( ai_core_1_init_hp_I_axi_m_arprot ),
				.ARID( ai_core_1_init_hp_I_axi_m_arid ),
				.ARREADY( ai_core_1_init_hp_I_axi_m_arready ),
				.RREADY( ai_core_1_init_hp_I_axi_m_rready ),
				.RVALID( ai_core_1_init_hp_I_axi_m_rvalid ),
				.RLAST( ai_core_1_init_hp_I_axi_m_rlast ),
				.RDATA(  ai_core_1_init_hp_I_axi_m_rdata ),
				.RRESP( ai_core_1_init_hp_I_axi_m_rresp ),
				.RID( ai_core_1_init_hp_I_axi_m_rid ),
				.AWVALID( ai_core_1_init_hp_I_axi_m_awvalid ),
				.AWADDR( ai_core_1_init_hp_I_axi_m_awaddr ),
				.AWLEN( ai_core_1_init_hp_I_axi_m_awlen),
				.AWSIZE( ai_core_1_init_hp_I_axi_m_awsize ),
				.AWBURST( ai_core_1_init_hp_I_axi_m_awburst ),
				.AWLOCK( ai_core_1_init_hp_I_axi_m_awlock ),
				.AWCACHE( ai_core_1_init_hp_I_axi_m_awcache ),
				.AWPROT( ai_core_1_init_hp_I_axi_m_awprot ),
				.AWID( ai_core_1_init_hp_I_axi_m_awid ),
				.AWREADY( ai_core_1_init_hp_I_axi_m_awready ),
				.WVALID( ai_core_1_init_hp_I_axi_m_wvalid ),
				.WLAST( ai_core_1_init_hp_I_axi_m_wlast ),
				.WDATA(  ai_core_1_init_hp_I_axi_m_wdata ),
				.WSTRB( ai_core_1_init_hp_I_axi_m_wstrb ),
				.WREADY( ai_core_1_init_hp_I_axi_m_wready),
				.BREADY( ai_core_1_init_hp_I_axi_m_bready ),
				.BVALID( ai_core_1_init_hp_I_axi_m_bvalid ),
				.BRESP( ai_core_1_init_hp_I_axi_m_bresp ),
				.BID( ai_core_1_init_hp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

//noc_init_lp_ai_core_1
bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (9),
				.WID_WIDTH  (9),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_lp_I_ai_core_1
				(
				.ACLK(aic_1_clk),
				.ARESETn(aic_1_rst_n),
				.ARVALID(ai_core_1_init_lp_I_axi_m_arvalid),
				.ARADDR(ai_core_1_init_lp_I_axi_m_araddr ),
				.ARLEN(ai_core_1_init_lp_I_axi_m_arlen),
				.ARSIZE( ai_core_1_init_lp_I_axi_m_arsize),
				.ARBURST( ai_core_1_init_lp_I_axi_m_arburst ),
				.ARLOCK( ai_core_1_init_lp_I_axi_m_arlock),
				.ARCACHE( ai_core_1_init_lp_I_axi_m_arcache ),
				.ARPROT( ai_core_1_init_lp_I_axi_m_arprot ),
				.ARID( ai_core_1_init_lp_I_axi_m_arid ),
				.ARREADY( ai_core_1_init_lp_I_axi_m_arready ),
				.RREADY( ai_core_1_init_lp_I_axi_m_rready ),
				.RVALID( ai_core_1_init_lp_I_axi_m_rvalid ),
				.RLAST( ai_core_1_init_lp_I_axi_m_rlast ),
				.RDATA(  ai_core_1_init_lp_I_axi_m_rdata ),
				.RRESP( ai_core_1_init_lp_I_axi_m_rresp ),
				.RID( ai_core_1_init_lp_I_axi_m_rid ),
				.AWVALID( ai_core_1_init_lp_I_axi_m_awvalid ),
				.AWADDR( ai_core_1_init_lp_I_axi_m_awaddr ),
				.AWLEN( ai_core_1_init_lp_I_axi_m_awlen),
				.AWSIZE( ai_core_1_init_lp_I_axi_m_awsize ),
				.AWBURST( ai_core_1_init_lp_I_axi_m_awburst ),
				.AWLOCK( ai_core_1_init_lp_I_axi_m_awlock ),
				.AWCACHE( ai_core_1_init_lp_I_axi_m_awcache ),
				.AWPROT( ai_core_1_init_lp_I_axi_m_awprot ),
				.AWID( ai_core_1_init_lp_I_axi_m_awid ),
				.AWREADY( ai_core_1_init_lp_I_axi_m_awready ),
				.WVALID( ai_core_1_init_lp_I_axi_m_wvalid ),
				.WLAST( ai_core_1_init_lp_I_axi_m_wlast ),
				.WDATA(  ai_core_1_init_lp_I_axi_m_wdata ),
				.WSTRB( ai_core_1_init_lp_I_axi_m_wstrb ),
				.WREADY( ai_core_1_init_lp_I_axi_m_wready),
				.BREADY( ai_core_1_init_lp_I_axi_m_bready ),
				.BVALID( ai_core_1_init_lp_I_axi_m_bvalid ),
				.BRESP( ai_core_1_init_lp_I_axi_m_bresp ),
				.BID( ai_core_1_init_lp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//// noc_Targ_lp_ai_core_1

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_targ_lp_I_ai_core_1
				(
				.ACLK(aic_1_clk),
				.ARESETn(aic_1_rst_n),
				.ARVALID(ai_core_1_targ_lp_T_axi_s_arvalid),
				.ARADDR(ai_core_1_targ_lp_T_axi_s_araddr ),
				.ARLEN(ai_core_1_targ_lp_T_axi_s_arlen),
				.ARSIZE( ai_core_1_targ_lp_T_axi_s_arsize),
				.ARBURST( ai_core_1_targ_lp_T_axi_s_arburst ),
				.ARLOCK( ai_core_1_targ_lp_T_axi_s_arlock),
				.ARCACHE( ai_core_1_targ_lp_T_axi_s_arcache ),
				.ARPROT( ai_core_1_targ_lp_T_axi_s_arprot ),
				.ARID( ai_core_1_targ_lp_T_axi_s_arid ),
				.ARREADY( ai_core_1_targ_lp_T_axi_s_arready ),
				.RREADY( ai_core_1_targ_lp_T_axi_s_rready ),
				.RVALID( ai_core_1_targ_lp_T_axi_s_rvalid ),
				.RLAST( ai_core_1_targ_lp_T_axi_s_rlast ),
				.RDATA(  ai_core_1_targ_lp_T_axi_s_rdata ),
				.RRESP( ai_core_1_targ_lp_T_axi_s_rresp ),
				.RID( ai_core_1_targ_lp_T_axi_s_rid ),
				.AWVALID( ai_core_1_targ_lp_T_axi_s_awvalid ),
				.AWADDR( ai_core_1_targ_lp_T_axi_s_awaddr ),
				.AWLEN( ai_core_1_targ_lp_T_axi_s_awlen),
				.AWSIZE( ai_core_1_targ_lp_T_axi_s_awsize ),
				.AWBURST( ai_core_1_targ_lp_T_axi_s_awburst ),
				.AWLOCK( ai_core_1_targ_lp_T_axi_s_awlock ),
				.AWCACHE( ai_core_1_targ_lp_T_axi_s_awcache ),
				.AWPROT( ai_core_1_targ_lp_T_axi_s_awprot ),
				.AWID( ai_core_1_targ_lp_T_axi_s_awid ),
				.AWREADY( ai_core_1_targ_lp_T_axi_s_awready ),
				.WVALID( ai_core_1_targ_lp_T_axi_s_wvalid ),
				.WLAST( ai_core_1_targ_lp_T_axi_s_wlast ),
				.WDATA(  ai_core_1_targ_lp_T_axi_s_wdata ),
				.WSTRB( ai_core_1_targ_lp_T_axi_s_wstrb ),
				.WREADY( ai_core_1_targ_lp_T_axi_s_wready),
				.BREADY( ai_core_1_targ_lp_T_axi_s_bready ),
				.BVALID( ai_core_1_targ_lp_T_axi_s_bvalid ),
				.BRESP( ai_core_1_targ_lp_T_axi_s_bresp ),
				.BID( ai_core_1_targ_lp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//noc_triton_hp_ai_core_2

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (9),
				.WID_WIDTH  (9),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_hp_I_ai_core_2
				(
				.ACLK(aic_2_clk),
				.ARESETn(aic_2_rst_n),
				.ARVALID(ai_core_2_init_hp_I_axi_m_arvalid),
				.ARADDR(ai_core_2_init_hp_I_axi_m_araddr ),
				.ARLEN(ai_core_2_init_hp_I_axi_m_arlen),
				.ARSIZE( ai_core_2_init_hp_I_axi_m_arsize),
				.ARBURST( ai_core_2_init_hp_I_axi_m_arburst ),
				.ARLOCK( ai_core_2_init_hp_I_axi_m_arlock),
				.ARCACHE( ai_core_2_init_hp_I_axi_m_arcache ),
				.ARPROT( ai_core_2_init_hp_I_axi_m_arprot ),
				.ARID( ai_core_2_init_hp_I_axi_m_arid ),
				.ARREADY( ai_core_2_init_hp_I_axi_m_arready ),
				.RREADY( ai_core_2_init_hp_I_axi_m_rready ),
				.RVALID( ai_core_2_init_hp_I_axi_m_rvalid ),
				.RLAST( ai_core_2_init_hp_I_axi_m_rlast ),
				.RDATA(  ai_core_2_init_hp_I_axi_m_rdata ),
				.RRESP( ai_core_2_init_hp_I_axi_m_rresp ),
				.RID( ai_core_2_init_hp_I_axi_m_rid ),
				.AWVALID( ai_core_2_init_hp_I_axi_m_awvalid ),
				.AWADDR( ai_core_2_init_hp_I_axi_m_awaddr ),
				.AWLEN( ai_core_2_init_hp_I_axi_m_awlen),
				.AWSIZE( ai_core_2_init_hp_I_axi_m_awsize ),
				.AWBURST( ai_core_2_init_hp_I_axi_m_awburst ),
				.AWLOCK( ai_core_2_init_hp_I_axi_m_awlock ),
				.AWCACHE( ai_core_2_init_hp_I_axi_m_awcache ),
				.AWPROT( ai_core_2_init_hp_I_axi_m_awprot ),
				.AWID( ai_core_2_init_hp_I_axi_m_awid ),
				.AWREADY( ai_core_2_init_hp_I_axi_m_awready ),
				.WVALID( ai_core_2_init_hp_I_axi_m_wvalid ),
				.WLAST( ai_core_2_init_hp_I_axi_m_wlast ),
				.WDATA(  ai_core_2_init_hp_I_axi_m_wdata ),
				.WSTRB( ai_core_2_init_hp_I_axi_m_wstrb ),
				.WREADY( ai_core_2_init_hp_I_axi_m_wready),
				.BREADY( ai_core_2_init_hp_I_axi_m_bready ),
				.BVALID( ai_core_2_init_hp_I_axi_m_bvalid ),
				.BRESP( ai_core_2_init_hp_I_axi_m_bresp ),
				.BID( ai_core_2_init_hp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

//noc_init_lp_ai_core_2
bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (9),
				.WID_WIDTH  (9),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_lp_I_ai_core_2
				(
				.ACLK(aic_2_clk),
				.ARESETn(aic_2_rst_n),
				.ARVALID(ai_core_2_init_lp_I_axi_m_arvalid),
				.ARADDR(ai_core_2_init_lp_I_axi_m_araddr ),
				.ARLEN(ai_core_2_init_lp_I_axi_m_arlen),
				.ARSIZE( ai_core_2_init_lp_I_axi_m_arsize),
				.ARBURST( ai_core_2_init_lp_I_axi_m_arburst ),
				.ARLOCK( ai_core_2_init_lp_I_axi_m_arlock),
				.ARCACHE( ai_core_2_init_lp_I_axi_m_arcache ),
				.ARPROT( ai_core_2_init_lp_I_axi_m_arprot ),
				.ARID( ai_core_2_init_lp_I_axi_m_arid ),
				.ARREADY( ai_core_2_init_lp_I_axi_m_arready ),
				.RREADY( ai_core_2_init_lp_I_axi_m_rready ),
				.RVALID( ai_core_2_init_lp_I_axi_m_rvalid ),
				.RLAST( ai_core_2_init_lp_I_axi_m_rlast ),
				.RDATA(  ai_core_2_init_lp_I_axi_m_rdata ),
				.RRESP( ai_core_2_init_lp_I_axi_m_rresp ),
				.RID( ai_core_2_init_lp_I_axi_m_rid ),
				.AWVALID( ai_core_2_init_lp_I_axi_m_awvalid ),
				.AWADDR( ai_core_2_init_lp_I_axi_m_awaddr ),
				.AWLEN( ai_core_2_init_lp_I_axi_m_awlen),
				.AWSIZE( ai_core_2_init_lp_I_axi_m_awsize ),
				.AWBURST( ai_core_2_init_lp_I_axi_m_awburst ),
				.AWLOCK( ai_core_2_init_lp_I_axi_m_awlock ),
				.AWCACHE( ai_core_2_init_lp_I_axi_m_awcache ),
				.AWPROT( ai_core_2_init_lp_I_axi_m_awprot ),
				.AWID( ai_core_2_init_lp_I_axi_m_awid ),
				.AWREADY( ai_core_2_init_lp_I_axi_m_awready ),
				.WVALID( ai_core_2_init_lp_I_axi_m_wvalid ),
				.WLAST( ai_core_2_init_lp_I_axi_m_wlast ),
				.WDATA(  ai_core_2_init_lp_I_axi_m_wdata ),
				.WSTRB( ai_core_2_init_lp_I_axi_m_wstrb ),
				.WREADY( ai_core_2_init_lp_I_axi_m_wready),
				.BREADY( ai_core_2_init_lp_I_axi_m_bready ),
				.BVALID( ai_core_2_init_lp_I_axi_m_bvalid ),
				.BRESP( ai_core_2_init_lp_I_axi_m_bresp ),
				.BID( ai_core_2_init_lp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//// noc_Targ_lp_ai_core_2

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
			  )
	AXI_Protocol_checker_noc_targ_lp_I_ai_core_2
				(
				.ACLK(aic_2_clk),
				.ARESETn(aic_2_rst_n),
				.ARVALID(ai_core_2_targ_lp_T_axi_s_arvalid),
				.ARADDR(ai_core_2_targ_lp_T_axi_s_araddr ),
				.ARLEN(ai_core_2_targ_lp_T_axi_s_arlen),
				.ARSIZE( ai_core_2_targ_lp_T_axi_s_arsize),
				.ARBURST( ai_core_2_targ_lp_T_axi_s_arburst ),
				.ARLOCK( ai_core_2_targ_lp_T_axi_s_arlock),
				.ARCACHE( ai_core_2_targ_lp_T_axi_s_arcache ),
				.ARPROT( ai_core_2_targ_lp_T_axi_s_arprot ),
				.ARID( ai_core_2_targ_lp_T_axi_s_arid ),
				.ARREADY( ai_core_2_targ_lp_T_axi_s_arready ),
				.RREADY( ai_core_2_targ_lp_T_axi_s_rready ),
				.RVALID( ai_core_2_targ_lp_T_axi_s_rvalid ),
				.RLAST( ai_core_2_targ_lp_T_axi_s_rlast ),
				.RDATA(  ai_core_2_targ_lp_T_axi_s_rdata ),
				.RRESP( ai_core_2_targ_lp_T_axi_s_rresp ),
				.RID( ai_core_2_targ_lp_T_axi_s_rid ),
				.AWVALID( ai_core_2_targ_lp_T_axi_s_awvalid ),
				.AWADDR( ai_core_2_targ_lp_T_axi_s_awaddr ),
				.AWLEN( ai_core_2_targ_lp_T_axi_s_awlen),
				.AWSIZE( ai_core_2_targ_lp_T_axi_s_awsize ),
				.AWBURST( ai_core_2_targ_lp_T_axi_s_awburst ),
				.AWLOCK( ai_core_2_targ_lp_T_axi_s_awlock ),
				.AWCACHE( ai_core_2_targ_lp_T_axi_s_awcache ),
				.AWPROT( ai_core_2_targ_lp_T_axi_s_awprot ),
				.AWID( ai_core_2_targ_lp_T_axi_s_awid ),
				.AWREADY( ai_core_2_targ_lp_T_axi_s_awready ),
				.WVALID( ai_core_2_targ_lp_T_axi_s_wvalid ),
				.WLAST( ai_core_2_targ_lp_T_axi_s_wlast ),
				.WDATA(  ai_core_2_targ_lp_T_axi_s_wdata ),
				.WSTRB( ai_core_2_targ_lp_T_axi_s_wstrb ),
				.WREADY( ai_core_2_targ_lp_T_axi_s_wready),
				.BREADY( ai_core_2_targ_lp_T_axi_s_bready ),
				.BVALID( ai_core_2_targ_lp_T_axi_s_bvalid ),
				.BRESP( ai_core_2_targ_lp_T_axi_s_bresp ),
				.BID( ai_core_2_targ_lp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

//triton_noc_hp_ai_core_3

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (9),
				.WID_WIDTH  (9),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_hp_I_ai_core_3
				(
				.ACLK(aic_3_clk),
				.ARESETn(aic_3_rst_n),
				.ARVALID(ai_core_3_init_hp_I_axi_m_arvalid),
				.ARADDR(ai_core_3_init_hp_I_axi_m_araddr ),
				.ARLEN(ai_core_3_init_hp_I_axi_m_arlen),
				.ARSIZE( ai_core_3_init_hp_I_axi_m_arsize),
				.ARBURST( ai_core_3_init_hp_I_axi_m_arburst ),
				.ARLOCK( ai_core_3_init_hp_I_axi_m_arlock),
				.ARCACHE( ai_core_3_init_hp_I_axi_m_arcache ),
				.ARPROT( ai_core_3_init_hp_I_axi_m_arprot ),
				.ARID( ai_core_3_init_hp_I_axi_m_arid ),
				.ARREADY( ai_core_3_init_hp_I_axi_m_arready ),
				.RREADY( ai_core_3_init_hp_I_axi_m_rready ),
				.RVALID( ai_core_3_init_hp_I_axi_m_rvalid ),
				.RLAST( ai_core_3_init_hp_I_axi_m_rlast ),
				.RDATA(  ai_core_3_init_hp_I_axi_m_rdata ),
				.RRESP( ai_core_3_init_hp_I_axi_m_rresp ),
				.RID( ai_core_3_init_hp_I_axi_m_rid ),
				.AWVALID( ai_core_3_init_hp_I_axi_m_awvalid ),
				.AWADDR( ai_core_3_init_hp_I_axi_m_awaddr ),
				.AWLEN( ai_core_3_init_hp_I_axi_m_awlen),
				.AWSIZE( ai_core_3_init_hp_I_axi_m_awsize ),
				.AWBURST( ai_core_3_init_hp_I_axi_m_awburst ),
				.AWLOCK( ai_core_3_init_hp_I_axi_m_awlock ),
				.AWCACHE( ai_core_3_init_hp_I_axi_m_awcache ),
				.AWPROT( ai_core_3_init_hp_I_axi_m_awprot ),
				.AWID( ai_core_3_init_hp_I_axi_m_awid ),
				.AWREADY( ai_core_3_init_hp_I_axi_m_awready ),
				.WVALID( ai_core_3_init_hp_I_axi_m_wvalid ),
				.WLAST( ai_core_3_init_hp_I_axi_m_wlast ),
				.WDATA(  ai_core_3_init_hp_I_axi_m_wdata ),
				.WSTRB( ai_core_3_init_hp_I_axi_m_wstrb ),
				.WREADY( ai_core_3_init_hp_I_axi_m_wready),
				.BREADY( ai_core_3_init_hp_I_axi_m_bready ),
				.BVALID( ai_core_3_init_hp_I_axi_m_bvalid ),
				.BRESP( ai_core_3_init_hp_I_axi_m_bresp ),
				.BID( ai_core_3_init_hp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

//noc_init_lp_ai_core_3
bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (9),
				.WID_WIDTH  (9),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_lp_I_ai_core_3
				(
				.ACLK(aic_3_clk),
				.ARESETn(aic_3_rst_n),
				.ARVALID(ai_core_3_init_lp_I_axi_m_arvalid),
				.ARADDR(ai_core_3_init_lp_I_axi_m_araddr ),
				.ARLEN(ai_core_3_init_lp_I_axi_m_arlen),
				.ARSIZE( ai_core_3_init_lp_I_axi_m_arsize),
				.ARBURST( ai_core_3_init_lp_I_axi_m_arburst ),
				.ARLOCK( ai_core_3_init_lp_I_axi_m_arlock),
				.ARCACHE( ai_core_3_init_lp_I_axi_m_arcache ),
				.ARPROT( ai_core_3_init_lp_I_axi_m_arprot ),
				.ARID( ai_core_3_init_lp_I_axi_m_arid ),
				.ARREADY( ai_core_3_init_lp_I_axi_m_arready ),
				.RREADY( ai_core_3_init_lp_I_axi_m_rready ),
				.RVALID( ai_core_3_init_lp_I_axi_m_rvalid ),
				.RLAST( ai_core_3_init_lp_I_axi_m_rlast ),
				.RDATA(  ai_core_3_init_lp_I_axi_m_rdata ),
				.RRESP( ai_core_3_init_lp_I_axi_m_rresp ),
				.RID( ai_core_3_init_lp_I_axi_m_rid ),
				.AWVALID( ai_core_3_init_lp_I_axi_m_awvalid ),
				.AWADDR( ai_core_3_init_lp_I_axi_m_awaddr ),
				.AWLEN( ai_core_3_init_lp_I_axi_m_awlen),
				.AWSIZE( ai_core_3_init_lp_I_axi_m_awsize ),
				.AWBURST( ai_core_3_init_lp_I_axi_m_awburst ),
				.AWLOCK( ai_core_3_init_lp_I_axi_m_awlock ),
				.AWCACHE( ai_core_3_init_lp_I_axi_m_awcache ),
				.AWPROT( ai_core_3_init_lp_I_axi_m_awprot ),
				.AWID( ai_core_3_init_lp_I_axi_m_awid ),
				.AWREADY( ai_core_3_init_lp_I_axi_m_awready ),
				.WVALID( ai_core_3_init_lp_I_axi_m_wvalid ),
				.WLAST( ai_core_3_init_lp_I_axi_m_wlast ),
				.WDATA(  ai_core_3_init_lp_I_axi_m_wdata ),
				.WSTRB( ai_core_3_init_lp_I_axi_m_wstrb ),
				.WREADY( ai_core_3_init_lp_I_axi_m_wready),
				.BREADY( ai_core_3_init_lp_I_axi_m_bready ),
				.BVALID( ai_core_3_init_lp_I_axi_m_bvalid ),
				.BRESP( ai_core_3_init_lp_I_axi_m_bresp ),
				.BID( ai_core_3_init_lp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//// noc_Targ_lp_ai_core_3

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_noc_targ_lp_I_ai_core_3
				(
				.ACLK(aic_3_clk),
				.ARESETn(aic_3_rst_n),
				.ARVALID(ai_core_3_targ_lp_T_axi_s_arvalid),
				.ARADDR(ai_core_3_targ_lp_T_axi_s_araddr ),
				.ARLEN(ai_core_3_targ_lp_T_axi_s_arlen),
				.ARSIZE( ai_core_3_targ_lp_T_axi_s_arsize),
				.ARBURST( ai_core_3_targ_lp_T_axi_s_arburst ),
				.ARLOCK( ai_core_3_targ_lp_T_axi_s_arlock),
				.ARCACHE( ai_core_3_targ_lp_T_axi_s_arcache ),
				.ARPROT( ai_core_3_targ_lp_T_axi_s_arprot ),
				.ARID( ai_core_3_targ_lp_T_axi_s_arid ),
				.ARREADY( ai_core_3_targ_lp_T_axi_s_arready ),
				.RREADY( ai_core_3_targ_lp_T_axi_s_rready ),
				.RVALID( ai_core_3_targ_lp_T_axi_s_rvalid ),
				.RLAST( ai_core_3_targ_lp_T_axi_s_rlast ),
				.RDATA(  ai_core_3_targ_lp_T_axi_s_rdata ),
				.RRESP( ai_core_3_targ_lp_T_axi_s_rresp ),
				.RID( ai_core_3_targ_lp_T_axi_s_rid ),
				.AWVALID( ai_core_3_targ_lp_T_axi_s_awvalid ),
				.AWADDR( ai_core_3_targ_lp_T_axi_s_awaddr ),
				.AWLEN( ai_core_3_targ_lp_T_axi_s_awlen),
				.AWSIZE( ai_core_3_targ_lp_T_axi_s_awsize ),
				.AWBURST( ai_core_3_targ_lp_T_axi_s_awburst ),
				.AWLOCK( ai_core_3_targ_lp_T_axi_s_awlock ),
				.AWCACHE( ai_core_3_targ_lp_T_axi_s_awcache ),
				.AWPROT( ai_core_3_targ_lp_T_axi_s_awprot ),
				.AWID( ai_core_3_targ_lp_T_axi_s_awid ),
				.AWREADY( ai_core_3_targ_lp_T_axi_s_awready ),
				.WVALID( ai_core_3_targ_lp_T_axi_s_wvalid ),
				.WLAST( ai_core_3_targ_lp_T_axi_s_wlast ),
				.WDATA(  ai_core_3_targ_lp_T_axi_s_wdata ),
				.WSTRB( ai_core_3_targ_lp_T_axi_s_wstrb ),
				.WREADY( ai_core_3_targ_lp_T_axi_s_wready),
				.BREADY( ai_core_3_targ_lp_T_axi_s_bready ),
				.BVALID( ai_core_3_targ_lp_T_axi_s_bvalid ),
				.BRESP( ai_core_3_targ_lp_T_axi_s_bresp ),
				.BID( ai_core_3_targ_lp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


// triton_noc_l2_hp_0


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (4),
				.WID_WIDTH  (4),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_l2_0_targ_hp_axi_s
				(
				.ACLK(l2_0_clk),
				.ARESETn(l2_0_rst_n),
				.ARVALID(l2_0_targ_hp_T_axi_s_arvalid),
				.ARADDR(l2_0_targ_hp_T_axi_s_araddr ),
				.ARLEN(l2_0_targ_hp_T_axi_s_arlen),
				.ARSIZE( l2_0_targ_hp_T_axi_s_arsize),
				.ARBURST( l2_0_targ_hp_T_axi_s_arburst ),
				.ARLOCK( l2_0_targ_hp_T_axi_s_arlock),
				.ARCACHE( l2_0_targ_hp_T_axi_s_arcache ),
				.ARPROT( l2_0_targ_hp_T_axi_s_arprot ),
				.ARID( l2_0_targ_hp_T_axi_s_arid ),
				.ARREADY( l2_0_targ_hp_T_axi_s_arready ),
				.RREADY( l2_0_targ_hp_T_axi_s_rready ),
				.RVALID( l2_0_targ_hp_T_axi_s_rvalid ),
				.RLAST( l2_0_targ_hp_T_axi_s_rlast ),
				.RDATA(  l2_0_targ_hp_T_axi_s_rdata ),
				.RRESP( l2_0_targ_hp_T_axi_s_rresp ),
				.RID( l2_0_targ_hp_T_axi_s_rid ),
				.AWVALID( l2_0_targ_hp_T_axi_s_awvalid ),
				.AWADDR( l2_0_targ_hp_T_axi_s_awaddr ),
				.AWLEN( l2_0_targ_hp_T_axi_s_awlen),
				.AWSIZE( l2_0_targ_hp_T_axi_s_awsize ),
				.AWBURST( l2_0_targ_hp_T_axi_s_awburst ),
				.AWLOCK( l2_0_targ_hp_T_axi_s_awlock ),
				.AWCACHE( l2_0_targ_hp_T_axi_s_awcache ),
				.AWPROT( l2_0_targ_hp_T_axi_s_awprot ),
				.AWID( l2_0_targ_hp_T_axi_s_awid ),
				.AWREADY( l2_0_targ_hp_T_axi_s_awready ),
				.WVALID( l2_0_targ_hp_T_axi_s_wvalid ),
				.WLAST( l2_0_targ_hp_T_axi_s_wlast ),
				.WDATA(  l2_0_targ_hp_T_axi_s_wdata ),
				.WSTRB( l2_0_targ_hp_T_axi_s_wstrb ),
				.WREADY( l2_0_targ_hp_T_axi_s_wready),
				.BREADY( l2_0_targ_hp_T_axi_s_bready ),
				.BVALID( l2_0_targ_hp_T_axi_s_bvalid ),
				.BRESP( l2_0_targ_hp_T_axi_s_bresp ),
				.BID( l2_0_targ_hp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

// l2_1_targ_hp


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (4),
				.WID_WIDTH  (4),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_l2_1_targ_hp_axi_s
				(
				.ACLK(l2_1_clk),
				.ARESETn(l2_1_rst_n),
				.ARVALID(l2_1_targ_hp_T_axi_s_arvalid),
				.ARADDR(l2_1_targ_hp_T_axi_s_araddr ),
				.ARLEN(l2_1_targ_hp_T_axi_s_arlen),
				.ARSIZE( l2_1_targ_hp_T_axi_s_arsize),
				.ARBURST( l2_1_targ_hp_T_axi_s_arburst ),
				.ARLOCK( l2_1_targ_hp_T_axi_s_arlock),
				.ARCACHE( l2_1_targ_hp_T_axi_s_arcache ),
				.ARPROT( l2_1_targ_hp_T_axi_s_arprot ),
				.ARID( l2_1_targ_hp_T_axi_s_arid ),
				.ARREADY( l2_1_targ_hp_T_axi_s_arready ),
				.RREADY( l2_1_targ_hp_T_axi_s_rready ),
				.RVALID( l2_1_targ_hp_T_axi_s_rvalid ),
				.RLAST( l2_1_targ_hp_T_axi_s_rlast ),
				.RDATA(  l2_1_targ_hp_T_axi_s_rdata ),
				.RRESP( l2_1_targ_hp_T_axi_s_rresp ),
				.RID( l2_1_targ_hp_T_axi_s_rid ),
				.AWVALID( l2_1_targ_hp_T_axi_s_awvalid ),
				.AWADDR( l2_1_targ_hp_T_axi_s_awaddr ),
				.AWLEN( l2_1_targ_hp_T_axi_s_awlen),
				.AWSIZE( l2_1_targ_hp_T_axi_s_awsize ),
				.AWBURST( l2_1_targ_hp_T_axi_s_awburst ),
				.AWLOCK( l2_1_targ_hp_T_axi_s_awlock ),
				.AWCACHE( l2_1_targ_hp_T_axi_s_awcache ),
				.AWPROT( l2_1_targ_hp_T_axi_s_awprot ),
				.AWID( l2_1_targ_hp_T_axi_s_awid ),
				.AWREADY( l2_1_targ_hp_T_axi_s_awready ),
				.WVALID( l2_1_targ_hp_T_axi_s_wvalid ),
				.WLAST( l2_1_targ_hp_T_axi_s_wlast ),
				.WDATA(  l2_1_targ_hp_T_axi_s_wdata ),
				.WSTRB( l2_1_targ_hp_T_axi_s_wstrb ),
				.WREADY( l2_1_targ_hp_T_axi_s_wready),
				.BREADY( l2_1_targ_hp_T_axi_s_bready ),
				.BVALID( l2_1_targ_hp_T_axi_s_bvalid ),
				.BRESP( l2_1_targ_hp_T_axi_s_bresp ),
				.BID( l2_1_targ_hp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//l2_2_targ_hp_T


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (4),
				.WID_WIDTH  (4),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_l2_2_targ_hp_axi_s
				(
				.ACLK(l2_2_clk),
				.ARESETn(l2_2_rst_n),
				.ARVALID(l2_2_targ_hp_T_axi_s_arvalid),
				.ARADDR(l2_2_targ_hp_T_axi_s_araddr ),
				.ARLEN(l2_2_targ_hp_T_axi_s_arlen),
				.ARSIZE( l2_2_targ_hp_T_axi_s_arsize),
				.ARBURST( l2_2_targ_hp_T_axi_s_arburst ),
				.ARLOCK( l2_2_targ_hp_T_axi_s_arlock),
				.ARCACHE( l2_2_targ_hp_T_axi_s_arcache ),
				.ARPROT( l2_2_targ_hp_T_axi_s_arprot ),
				.ARID( l2_2_targ_hp_T_axi_s_arid ),
				.ARREADY( l2_2_targ_hp_T_axi_s_arready ),
				.RREADY( l2_2_targ_hp_T_axi_s_rready ),
				.RVALID( l2_2_targ_hp_T_axi_s_rvalid ),
				.RLAST( l2_2_targ_hp_T_axi_s_rlast ),
				.RDATA(  l2_2_targ_hp_T_axi_s_rdata ),
				.RRESP( l2_2_targ_hp_T_axi_s_rresp ),
				.RID( l2_2_targ_hp_T_axi_s_rid ),
				.AWVALID( l2_2_targ_hp_T_axi_s_awvalid ),
				.AWADDR( l2_2_targ_hp_T_axi_s_awaddr ),
				.AWLEN( l2_2_targ_hp_T_axi_s_awlen),
				.AWSIZE( l2_2_targ_hp_T_axi_s_awsize ),
				.AWBURST( l2_2_targ_hp_T_axi_s_awburst ),
				.AWLOCK( l2_2_targ_hp_T_axi_s_awlock ),
				.AWCACHE( l2_2_targ_hp_T_axi_s_awcache ),
				.AWPROT( l2_2_targ_hp_T_axi_s_awprot ),
				.AWID( l2_2_targ_hp_T_axi_s_awid ),
				.AWREADY( l2_2_targ_hp_T_axi_s_awready ),
				.WVALID( l2_2_targ_hp_T_axi_s_wvalid ),
				.WLAST( l2_2_targ_hp_T_axi_s_wlast ),
				.WDATA(  l2_2_targ_hp_T_axi_s_wdata ),
				.WSTRB( l2_2_targ_hp_T_axi_s_wstrb ),
				.WREADY( l2_2_targ_hp_T_axi_s_wready),
				.BREADY( l2_2_targ_hp_T_axi_s_bready ),
				.BVALID( l2_2_targ_hp_T_axi_s_bvalid ),
				.BRESP( l2_2_targ_hp_T_axi_s_bresp ),
				.BID( l2_2_targ_hp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


// l2_3_targ_hp_T


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (4),
				.WID_WIDTH  (4),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_l2_3_targ_hp_axi_s
				(
				.ACLK(l2_3_clk),
				.ARESETn(l2_3_rst_n),
				.ARVALID(l2_3_targ_hp_T_axi_s_arvalid),
				.ARADDR(l2_3_targ_hp_T_axi_s_araddr ),
				.ARLEN(l2_3_targ_hp_T_axi_s_arlen),
				.ARSIZE( l2_3_targ_hp_T_axi_s_arsize),
				.ARBURST( l2_3_targ_hp_T_axi_s_arburst ),
				.ARLOCK( l2_3_targ_hp_T_axi_s_arlock),
				.ARCACHE( l2_3_targ_hp_T_axi_s_arcache ),
				.ARPROT( l2_3_targ_hp_T_axi_s_arprot ),
				.ARID( l2_3_targ_hp_T_axi_s_arid ),
				.ARREADY( l2_3_targ_hp_T_axi_s_arready ),
				.RREADY( l2_3_targ_hp_T_axi_s_rready ),
				.RVALID( l2_3_targ_hp_T_axi_s_rvalid ),
				.RLAST( l2_3_targ_hp_T_axi_s_rlast ),
				.RDATA(  l2_3_targ_hp_T_axi_s_rdata ),
				.RRESP( l2_3_targ_hp_T_axi_s_rresp ),
				.RID( l2_3_targ_hp_T_axi_s_rid ),
				.AWVALID( l2_3_targ_hp_T_axi_s_awvalid ),
				.AWADDR( l2_3_targ_hp_T_axi_s_awaddr ),
				.AWLEN( l2_3_targ_hp_T_axi_s_awlen),
				.AWSIZE( l2_3_targ_hp_T_axi_s_awsize ),
				.AWBURST( l2_3_targ_hp_T_axi_s_awburst ),
				.AWLOCK( l2_3_targ_hp_T_axi_s_awlock ),
				.AWCACHE( l2_3_targ_hp_T_axi_s_awcache ),
				.AWPROT( l2_3_targ_hp_T_axi_s_awprot ),
				.AWID( l2_3_targ_hp_T_axi_s_awid ),
				.AWREADY( l2_3_targ_hp_T_axi_s_awready ),
				.WVALID( l2_3_targ_hp_T_axi_s_wvalid ),
				.WLAST( l2_3_targ_hp_T_axi_s_wlast ),
				.WDATA(  l2_3_targ_hp_T_axi_s_wdata ),
				.WSTRB( l2_3_targ_hp_T_axi_s_wstrb ),
				.WREADY( l2_3_targ_hp_T_axi_s_wready),
				.BREADY( l2_3_targ_hp_T_axi_s_bready ),
				.BVALID( l2_3_targ_hp_T_axi_s_bvalid ),
				.BRESP( l2_3_targ_hp_T_axi_s_bresp ),
				.BID( l2_3_targ_hp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//sys_ctrl_init_lp_I_axi


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_sys_ctrl_init_lp_axi_m
				(
				.ACLK(sys_ctrl_clk),
				.ARESETn(sys_ctrl_rst_n),
				.ARVALID(sys_ctrl_init_lp_I_axi_m_arvalid),
				.ARADDR(sys_ctrl_init_lp_I_axi_m_araddr ),
				.ARLEN(sys_ctrl_init_lp_I_axi_m_arlen),
				.ARSIZE( sys_ctrl_init_lp_I_axi_m_arsize),
				.ARBURST( sys_ctrl_init_lp_I_axi_m_arburst ),
				.ARLOCK( sys_ctrl_init_lp_I_axi_m_arlock),
				.ARCACHE( sys_ctrl_init_lp_I_axi_m_arcache ),
				.ARPROT( sys_ctrl_init_lp_I_axi_m_arprot ),
				.ARID( sys_ctrl_init_lp_I_axi_m_arid ),
				.ARREADY( sys_ctrl_init_lp_I_axi_m_arready ),
				.RREADY( sys_ctrl_init_lp_I_axi_m_rready ),
				.RVALID( sys_ctrl_init_lp_I_axi_m_rvalid ),
				.RLAST( sys_ctrl_init_lp_I_axi_m_rlast ),
				.RDATA(  sys_ctrl_init_lp_I_axi_m_rdata ),
				.RRESP( sys_ctrl_init_lp_I_axi_m_rresp ),
				.RID( sys_ctrl_init_lp_I_axi_m_rid ),
				.AWVALID( sys_ctrl_init_lp_I_axi_m_awvalid ),
				.AWADDR( sys_ctrl_init_lp_I_axi_m_awaddr ),
				.AWLEN( sys_ctrl_init_lp_I_axi_m_awlen),
				.AWSIZE( sys_ctrl_init_lp_I_axi_m_awsize ),
				.AWBURST( sys_ctrl_init_lp_I_axi_m_awburst ),
				.AWLOCK( sys_ctrl_init_lp_I_axi_m_awlock ),
				.AWCACHE( sys_ctrl_init_lp_I_axi_m_awcache ),
				.AWPROT( sys_ctrl_init_lp_I_axi_m_awprot ),
				.AWID( sys_ctrl_init_lp_I_axi_m_awid ),
				.AWREADY( sys_ctrl_init_lp_I_axi_m_awready ),
				.WVALID( sys_ctrl_init_lp_I_axi_m_wvalid ),
				.WLAST( sys_ctrl_init_lp_I_axi_m_wlast ),
				.WDATA(  sys_ctrl_init_lp_I_axi_m_wdata ),
				.WSTRB( sys_ctrl_init_lp_I_axi_m_wstrb ),
				.WREADY( sys_ctrl_init_lp_I_axi_m_wready),
				.BREADY( sys_ctrl_init_lp_I_axi_m_bready ),
				.BVALID( sys_ctrl_init_lp_I_axi_m_bvalid ),
				.BRESP( sys_ctrl_init_lp_I_axi_m_bresp ),
				.BID( sys_ctrl_init_lp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//sys_ctrl_targ_lp_T

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (4),
				.WID_WIDTH  (4),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_sys_ctrl_targ_lp_axi_s
				(
				.ACLK(sys_ctrl_clk),
				.ARESETn(sys_ctrl_rst_n),
				.ARVALID(sys_ctrl_targ_lp_T_axi_s_arvalid),
				.ARADDR(sys_ctrl_targ_lp_T_axi_s_araddr ),
				.ARLEN(sys_ctrl_targ_lp_T_axi_s_arlen),
				.ARSIZE( sys_ctrl_targ_lp_T_axi_s_arsize),
				.ARBURST( sys_ctrl_targ_lp_T_axi_s_arburst ),
				.ARLOCK( sys_ctrl_targ_lp_T_axi_s_arlock),
				.ARCACHE( sys_ctrl_targ_lp_T_axi_s_arcache ),
				.ARPROT( sys_ctrl_targ_lp_T_axi_s_arprot ),
				.ARID( sys_ctrl_targ_lp_T_axi_s_arid ),
				.ARREADY( sys_ctrl_targ_lp_T_axi_s_arready ),
				.RREADY( sys_ctrl_targ_lp_T_axi_s_rready ),
				.RVALID( sys_ctrl_targ_lp_T_axi_s_rvalid ),
				.RLAST( sys_ctrl_targ_lp_T_axi_s_rlast ),
				.RDATA(  sys_ctrl_targ_lp_T_axi_s_rdata ),
				.RRESP( sys_ctrl_targ_lp_T_axi_s_rresp ),
				.RID( sys_ctrl_targ_lp_T_axi_s_rid ),
				.AWVALID( sys_ctrl_targ_lp_T_axi_s_awvalid ),
				.AWADDR( sys_ctrl_targ_lp_T_axi_s_awaddr ),
				.AWLEN( sys_ctrl_targ_lp_T_axi_s_awlen),
				.AWSIZE( sys_ctrl_targ_lp_T_axi_s_awsize ),
				.AWBURST( sys_ctrl_targ_lp_T_axi_s_awburst ),
				.AWLOCK( sys_ctrl_targ_lp_T_axi_s_awlock ),
				.AWCACHE( sys_ctrl_targ_lp_T_axi_s_awcache ),
				.AWPROT( sys_ctrl_targ_lp_T_axi_s_awprot ),
				.AWID( sys_ctrl_targ_lp_T_axi_s_awid ),
				.AWREADY( sys_ctrl_targ_lp_T_axi_s_awready ),
				.WVALID( sys_ctrl_targ_lp_T_axi_s_wvalid ),
				.WLAST( sys_ctrl_targ_lp_T_axi_s_wlast ),
				.WDATA(  sys_ctrl_targ_lp_T_axi_s_wdata ),
				.WSTRB( sys_ctrl_targ_lp_T_axi_s_wstrb ),
				.WREADY( sys_ctrl_targ_lp_T_axi_s_wready),
				.BREADY( sys_ctrl_targ_lp_T_axi_s_bready ),
				.BVALID( sys_ctrl_targ_lp_T_axi_s_bvalid ),
				.BRESP( sys_ctrl_targ_lp_T_axi_s_bresp ),
				.BID( sys_ctrl_targ_lp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);



//sys_dma_0_init_hp


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_sys_dma_0_init_hp_axi_m
				(
				.ACLK(sys_dma_clk),
				.ARESETn(sys_dma_rst_n),
				.ARVALID(sys_dma_0_init_hp_I_axi_m_arvalid),
				.ARADDR(sys_dma_0_init_hp_I_axi_m_araddr ),
				.ARLEN(sys_dma_0_init_hp_I_axi_m_arlen),
				.ARSIZE( sys_dma_0_init_hp_I_axi_m_arsize),
				.ARBURST( sys_dma_0_init_hp_I_axi_m_arburst ),
				.ARLOCK( sys_dma_0_init_hp_I_axi_m_arlock),
				.ARCACHE( sys_dma_0_init_hp_I_axi_m_arcache ),
				.ARPROT( sys_dma_0_init_hp_I_axi_m_arprot ),
				.ARID( sys_dma_0_init_hp_I_axi_m_arid ),
				.ARREADY( sys_dma_0_init_hp_I_axi_m_arready ),
				.RREADY( sys_dma_0_init_hp_I_axi_m_rready ),
				.RVALID( sys_dma_0_init_hp_I_axi_m_rvalid ),
				.RLAST( sys_dma_0_init_hp_I_axi_m_rlast ),
				.RDATA(  sys_dma_0_init_hp_I_axi_m_rdata ),
				.RRESP( sys_dma_0_init_hp_I_axi_m_rresp ),
				.RID( sys_dma_0_init_hp_I_axi_m_rid ),
				.AWVALID( sys_dma_0_init_hp_I_axi_m_awvalid ),
				.AWADDR( sys_dma_0_init_hp_I_axi_m_awaddr ),
				.AWLEN( sys_dma_0_init_hp_I_axi_m_awlen),
				.AWSIZE( sys_dma_0_init_hp_I_axi_m_awsize ),
				.AWBURST( sys_dma_0_init_hp_I_axi_m_awburst ),
				.AWLOCK( sys_dma_0_init_hp_I_axi_m_awlock ),
				.AWCACHE( sys_dma_0_init_hp_I_axi_m_awcache ),
				.AWPROT( sys_dma_0_init_hp_I_axi_m_awprot ),
				.AWID( sys_dma_0_init_hp_I_axi_m_awid ),
				.AWREADY( sys_dma_0_init_hp_I_axi_m_awready ),
				.WVALID( sys_dma_0_init_hp_I_axi_m_wvalid ),
				.WLAST( sys_dma_0_init_hp_I_axi_m_wlast ),
				.WDATA(  sys_dma_0_init_hp_I_axi_m_wdata ),
				.WSTRB( sys_dma_0_init_hp_I_axi_m_wstrb ),
				.WREADY( sys_dma_0_init_hp_I_axi_m_wready),
				.BREADY( sys_dma_0_init_hp_I_axi_m_bready ),
				.BVALID( sys_dma_0_init_hp_I_axi_m_bvalid ),
				.BRESP( sys_dma_0_init_hp_I_axi_m_bresp ),
				.BID( sys_dma_0_init_hp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//sys_dma_1_hp_axi_m

bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_sys_dma_1_init_hp_axi_m
				(
				.ACLK(sys_dma_clk),
				.ARESETn(sys_dma_rst_n),
				.ARVALID(sys_dma_1_init_hp_I_axi_m_arvalid),
				.ARADDR(sys_dma_1_init_hp_I_axi_m_araddr ),
				.ARLEN(sys_dma_1_init_hp_I_axi_m_arlen),
				.ARSIZE( sys_dma_1_init_hp_I_axi_m_arsize),
				.ARBURST( sys_dma_1_init_hp_I_axi_m_arburst ),
				.ARLOCK( sys_dma_1_init_hp_I_axi_m_arlock),
				.ARCACHE( sys_dma_1_init_hp_I_axi_m_arcache ),
				.ARPROT( sys_dma_1_init_hp_I_axi_m_arprot ),
				.ARID( sys_dma_1_init_hp_I_axi_m_arid ),
				.ARREADY( sys_dma_1_init_hp_I_axi_m_arready ),
				.RREADY( sys_dma_1_init_hp_I_axi_m_rready ),
				.RVALID( sys_dma_1_init_hp_I_axi_m_rvalid ),
				.RLAST( sys_dma_1_init_hp_I_axi_m_rlast ),
				.RDATA(  sys_dma_1_init_hp_I_axi_m_rdata ),
				.RRESP( sys_dma_1_init_hp_I_axi_m_rresp ),
				.RID( sys_dma_1_init_hp_I_axi_m_rid ),
				.AWVALID( sys_dma_1_init_hp_I_axi_m_awvalid ),
				.AWADDR( sys_dma_1_init_hp_I_axi_m_awaddr ),
				.AWLEN( sys_dma_1_init_hp_I_axi_m_awlen),
				.AWSIZE( sys_dma_1_init_hp_I_axi_m_awsize ),
				.AWBURST( sys_dma_1_init_hp_I_axi_m_awburst ),
				.AWLOCK( sys_dma_1_init_hp_I_axi_m_awlock ),
				.AWCACHE( sys_dma_1_init_hp_I_axi_m_awcache ),
				.AWPROT( sys_dma_1_init_hp_I_axi_m_awprot ),
				.AWID( sys_dma_1_init_hp_I_axi_m_awid ),
				.AWREADY( sys_dma_1_init_hp_I_axi_m_awready ),
				.WVALID( sys_dma_1_init_hp_I_axi_m_wvalid ),
				.WLAST( sys_dma_1_init_hp_I_axi_m_wlast ),
				.WDATA(  sys_dma_1_init_hp_I_axi_m_wdata ),
				.WSTRB( sys_dma_1_init_hp_I_axi_m_wstrb ),
				.WREADY( sys_dma_1_init_hp_I_axi_m_wready),
				.BREADY( sys_dma_1_init_hp_I_axi_m_bready ),
				.BVALID( sys_dma_1_init_hp_I_axi_m_bvalid ),
				.BRESP( sys_dma_1_init_hp_I_axi_m_bresp ),
				.BID( sys_dma_1_init_hp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

//pcie_init_hp_I_axi_m


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_pcie_init_hp_I_axi_m
				(
				.ACLK(pcie_mst_clk),
				.ARESETn(pcie_mst_rst_n),
				.ARVALID(pcie_init_hp_I_axi_m_arvalid),
				.ARADDR(pcie_init_hp_I_axi_m_araddr ),
				.ARLEN(pcie_init_hp_I_axi_m_arlen),
				.ARSIZE( pcie_init_hp_I_axi_m_arsize),
				.ARBURST( pcie_init_hp_I_axi_m_arburst ),
				.ARLOCK( pcie_init_hp_I_axi_m_arlock),
				.ARCACHE( pcie_init_hp_I_axi_m_arcache ),
				.ARPROT( pcie_init_hp_I_axi_m_arprot ),
				.ARID( pcie_init_hp_I_axi_m_arid ),
				.ARREADY( pcie_init_hp_I_axi_m_arready ),
				.RREADY( pcie_init_hp_I_axi_m_rready ),
				.RVALID( pcie_init_hp_I_axi_m_rvalid ),
				.RLAST( pcie_init_hp_I_axi_m_rlast ),
				.RDATA(  pcie_init_hp_I_axi_m_rdata ),
				.RRESP( pcie_init_hp_I_axi_m_rresp ),
				.RID( pcie_init_hp_I_axi_m_rid ),
				.AWVALID( pcie_init_hp_I_axi_m_awvalid ),
				.AWADDR( pcie_init_hp_I_axi_m_awaddr ),
				.AWLEN( pcie_init_hp_I_axi_m_awlen),
				.AWSIZE( pcie_init_hp_I_axi_m_awsize ),
				.AWBURST( pcie_init_hp_I_axi_m_awburst ),
				.AWLOCK( pcie_init_hp_I_axi_m_awlock ),
				.AWCACHE( pcie_init_hp_I_axi_m_awcache ),
				.AWPROT( pcie_init_hp_I_axi_m_awprot ),
				.AWID( pcie_init_hp_I_axi_m_awid ),
				.AWREADY( pcie_init_hp_I_axi_m_awready ),
				.WVALID( pcie_init_hp_I_axi_m_wvalid ),
				.WLAST( pcie_init_hp_I_axi_m_wlast ),
				.WDATA(  pcie_init_hp_I_axi_m_wdata ),
				.WSTRB( pcie_init_hp_I_axi_m_wstrb ),
				.WREADY( pcie_init_hp_I_axi_m_wready),
				.BREADY( pcie_init_hp_I_axi_m_bready ),
				.BVALID( pcie_init_hp_I_axi_m_bvalid ),
				.BRESP( pcie_init_hp_I_axi_m_bresp ),
				.BID( pcie_init_hp_I_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);



//pcie_targ_dbi_T_axi_s


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(32),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (4),
				.WID_WIDTH  (4),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_pcie_targ_dbi_T_axi_s
				(
				.ACLK(pcie_dbi_clk),
				.ARESETn(pcie_dbi_rst_n),
				.ARVALID(pcie_targ_dbi_T_axi_s_arvalid),
				.ARADDR(pcie_targ_dbi_T_axi_s_araddr ),
				.ARLEN(pcie_targ_dbi_T_axi_s_arlen),
				.ARSIZE( pcie_targ_dbi_T_axi_s_arsize),
				.ARBURST( pcie_targ_dbi_T_axi_s_arburst ),
				.ARLOCK( pcie_targ_dbi_T_axi_s_arlock),
				.ARCACHE( pcie_targ_dbi_T_axi_s_arcache ),
				.ARPROT( pcie_targ_dbi_T_axi_s_arprot ),
				.ARID( pcie_targ_dbi_T_axi_s_arid ),
				.ARREADY( pcie_targ_dbi_T_axi_s_arready ),
				.RREADY( pcie_targ_dbi_T_axi_s_rready ),
				.RVALID( pcie_targ_dbi_T_axi_s_rvalid ),
				.RLAST( pcie_targ_dbi_T_axi_s_rlast ),
				.RDATA(  pcie_targ_dbi_T_axi_s_rdata ),
				.RRESP( pcie_targ_dbi_T_axi_s_rresp ),
				.RID( pcie_targ_dbi_T_axi_s_rid ),
				.AWVALID( pcie_targ_dbi_T_axi_s_awvalid ),
				.AWADDR( pcie_targ_dbi_T_axi_s_awaddr ),
				.AWLEN( pcie_targ_dbi_T_axi_s_awlen),
				.AWSIZE( pcie_targ_dbi_T_axi_s_awsize ),
				.AWBURST( pcie_targ_dbi_T_axi_s_awburst ),
				.AWLOCK( pcie_targ_dbi_T_axi_s_awlock ),
				.AWCACHE( pcie_targ_dbi_T_axi_s_awcache ),
				.AWPROT( pcie_targ_dbi_T_axi_s_awprot ),
				.AWID( pcie_targ_dbi_T_axi_s_awid ),
				.AWREADY( pcie_targ_dbi_T_axi_s_awready ),
				.WVALID( pcie_targ_dbi_T_axi_s_wvalid ),
				.WLAST( pcie_targ_dbi_T_axi_s_wlast ),
				.WDATA(  pcie_targ_dbi_T_axi_s_wdata ),
				.WSTRB( pcie_targ_dbi_T_axi_s_wstrb ),
				.WREADY( pcie_targ_dbi_T_axi_s_wready),
				.BREADY( pcie_targ_dbi_T_axi_s_bready ),
				.BVALID( pcie_targ_dbi_T_axi_s_bvalid ),
				.BRESP( pcie_targ_dbi_T_axi_s_bresp ),
				.BID( pcie_targ_dbi_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);



//pcie_targ_lp_I_axi_s


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(64),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (6),
				.WID_WIDTH  (6),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_pcie_targ_lp_T_axi_s
				(
				.ACLK(pcie_slv_clk),
				.ARESETn(pcie_slv_rst_n),
				.ARVALID(pcie_targ_lp_T_axi_s_arvalid),
				.ARADDR(pcie_targ_lp_T_axi_s_araddr ),
				.ARLEN(pcie_targ_lp_T_axi_s_arlen),
				.ARSIZE( pcie_targ_lp_T_axi_s_arsize),
				.ARBURST( pcie_targ_lp_T_axi_s_arburst ),
				.ARLOCK( pcie_targ_lp_T_axi_s_arlock),
				.ARCACHE( pcie_targ_lp_T_axi_s_arcache ),
				.ARPROT( pcie_targ_lp_T_axi_s_arprot ),
				.ARID( pcie_targ_lp_T_axi_s_arid ),
				.ARREADY( pcie_targ_lp_T_axi_s_arready ),
				.RREADY( pcie_targ_lp_T_axi_s_rready ),
				.RVALID( pcie_targ_lp_T_axi_s_rvalid ),
				.RLAST( pcie_targ_lp_T_axi_s_rlast ),
				.RDATA(  pcie_targ_lp_T_axi_s_rdata ),
				.RRESP( pcie_targ_lp_T_axi_s_rresp ),
				.RID( pcie_targ_lp_T_axi_s_rid ),
				.AWVALID( pcie_targ_lp_T_axi_s_awvalid ),
				.AWADDR( pcie_targ_lp_T_axi_s_awaddr ),
				.AWLEN( pcie_targ_lp_T_axi_s_awlen),
				.AWSIZE( pcie_targ_lp_T_axi_s_awsize ),
				.AWBURST( pcie_targ_lp_T_axi_s_awburst ),
				.AWLOCK( pcie_targ_lp_T_axi_s_awlock ),
				.AWCACHE( pcie_targ_lp_T_axi_s_awcache ),
				.AWPROT( pcie_targ_lp_T_axi_s_awprot ),
				.AWID( pcie_targ_lp_T_axi_s_awid ),
				.AWREADY( pcie_targ_lp_T_axi_s_awready ),
				.WVALID( pcie_targ_lp_T_axi_s_wvalid ),
				.WLAST( pcie_targ_lp_T_axi_s_wlast ),
				.WDATA(  pcie_targ_lp_T_axi_s_wdata ),
				.WSTRB( pcie_targ_lp_T_axi_s_wstrb ),
				.WREADY( pcie_targ_lp_T_axi_s_wready),
				.BREADY( pcie_targ_lp_T_axi_s_bready ),
				.BVALID( pcie_targ_lp_T_axi_s_bvalid ),
				.BRESP( pcie_targ_lp_T_axi_s_bresp ),
				.BID( pcie_targ_lp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


//ddrc_targ_mp_T_axi_s


bind triton_noc_p Axi4PC # (
				.DATA_WIDTH(512),
                .ADDR_WIDTH(36),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (8),
				.WID_WIDTH  (8),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
				.AWREADY_MAXWAITS ( 256 ),
        .ARREADY_MAXWAITS ( 256 ),
        .WREADY_MAXWAITS ( 256 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_Protocol_checker_ddrc_targ_mp_T_axi_s
				(
				.ACLK(ddr_axi_clk),
				.ARESETn(ddr_axi_rst_n),
				.ARVALID(ddrc_targ_mp_T_axi_s_arvalid),
				.ARADDR(ddrc_targ_mp_T_axi_s_araddr ),
				.ARLEN(ddrc_targ_mp_T_axi_s_arlen),
				.ARSIZE( ddrc_targ_mp_T_axi_s_arsize),
				.ARBURST( ddrc_targ_mp_T_axi_s_arburst ),
				.ARLOCK( ddrc_targ_mp_T_axi_s_arlock),
				.ARCACHE( ddrc_targ_mp_T_axi_s_arcache ),
				.ARPROT( ddrc_targ_mp_T_axi_s_arprot ),
				.ARID( ddrc_targ_mp_T_axi_s_arid ),
				.ARREADY( ddrc_targ_mp_T_axi_s_arready ),
				.RREADY( ddrc_targ_mp_T_axi_s_rready ),
				.RVALID( ddrc_targ_mp_T_axi_s_rvalid ),
				.RLAST( ddrc_targ_mp_T_axi_s_rlast ),
				.RDATA(  ddrc_targ_mp_T_axi_s_rdata ),
				.RRESP( ddrc_targ_mp_T_axi_s_rresp ),
				.RID( ddrc_targ_mp_T_axi_s_rid ),
				.AWVALID( ddrc_targ_mp_T_axi_s_awvalid ),
				.AWADDR( ddrc_targ_mp_T_axi_s_awaddr ),
				.AWLEN( ddrc_targ_mp_T_axi_s_awlen),
				.AWSIZE( ddrc_targ_mp_T_axi_s_awsize ),
				.AWBURST( ddrc_targ_mp_T_axi_s_awburst ),
				.AWLOCK( ddrc_targ_mp_T_axi_s_awlock ),
				.AWCACHE( ddrc_targ_mp_T_axi_s_awcache ),
				.AWPROT( ddrc_targ_mp_T_axi_s_awprot ),
				.AWID( ddrc_targ_mp_T_axi_s_awid ),
				.AWREADY( ddrc_targ_mp_T_axi_s_awready ),
				.WVALID( ddrc_targ_mp_T_axi_s_wvalid ),
				.WLAST( ddrc_targ_mp_T_axi_s_wlast ),
				.WDATA(  ddrc_targ_mp_T_axi_s_wdata ),
				.WSTRB( ddrc_targ_mp_T_axi_s_wstrb ),
				.WREADY( ddrc_targ_mp_T_axi_s_wready),
				.BREADY( ddrc_targ_mp_T_axi_s_bready ),
				.BVALID( ddrc_targ_mp_T_axi_s_bvalid ),
				.BRESP( ddrc_targ_mp_T_axi_s_bresp ),
				.BID( ddrc_targ_mp_T_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);
