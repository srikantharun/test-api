// (C) Copyright Axelera AI 2022
// All Rights Reserved
// *** Axelera AI Confidential ***

// Description: eFUSE wrapper.

// Module declaration

module soc_mgmt_bus_fabric_wrapper (
   // Ports for Interface ACLK
   input  wire          i_aclk                                    ,
   // Ports for Interface ARESETn,
   input  wire          i_aresetn                                 ,
   // Ports for Interface PCLK,
   input  wire          i_pclk                                    ,
   // Ports for Interface PRESETn,
   input  wire          i_presetn                                 ,
   // Ports for Interface ext_axi_x2h_HCLK,
   input  wire          i_hclk                                    ,
   // Ports for Interface ext_axi_x2h_HRESETn,
   input  wire          i_hresetn                                 ,
    // port for MBIST APB if
   input  logic [31:0]  i_mbist_prdata                            ,
   input  logic         i_apb_mbist_pready                        ,
   input  logic         i_apb_mbist_pslverr                       ,
   output logic [31:0]  o_mbist_paddr                             ,
   output logic         o_mbist_penable                           ,
   output logic         o_mbist_psel                              ,
   output logic [31:0]  o_mbist_pwdata                            ,
   output logic         o_mbist_pwrite                            ,
   // Ports for Interface ex_axi_x2p_s_tms_csr,
   input  logic [31:0]  i_apb_tms_prdata                          ,
   input  logic         i_apb_tms_pready                          ,
   input  logic         i_apb_tms_pslverr                         ,
   output logic [31:0]  o_apb_tms_csr_paddr                       ,
   output logic         o_apb_tms_csr_penable                     ,
   output logic         o_apb_tms_csr_psel                        ,
   output logic [31:0]  o_apb_tms_csr_pwdata                      ,
   output logic         o_apb_tms_csr_pwrite                      ,
   // OTP and ROT AO APB Interface
   input  logic [31:0]  i_apb_rot_ao_and_otp_prdata               ,
   input  logic         i_apb_rot_ao_and_otp_pready               ,
   input  logic         i_apb_rot_ao_and_otp_pslverr              ,
   output logic [31:0]  o_apb_rot_ao_and_otp_paddr                ,
   output logic         o_apb_rot_ao_and_otp_penable              ,
   output logic         o_apb_rot_ao_and_otp_psel                 ,
   output logic [31:0]  o_apb_rot_ao_and_otp_pwdata               ,
   output logic         o_apb_rot_ao_and_otp_pwrite               ,
   // Ports for Interface ex_o_rtc_Intr,
   output logic         o_ex_o_rtc_intr_irq                       ,
   // Ports for Interface ex_o_wdt_Intr,
   output logic         o_ex_o_wdt_intr_irq                       ,
   // Ports for Interface ex_smu_axi_fabric_lt_axi_dbgr_m
   input  logic         i_ex_smu_axi_fabric_lt_axi_dbgr_m_arready ,
   input  logic         i_ex_smu_axi_fabric_lt_axi_dbgr_m_awready ,
   input  logic [3:0]   i_ex_smu_axi_fabric_lt_axi_dbgr_m_bid     ,
   input  logic [1:0]   i_ex_smu_axi_fabric_lt_axi_dbgr_m_bresp   ,
   input  logic         i_ex_smu_axi_fabric_lt_axi_dbgr_m_bvalid  ,
   input  logic [63:0]  i_ex_smu_axi_fabric_lt_axi_dbgr_m_rdata   ,
   input  logic [3:0]   i_ex_smu_axi_fabric_lt_axi_dbgr_m_rid     ,
   input  logic         i_ex_smu_axi_fabric_lt_axi_dbgr_m_rlast   ,
   input  logic [1:0]   i_ex_smu_axi_fabric_lt_axi_dbgr_m_rresp   ,
   input  logic         i_ex_smu_axi_fabric_lt_axi_dbgr_m_rvalid  ,
   input  logic         i_ex_smu_axi_fabric_lt_axi_dbgr_m_wready  ,
   output logic [39:0]  o_ex_smu_axi_fabric_lt_axi_dbgr_m_araddr  ,
   output logic [1:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_arburst ,
   output logic [3:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_arcache ,
   output logic [3:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_arid    ,
   output logic [7:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_arlen   ,
   output logic         o_ex_smu_axi_fabric_lt_axi_dbgr_m_arlock  ,
   output logic [2:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_arprot  ,
   output logic [2:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_arsize  ,
   output logic         o_ex_smu_axi_fabric_lt_axi_dbgr_m_arvalid ,
   output logic [39:0]  o_ex_smu_axi_fabric_lt_axi_dbgr_m_awaddr  ,
   output logic [1:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_awburst ,
   output logic [3:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_awcache ,
   output logic [3:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_awid    ,
   output logic [7:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_awlen   ,
   output logic         o_ex_smu_axi_fabric_lt_axi_dbgr_m_awlock  ,
   output logic [2:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_awprot  ,
   output logic [2:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_awsize  ,
   output logic         o_ex_smu_axi_fabric_lt_axi_dbgr_m_awvalid ,
   output logic         o_ex_smu_axi_fabric_lt_axi_dbgr_m_bready  ,
   output logic         o_ex_smu_axi_fabric_lt_axi_dbgr_m_rready  ,
   output logic [63:0]  o_ex_smu_axi_fabric_lt_axi_dbgr_m_wdata   ,
   output logic         o_ex_smu_axi_fabric_lt_axi_dbgr_m_wlast   ,
   output logic [7:0]   o_ex_smu_axi_fabric_lt_axi_dbgr_m_wstrb   ,
   output logic         o_ex_smu_axi_fabric_lt_axi_dbgr_m_wvalid  ,
   // Ports for Interface ext_axi_x2h_m_kse_,
   input  logic [31:0]  i_ext_axi_x2h_m_kse_hrdata                ,
   input  logic         i_ext_axi_x2h_m_kse_hready                ,
   input  logic [1:0]   i_ext_axi_x2h_m_kse_hresp                 ,
   output logic [31:0]  o_ext_axi_x2h_m_kse_haddr                 ,
   output logic [2:0]   o_ext_axi_x2h_m_kse_hburst                ,
   output logic         o_ext_axi_x2h_m_kse_hlock                 ,
   output logic [3:0]   o_ext_axi_x2h_m_kse_hprot                 ,
   output logic [2:0]   o_ext_axi_x2h_m_kse_hsize                 ,
   output logic [1:0]   o_ext_axi_x2h_m_kse_htrans                ,
   output logic [31:0]  o_ext_axi_x2h_m_kse_hwdata                ,
   output logic         o_ext_axi_x2h_m_kse_hwrite                ,
   // Ports for Interface ext_smu_fabric_lt_axi_s,
   input  logic [39:0]  i_ext_smu_fabric_lt_axi_s_araddr          ,
   input  logic [1:0]   i_ext_smu_fabric_lt_axi_s_arburst         ,
   input  logic [3:0]   i_ext_smu_fabric_lt_axi_s_arcache         ,
   input  logic [3:0]   i_ext_smu_fabric_lt_axi_s_arid            ,
   input  logic [7:0]   i_ext_smu_fabric_lt_axi_s_arlen           ,
   input  logic         i_ext_smu_fabric_lt_axi_s_arlock          ,
   input  logic [2:0]   i_ext_smu_fabric_lt_axi_s_arprot          ,
   input  logic [2:0]   i_ext_smu_fabric_lt_axi_s_arsize          ,
   input  logic         i_ext_smu_fabric_lt_axi_s_arvalid         ,
   input  logic [39:0]  i_ext_smu_fabric_lt_axi_s_awaddr          ,
   input  logic [1:0]   i_ext_smu_fabric_lt_axi_s_awburst         ,
   input  logic [3:0]   i_ext_smu_fabric_lt_axi_s_awcache         ,
   input  logic [3:0]   i_ext_smu_fabric_lt_axi_s_awid            ,
   input  logic [7:0]   i_ext_smu_fabric_lt_axi_s_awlen           ,
   input  logic         i_ext_smu_fabric_lt_axi_s_awlock          ,
   input  logic [2:0]   i_ext_smu_fabric_lt_axi_s_awprot          ,
   input  logic [2:0]   i_ext_smu_fabric_lt_axi_s_awsize          ,
   input  logic         i_ext_smu_fabric_lt_axi_s_awvalid         ,
   input  logic         i_ext_smu_fabric_lt_axi_s_bready          ,
   input  logic         i_ext_smu_fabric_lt_axi_s_rready          ,
   input  logic [63:0]  i_ext_smu_fabric_lt_axi_s_wdata           ,
   input  logic         i_ext_smu_fabric_lt_axi_s_wlast           ,
   input  logic [7:0]   i_ext_smu_fabric_lt_axi_s_wstrb           ,
   input  logic         i_ext_smu_fabric_lt_axi_s_wvalid          ,
   output logic         o_ext_smu_fabric_lt_axi_s_arready         ,
   output logic         o_ext_smu_fabric_lt_axi_s_awready         ,
   output logic [3:0]   o_ext_smu_fabric_lt_axi_s_bid             ,
   output logic [1:0]   o_ext_smu_fabric_lt_axi_s_bresp           ,
   output logic         o_ext_smu_fabric_lt_axi_s_bvalid          ,
   output logic [63:0]  o_ext_smu_fabric_lt_axi_s_rdata           ,
   output logic [3:0]   o_ext_smu_fabric_lt_axi_s_rid             ,
   output logic         o_ext_smu_fabric_lt_axi_s_rlast           ,
   output logic [1:0]   o_ext_smu_fabric_lt_axi_s_rresp           ,
   output logic         o_ext_smu_fabric_lt_axi_s_rvalid          ,
   output logic         o_ext_smu_fabric_lt_axi_s_wready          ,
   // Ports for Manually exported pins
   input  wire          i_rtc_rtc_clk                             ,
   input  wire          i_rtc_rtc_fpclk                           ,
   input  wire          i_rtc_rtc_rst_n                           ,
   input  logic         i_rtc_scan_mode                           ,
   input  logic         i_wdt_scan_mode                           ,
   input  logic         i_wdt_speed_up                            ,
   input  logic         i_wdt_pause                               ,
   output logic         o_wdt_wdt_sys_rst                         ,
   output logic         o_smu_axi_fabric_dbg_active_trans         ,
   output logic [39:0]  o_smu_axi_fabric_dbg_araddr_s0            ,
   output logic [1:0]   o_smu_axi_fabric_dbg_arburst_s0           ,
   output logic [3:0]   o_smu_axi_fabric_dbg_arcache_s0           ,
   output logic [3:0]   o_smu_axi_fabric_dbg_arid_s0              ,
   output logic [7:0]   o_smu_axi_fabric_dbg_arlen_s0             ,
   output logic         o_smu_axi_fabric_dbg_arlock_s0            ,
   output logic [2:0]   o_smu_axi_fabric_dbg_arprot_s0            ,
   output logic         o_smu_axi_fabric_dbg_arready_s0           ,
   output logic [2:0]   o_smu_axi_fabric_dbg_arsize_s0            ,
   output logic         o_smu_axi_fabric_dbg_arvalid_s0           ,
   output logic [39:0]  o_smu_axi_fabric_dbg_awaddr_s0            ,
   output logic [1:0]   o_smu_axi_fabric_dbg_awburst_s0           ,
   output logic [3:0]   o_smu_axi_fabric_dbg_awcache_s0           ,
   output logic [3:0]   o_smu_axi_fabric_dbg_awid_s0              ,
   output logic [7:0]   o_smu_axi_fabric_dbg_awlen_s0             ,
   output logic         o_smu_axi_fabric_dbg_awlock_s0            ,
   output logic [2:0]   o_smu_axi_fabric_dbg_awprot_s0            ,
   output logic         o_smu_axi_fabric_dbg_awready_s0           ,
   output logic [2:0]   o_smu_axi_fabric_dbg_awsize_s0            ,
   output logic         o_smu_axi_fabric_dbg_awvalid_s0           ,
   output logic [3:0]   o_smu_axi_fabric_dbg_bid_s0               ,
   output logic         o_smu_axi_fabric_dbg_bready_s0            ,
   output logic [1:0]   o_smu_axi_fabric_dbg_bresp_s0             ,
   output logic         o_smu_axi_fabric_dbg_bvalid_s0            ,
   output logic [63:0]  o_smu_axi_fabric_dbg_rdata_s0             ,
   output logic [3:0]   o_smu_axi_fabric_dbg_rid_s0               ,
   output logic         o_smu_axi_fabric_dbg_rlast_s0             ,
   output logic         o_smu_axi_fabric_dbg_rready_s0            ,
   output logic [1:0]   o_smu_axi_fabric_dbg_rresp_s0             ,
   output logic         o_smu_axi_fabric_dbg_rvalid_s0            ,
   output logic [63:0]  o_smu_axi_fabric_dbg_wdata_s0             ,
   output logic [3:0]   o_smu_axi_fabric_dbg_wid_s0               ,
   output logic         o_smu_axi_fabric_dbg_wlast_s0             ,
   output logic         o_smu_axi_fabric_dbg_wready_s0            ,
   output logic [7:0]   o_smu_axi_fabric_dbg_wstrb_s0             ,
   output logic         o_smu_axi_fabric_dbg_wvalid_s0
);


  //============================================================================
  smu_fabric_subsys u_smu_fabric_subsys (
    .aclk                                        ( i_aclk                                        ),
    .aresetn                                     ( i_aresetn                                     ),
    .hclk                                        ( i_hclk                                        ),
    .hresetn                                     ( i_hresetn                                     ),
    .pclk                                        ( i_pclk                                        ),
    .presetn                                     ( i_presetn                                     ),
    // Ports for Interface ex_apb_mbist
    .ex_apb_mbist_prdata                         ( i_mbist_prdata                                ),
    .ex_apb_mbist_pready                         ( i_apb_mbist_pready                            ),
    .ex_apb_mbist_pslverr                        ( i_apb_mbist_pslverr                           ),
    .ex_apb_mbist_paddr                          ( o_mbist_paddr                                 ),
    .ex_apb_mbist_penable                        ( o_mbist_penable                               ),
    .ex_apb_mbist_psel                           ( o_mbist_psel                                  ),
    .ex_apb_mbist_pwdata                         ( o_mbist_pwdata                                ),
    .ex_apb_mbist_pwrite                         ( o_mbist_pwrite                                ),
    // Ports for Interface ex_i_apb_rot_
    .ex_i_apb_tms_prdata                         ( i_apb_tms_prdata                             ),
    .ex_i_apb_tms_pready                         ( i_apb_tms_pready                             ),
    .ex_i_apb_tms_pslverr                        ( i_apb_tms_pslverr                            ),
    .ex_i_apb_tms_paddr                          ( o_apb_tms_csr_paddr                          ),
    .ex_i_apb_tms_penable                        ( o_apb_tms_csr_penable                        ),
    .ex_i_apb_tms_psel                           ( o_apb_tms_csr_psel                           ),
    .ex_i_apb_tms_pwdata                         ( o_apb_tms_csr_pwdata                         ),
    .ex_i_apb_tms_pwrite                         ( o_apb_tms_csr_pwrite                         ),
    // Ports for Interface ex_i_axi_x2p_otp
    .ex_i_axi_x2p_otp_prdata                     ( i_apb_rot_ao_and_otp_prdata                   ),
    .ex_i_axi_x2p_otp_pready                     ( i_apb_rot_ao_and_otp_pready                   ),
    .ex_i_axi_x2p_otp_pslverr                    ( i_apb_rot_ao_and_otp_pslverr                  ),
    .ex_i_axi_x2p_otp_paddr                      ( o_apb_rot_ao_and_otp_paddr                    ),
    .ex_i_axi_x2p_otp_penable                    ( o_apb_rot_ao_and_otp_penable                  ),
    .ex_i_axi_x2p_otp_psel                       ( o_apb_rot_ao_and_otp_psel                     ),
    .ex_i_axi_x2p_otp_pwdata                     ( o_apb_rot_ao_and_otp_pwdata                   ),
    .ex_i_axi_x2p_otp_pwrite                     ( o_apb_rot_ao_and_otp_pwrite                   ),

    .ex_o_rtc_Intr_irq                           ( o_ex_o_rtc_intr_irq                           ),
    .ex_o_wdt_Intr_irq                           ( o_ex_o_wdt_intr_irq                           ),

    // LT AXI Debugger master interface
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arready     ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_arready     ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awready     ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_awready     ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_bid         ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_bid         ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_bresp       ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_bresp       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_bvalid      ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_bvalid      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_rdata       ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_rdata       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_rid         ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_rid         ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_rlast       ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_rlast       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_rresp       ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_rresp       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_rvalid      ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_rvalid      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_wready      ( i_ex_smu_axi_fabric_lt_axi_dbgr_m_wready      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_araddr      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_araddr      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arburst     ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_arburst     ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arcache     ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_arcache     ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arid        ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_arid        ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arlen       ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_arlen       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arlock      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_arlock      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arprot      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_arprot      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arsize      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_arsize      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_arvalid     ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_arvalid     ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awaddr      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awaddr      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awburst     ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awburst     ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awcache     ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awcache     ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awid        ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awid        ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awlen       ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awlen       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awlock      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awlock      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awprot      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awprot      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awsize      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awsize      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_awvalid     ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_awvalid     ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_bready      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_bready      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_rready      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_rready      ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_wdata       ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_wdata       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_wlast       ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_wlast       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_wstrb       ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_wstrb       ),
    .ex_smu_axi_fabric_lt_axi_dbgr_m_wvalid      ( o_ex_smu_axi_fabric_lt_axi_dbgr_m_wvalid      ),
    // Ports for Interface ext_axi_x2h_m_kse_
    .ext_axi_x2h_m_kse_hrdata                    ( i_ext_axi_x2h_m_kse_hrdata                    ),
    .ext_axi_x2h_m_kse_hready                    ( i_ext_axi_x2h_m_kse_hready                    ),
    .ext_axi_x2h_m_kse_hresp                     ( i_ext_axi_x2h_m_kse_hresp                     ),
    .ext_axi_x2h_m_kse_haddr                     ( o_ext_axi_x2h_m_kse_haddr                     ),
    .ext_axi_x2h_m_kse_hburst                    ( o_ext_axi_x2h_m_kse_hburst                    ),
    .ext_axi_x2h_m_kse_hlock                     ( o_ext_axi_x2h_m_kse_hlock                     ),
    .ext_axi_x2h_m_kse_hprot                     ( o_ext_axi_x2h_m_kse_hprot                     ),
    .ext_axi_x2h_m_kse_hsize                     ( o_ext_axi_x2h_m_kse_hsize                     ),
    .ext_axi_x2h_m_kse_htrans                    ( o_ext_axi_x2h_m_kse_htrans                    ),
    .ext_axi_x2h_m_kse_hwdata                    ( o_ext_axi_x2h_m_kse_hwdata                    ),
    .ext_axi_x2h_m_kse_hwrite                    ( o_ext_axi_x2h_m_kse_hwrite                    ),
    // Ports for Interface ext_smu_fabric_lt_axi_s
    .ext_smu_fabric_lt_axi_s_araddr              ( i_ext_smu_fabric_lt_axi_s_araddr              ),
    .ext_smu_fabric_lt_axi_s_arburst             ( i_ext_smu_fabric_lt_axi_s_arburst             ),
    .ext_smu_fabric_lt_axi_s_arcache             ( i_ext_smu_fabric_lt_axi_s_arcache             ),
    .ext_smu_fabric_lt_axi_s_arid                ( i_ext_smu_fabric_lt_axi_s_arid                ),
    .ext_smu_fabric_lt_axi_s_arlen               ( i_ext_smu_fabric_lt_axi_s_arlen               ),
    .ext_smu_fabric_lt_axi_s_arlock              ( i_ext_smu_fabric_lt_axi_s_arlock              ),
    .ext_smu_fabric_lt_axi_s_arprot              ( i_ext_smu_fabric_lt_axi_s_arprot              ),
    .ext_smu_fabric_lt_axi_s_arsize              ( i_ext_smu_fabric_lt_axi_s_arsize              ),
    .ext_smu_fabric_lt_axi_s_arvalid             ( i_ext_smu_fabric_lt_axi_s_arvalid             ),
    .ext_smu_fabric_lt_axi_s_awaddr              ( i_ext_smu_fabric_lt_axi_s_awaddr              ),
    .ext_smu_fabric_lt_axi_s_awburst             ( i_ext_smu_fabric_lt_axi_s_awburst             ),
    .ext_smu_fabric_lt_axi_s_awcache             ( i_ext_smu_fabric_lt_axi_s_awcache             ),
    .ext_smu_fabric_lt_axi_s_awid                ( i_ext_smu_fabric_lt_axi_s_awid                ),
    .ext_smu_fabric_lt_axi_s_awlen               ( i_ext_smu_fabric_lt_axi_s_awlen               ),
    .ext_smu_fabric_lt_axi_s_awlock              ( i_ext_smu_fabric_lt_axi_s_awlock              ),
    .ext_smu_fabric_lt_axi_s_awprot              ( i_ext_smu_fabric_lt_axi_s_awprot              ),
    .ext_smu_fabric_lt_axi_s_awsize              ( i_ext_smu_fabric_lt_axi_s_awsize              ),
    .ext_smu_fabric_lt_axi_s_awvalid             ( i_ext_smu_fabric_lt_axi_s_awvalid             ),
    .ext_smu_fabric_lt_axi_s_bready              ( i_ext_smu_fabric_lt_axi_s_bready              ),
    .ext_smu_fabric_lt_axi_s_rready              ( i_ext_smu_fabric_lt_axi_s_rready              ),
    .ext_smu_fabric_lt_axi_s_wdata               ( i_ext_smu_fabric_lt_axi_s_wdata               ),
    .ext_smu_fabric_lt_axi_s_wlast               ( i_ext_smu_fabric_lt_axi_s_wlast               ),
    .ext_smu_fabric_lt_axi_s_wstrb               ( i_ext_smu_fabric_lt_axi_s_wstrb               ),
    .ext_smu_fabric_lt_axi_s_wvalid              ( i_ext_smu_fabric_lt_axi_s_wvalid              ),
    .ext_smu_fabric_lt_axi_s_arready             ( o_ext_smu_fabric_lt_axi_s_arready             ),
    .ext_smu_fabric_lt_axi_s_awready             ( o_ext_smu_fabric_lt_axi_s_awready             ),
    .ext_smu_fabric_lt_axi_s_bid                 ( o_ext_smu_fabric_lt_axi_s_bid                 ),
    .ext_smu_fabric_lt_axi_s_bresp               ( o_ext_smu_fabric_lt_axi_s_bresp               ),
    .ext_smu_fabric_lt_axi_s_bvalid              ( o_ext_smu_fabric_lt_axi_s_bvalid              ),
    .ext_smu_fabric_lt_axi_s_rdata               ( o_ext_smu_fabric_lt_axi_s_rdata               ),
    .ext_smu_fabric_lt_axi_s_rid                 ( o_ext_smu_fabric_lt_axi_s_rid                 ),
    .ext_smu_fabric_lt_axi_s_rlast               ( o_ext_smu_fabric_lt_axi_s_rlast               ),
    .ext_smu_fabric_lt_axi_s_rresp               ( o_ext_smu_fabric_lt_axi_s_rresp               ),
    .ext_smu_fabric_lt_axi_s_rvalid              ( o_ext_smu_fabric_lt_axi_s_rvalid              ),
    .ext_smu_fabric_lt_axi_s_wready              ( o_ext_smu_fabric_lt_axi_s_wready              ),

    .i_rtc_rtc_clk                               ( i_rtc_rtc_clk                                 ),
    .i_rtc_rtc_fpclk                             ( i_rtc_rtc_fpclk                               ),
    .i_rtc_rtc_rst_n                             ( i_rtc_rtc_rst_n                               ),
    .i_rtc_scan_mode                             ( i_rtc_scan_mode                               ),
    .i_wdt_scan_mode                             ( i_wdt_scan_mode                               ),
    .i_wdt_speed_up                              ( i_wdt_speed_up                                ),
    .i_wdt_pause                                 ( i_wdt_pause                                   ),
    .i_wdt_wdt_sys_rst                           ( o_wdt_wdt_sys_rst                             ),
    .smu_axi_fabric_dbg_active_trans             ( o_smu_axi_fabric_dbg_active_trans             ),
    .smu_axi_fabric_dbg_araddr_s0                ( o_smu_axi_fabric_dbg_araddr_s0                ),
    .smu_axi_fabric_dbg_arburst_s0               ( o_smu_axi_fabric_dbg_arburst_s0               ),
    .smu_axi_fabric_dbg_arcache_s0               ( o_smu_axi_fabric_dbg_arcache_s0               ),
    .smu_axi_fabric_dbg_arid_s0                  ( o_smu_axi_fabric_dbg_arid_s0                  ),
    .smu_axi_fabric_dbg_arlen_s0                 ( o_smu_axi_fabric_dbg_arlen_s0                 ),
    .smu_axi_fabric_dbg_arlock_s0                ( o_smu_axi_fabric_dbg_arlock_s0                ),
    .smu_axi_fabric_dbg_arprot_s0                ( o_smu_axi_fabric_dbg_arprot_s0                ),
    .smu_axi_fabric_dbg_arready_s0               ( o_smu_axi_fabric_dbg_arready_s0               ),
    .smu_axi_fabric_dbg_arsize_s0                ( o_smu_axi_fabric_dbg_arsize_s0                ),
    .smu_axi_fabric_dbg_arvalid_s0               ( o_smu_axi_fabric_dbg_arvalid_s0               ),
    .smu_axi_fabric_dbg_awaddr_s0                ( o_smu_axi_fabric_dbg_awaddr_s0                ),
    .smu_axi_fabric_dbg_awburst_s0               ( o_smu_axi_fabric_dbg_awburst_s0               ),
    .smu_axi_fabric_dbg_awcache_s0               ( o_smu_axi_fabric_dbg_awcache_s0               ),
    .smu_axi_fabric_dbg_awid_s0                  ( o_smu_axi_fabric_dbg_awid_s0                  ),
    .smu_axi_fabric_dbg_awlen_s0                 ( o_smu_axi_fabric_dbg_awlen_s0                 ),
    .smu_axi_fabric_dbg_awlock_s0                ( o_smu_axi_fabric_dbg_awlock_s0                ),
    .smu_axi_fabric_dbg_awprot_s0                ( o_smu_axi_fabric_dbg_awprot_s0                ),
    .smu_axi_fabric_dbg_awready_s0               ( o_smu_axi_fabric_dbg_awready_s0               ),
    .smu_axi_fabric_dbg_awsize_s0                ( o_smu_axi_fabric_dbg_awsize_s0                ),
    .smu_axi_fabric_dbg_awvalid_s0               ( o_smu_axi_fabric_dbg_awvalid_s0               ),
    .smu_axi_fabric_dbg_bid_s0                   ( o_smu_axi_fabric_dbg_bid_s0                   ),
    .smu_axi_fabric_dbg_bready_s0                ( o_smu_axi_fabric_dbg_bready_s0                ),
    .smu_axi_fabric_dbg_bresp_s0                 ( o_smu_axi_fabric_dbg_bresp_s0                 ),
    .smu_axi_fabric_dbg_bvalid_s0                ( o_smu_axi_fabric_dbg_bvalid_s0                ),
    .smu_axi_fabric_dbg_rdata_s0                 ( o_smu_axi_fabric_dbg_rdata_s0                 ),
    .smu_axi_fabric_dbg_rid_s0                   ( o_smu_axi_fabric_dbg_rid_s0                   ),
    .smu_axi_fabric_dbg_rlast_s0                 ( o_smu_axi_fabric_dbg_rlast_s0                 ),
    .smu_axi_fabric_dbg_rready_s0                ( o_smu_axi_fabric_dbg_rready_s0                ),
    .smu_axi_fabric_dbg_rresp_s0                 ( o_smu_axi_fabric_dbg_rresp_s0                 ),
    .smu_axi_fabric_dbg_rvalid_s0                ( o_smu_axi_fabric_dbg_rvalid_s0                ),
    .smu_axi_fabric_dbg_wdata_s0                 ( o_smu_axi_fabric_dbg_wdata_s0                 ),
    .smu_axi_fabric_dbg_wid_s0                   ( o_smu_axi_fabric_dbg_wid_s0                   ),
    .smu_axi_fabric_dbg_wlast_s0                 ( o_smu_axi_fabric_dbg_wlast_s0                 ),
    .smu_axi_fabric_dbg_wready_s0                ( o_smu_axi_fabric_dbg_wready_s0                ),
    .smu_axi_fabric_dbg_wstrb_s0                 ( o_smu_axi_fabric_dbg_wstrb_s0                 ),
    .smu_axi_fabric_dbg_wvalid_s0                ( o_smu_axi_fabric_dbg_wvalid_s0                )
  );

endmodule
