// (C) Copyright Axelera AI 2023
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description:  Verification Utility Package
//  Put here common classes useful for verification
// Owner: Raymond Garcia <raymond.garcia@axelera.ai>

package v_utils_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "v_object.sv"
    `include "register_access.sv"
endpackage
