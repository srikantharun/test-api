 const phy_init_data_t phy_init_devinit_skiptrain_details[string][] = '{
                  
//[dwc_ddrphy_phyinit_userCustom_A_bringupPower] Start of dwc_ddrphy_phyinit_userCustom_A_bringupPower()
//[dwc_ddrphy_phyinit_userCustom_A_bringupPower] End of dwc_ddrphy_phyinit_userCustom_A_bringupPower()
 
                  
//[dwc_ddrphy_phyinit_userCustom_B_startClockResetPhy] Start of dwc_ddrphy_phyinit_userCustom_B_startClockResetPhy()
//[dwc_ddrphy_phyinit_userCustom_B_startClockResetPhy] End of dwc_ddrphy_phyinit_userCustom_B_startClockResetPhy()
 
   "C" : '{                 
//[phyinit_C_initPhyConfig] Start of dwc_ddrphy_phyinit_C_initPhyConfig()
                          '{ step_type : REG_WRITE, reg_addr : 32'h30022, value : 32'h2}, //[dwc_ddrphy_phyinit_programMemResetL] Programming MemResetL AC0 to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h31022, value : 32'h2}, //[dwc_ddrphy_phyinit_programMemResetL] Programming MemResetL AC1 to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4070, value : 32'hff}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=0, Programming HMAC 4  TxImpedanceAC::CS to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h5070, value : 32'h77}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=0, Programming HMAC 5  TxImpedanceAC::CK to 0x77
                          '{ step_type : REG_WRITE, reg_addr : 32'hb070, value : 32'hff}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=0, Programming HMAC 11 TxImpedanceAC::CS to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'hc070, value : 32'h77}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=0, Programming HMAC 12 TxImpedanceAC::CK to 0x77
                          '{ step_type : REG_WRITE, reg_addr : 32'h104070, value : 32'hff}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=1, Programming HMAC 4  TxImpedanceAC::CS to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h105070, value : 32'h77}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=1, Programming HMAC 5  TxImpedanceAC::CK to 0x77
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b070, value : 32'hff}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=1, Programming HMAC 11 TxImpedanceAC::CS to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c070, value : 32'h77}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=1, Programming HMAC 12 TxImpedanceAC::CK to 0x77
                          '{ step_type : REG_WRITE, reg_addr : 32'h204070, value : 32'hff}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=2, Programming HMAC 4  TxImpedanceAC::CS to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h205070, value : 32'h77}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=2, Programming HMAC 5  TxImpedanceAC::CK to 0x77
                          '{ step_type : REG_WRITE, reg_addr : 32'h20b070, value : 32'hff}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=2, Programming HMAC 11 TxImpedanceAC::CS to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h20c070, value : 32'h77}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=2, Programming HMAC 12 TxImpedanceAC::CK to 0x77
                          '{ step_type : REG_WRITE, reg_addr : 32'h304070, value : 32'hff}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=3, Programming HMAC 4  TxImpedanceAC::CS to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h305070, value : 32'h77}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=3, Programming HMAC 5  TxImpedanceAC::CK to 0x77
                          '{ step_type : REG_WRITE, reg_addr : 32'h30b070, value : 32'hff}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=3, Programming HMAC 11 TxImpedanceAC::CS to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h30c070, value : 32'h77}, //[dwc_ddrphy_phyinit_PowerUp] Pstate=3, Programming HMAC 12 TxImpedanceAC::CK to 0x77
                          '{ step_type : REG_WRITE, reg_addr : 32'h5, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC0 Instance0 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC1 Instance1 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC2 Instance2 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC3 Instance3 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h4005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC4 Instance4 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h5005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC5 Instance5 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h7005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC0 Instance7 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h8005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC1 Instance8 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h9005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC2 Instance9 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'ha005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC3 Instance10 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'hb005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC4 Instance11 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'hc005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC5 Instance12 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'ha0308, value : 32'h2}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMZCAL TxPowerDownZCAL to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'ha0002, value : 32'h1}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMZCAL ZcalPowerCtl.RxPowerDown to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he0046, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownLn0 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he0047, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownLn1 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he0048, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownLn2 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he0049, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownLn3 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he1046, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn0 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he1047, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn1 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he1048, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn2 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he1049, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn3 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he104a, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn4 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he004b, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownDQS TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he104b, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownDQS TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he2046, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownLn0 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he2047, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownLn1 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he2048, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownLn2 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he2049, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownLn3 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he3046, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn0 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he3047, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn1 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he3048, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn2 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he3049, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn3 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he304a, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn4 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he204b, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownDQS TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he304b, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownDQS TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he4046, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownLn0 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he4047, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownLn1 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he4048, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownLn2 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he4049, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownLn3 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he5046, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn0 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he5047, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn1 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he5048, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn2 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he5049, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn3 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he504a, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn4 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he404b, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownDQS TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he504b, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownDQS TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he6046, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownLn0 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he6047, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownLn1 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he6048, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownLn2 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he6049, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownLn3 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he7046, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn0 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he7047, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn1 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he7048, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn2 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he7049, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn3 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he704a, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn4 TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he604b, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownDQS TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'he704b, value : 32'h6}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownDQS TxPowerDown to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h30020, value : 32'h1}, //[dwc_ddrphy_phyinit_PowerUp] Programming PorControl::PwrOkDlyCtrl to 1'b1
                          '{ step_type : REG_WRITE, reg_addr : 32'h31020, value : 32'h1},
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 16},
//Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 16 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'h5, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC0 Instance0 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC1 Instance1 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC2 Instance2 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC3 Instance3 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h4005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC4 Instance4 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h5005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX0 HMAC5 Instance5 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h7005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC0 Instance7 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h8005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC1 Instance8 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h9005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC2 Instance9 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'ha005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC3 Instance10 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'hb005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC4 Instance11 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'hc005, value : 32'h3}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming ACX1 HMAC5 Instance12 RxPowerDownAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'ha0308, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMZCAL TxPowerDownZCAL to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'ha0002, value : 32'h1}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMZCAL ZcalPowerCtl.RxPowerDown to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he0046, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownLn0 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he0047, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownLn1 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he0048, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownLn2 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he0049, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownLn3 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he1046, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn0 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he1047, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn1 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he1048, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn2 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he1049, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn3 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he104a, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownLn4 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he004b, value : 32'h2}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX0 DxRxPowerDownDQS TxPowerDown to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'he104b, value : 32'h4}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE0 DX1 DxRxPowerDownDQS TxPowerDown to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he2046, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownLn0 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he2047, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownLn1 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he2048, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownLn2 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he2049, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownLn3 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he3046, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn0 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he3047, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn1 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he3048, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn2 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he3049, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn3 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he304a, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownLn4 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he204b, value : 32'h2}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX0 DxRxPowerDownDQS TxPowerDown to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'he304b, value : 32'h4}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE1 DX1 DxRxPowerDownDQS TxPowerDown to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he4046, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownLn0 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he4047, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownLn1 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he4048, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownLn2 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he4049, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownLn3 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he5046, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn0 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he5047, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn1 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he5048, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn2 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he5049, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn3 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he504a, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownLn4 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he404b, value : 32'h2}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX0 DxRxPowerDownDQS TxPowerDown to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'he504b, value : 32'h4}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE2 DX1 DxRxPowerDownDQS TxPowerDown to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he6046, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownLn0 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he6047, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownLn1 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he6048, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownLn2 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he6049, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownLn3 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he7046, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn0 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he7047, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn1 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he7048, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn2 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he7049, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn3 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he704a, value : 32'h0}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownLn4 TxPowerDown to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he604b, value : 32'h2}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX0 DxRxPowerDownDQS TxPowerDown to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'he704b, value : 32'h4}, //[dwc_ddrphy_phyinit_setTxRxPowerDown] Programming HMDBYTE3 DX1 DxRxPowerDownDQS TxPowerDown to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h200a5, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming LP5Mode to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h10097, value : 32'h7ff}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE0 DxOdtEn to 0x7ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h11097, value : 32'h7ff}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE1 DxOdtEn to 0x7ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h12097, value : 32'h7ff}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE2 DxOdtEn to 0x7ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h13097, value : 32'h7ff}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE3 DxOdtEn to 0x7ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE0. TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE0. TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE1. TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE1. TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE2. TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE2. TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE3. TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming DBYTE3. TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb0303, value : 32'h9}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ZCalRate::ZCalOnce to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'ha0302, value : 32'h26}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ZCalCompVref::ZCalDACRangeSel to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb0301, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ZCalBaseCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb030f, value : 32'h1d}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ZCalAnaSettlingTime to 0x1d
                          '{ step_type : REG_WRITE, reg_addr : 32'h300ae, value : 32'h1880}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming AC0.AcLnDisable to 0x1880
                          '{ step_type : REG_WRITE, reg_addr : 32'h300ad, value : 32'h1880}, //phyinit_io_write: 0x300ae, 0x1880
                          '{ step_type : REG_WRITE, reg_addr : 32'h300ac, value : 32'h1880}, //phyinit_io_write: 0x300ad, 0x1880
                          '{ step_type : REG_WRITE, reg_addr : 32'h310ae, value : 32'h1880}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming AC1.AcLnDisable to 0x1880
                          '{ step_type : REG_WRITE, reg_addr : 32'h310ad, value : 32'h1880}, //phyinit_io_write: 0x310ae, 0x1880
                          '{ step_type : REG_WRITE, reg_addr : 32'h310ac, value : 32'h1880}, //phyinit_io_write: 0x310ad, 0x1880
                          '{ step_type : REG_WRITE, reg_addr : 32'h100a3, value : 32'h833}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming PptCtlStatic to 0x833
                          '{ step_type : REG_WRITE, reg_addr : 32'h110a3, value : 32'h83f}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming PptCtlStatic to 0x83f
                          '{ step_type : REG_WRITE, reg_addr : 32'h120a3, value : 32'h833}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming PptCtlStatic to 0x833
                          '{ step_type : REG_WRITE, reg_addr : 32'h130a3, value : 32'h83f}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming PptCtlStatic to 0x83f
                          '{ step_type : REG_WRITE, reg_addr : 32'hc00f0, value : 32'h1111}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat[3]=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h90730, value : 32'h688}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat_dp[3]=3
                          '{ step_type : REG_WRITE, reg_addr : 32'hc00f1, value : 32'h2222}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat[7]=2
                          '{ step_type : REG_WRITE, reg_addr : 32'h90731, value : 32'h688}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat_dp[7]=3
                          '{ step_type : REG_WRITE, reg_addr : 32'hc00f2, value : 32'h7777}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat[11]=7
                          '{ step_type : REG_WRITE, reg_addr : 32'h90732, value : 32'h688}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat_dp[11]=3
                          '{ step_type : REG_WRITE, reg_addr : 32'hc00f3, value : 32'h34}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat[15]=0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90733, value : 32'h2d}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat_dp[15]=0
                          '{ step_type : REG_WRITE, reg_addr : 32'hc00f4, value : 32'h5555}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat[19]=5
                          '{ step_type : REG_WRITE, reg_addr : 32'h90734, value : 32'h688}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat_dp[19]=3
                          '{ step_type : REG_WRITE, reg_addr : 32'hc00f7, value : 32'hf000}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat[31]=15
                          '{ step_type : REG_WRITE, reg_addr : 32'h90737, value : 32'ha00}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat_dp[31]=5
                          '{ step_type : REG_WRITE, reg_addr : 32'h9071f, value : 32'h4}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming xlat_dp[63]=0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90829, value : 32'hf}, //phyinit_io_write: 0x9071f, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h20007, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming MASTER.PubDbyteDisable to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he007a, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE 0 DX4 RxModeX8Sel to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he107a, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE 0 DX5 RxModeX8Sel to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he207a, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE 1 DX4 RxModeX8Sel to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he307a, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE 1 DX5 RxModeX8Sel to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he407a, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE 2 DX4 RxModeX8Sel to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he507a, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE 2 DX5 RxModeX8Sel to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he607a, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE 3 DX4 RxModeX8Sel to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he707a, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE 3 DX5 RxModeX8Sel to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h61e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC0 Instance0 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h161e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC1 Instance1 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h261e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC2 Instance2 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h361e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC3 Instance3 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h461e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC4 Instance4 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h561e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC5 Instance5 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h761e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC0 Instance7 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h861e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC1 Instance8 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h961e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC2 Instance9 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'ha61e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC3 Instance10 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb61e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC4 Instance11 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hc61e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC5 Instance12 PclkDCAClkGaterEnAC/DB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10e1f, value : 32'h0}, //phyinit_io_write: 0xc61e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11e1f, value : 32'h0}, //phyinit_io_write: 0x10e1f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h12e1f, value : 32'h0}, //phyinit_io_write: 0x11e1f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h13e1f, value : 32'h0}, //phyinit_io_write: 0x12e1f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30807, value : 32'hee66}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming PclkDCANextFineOnCoarseAC/DB Full Search to 0xee66
                          '{ step_type : REG_WRITE, reg_addr : 32'h31807, value : 32'hee66}, //phyinit_io_write: 0x30807, 0xee66
                          '{ step_type : REG_WRITE, reg_addr : 32'h10807, value : 32'hee66}, //phyinit_io_write: 0x31807, 0xee66
                          '{ step_type : REG_WRITE, reg_addr : 32'h11807, value : 32'hee66}, //phyinit_io_write: 0x10807, 0xee66
                          '{ step_type : REG_WRITE, reg_addr : 32'h12807, value : 32'hee66}, //phyinit_io_write: 0x11807, 0xee66
                          '{ step_type : REG_WRITE, reg_addr : 32'h13807, value : 32'hee66}, //phyinit_io_write: 0x12807, 0xee66
                          '{ step_type : REG_WRITE, reg_addr : 32'h300a0, value : 32'h3fff}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming AC0.AsyncAcTxMode to 0x3fff
                          '{ step_type : REG_WRITE, reg_addr : 32'h310a0, value : 32'h3fff}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming AC1.AsyncAcTxMode to 0x3fff
                          '{ step_type : REG_WRITE, reg_addr : 32'h10089, value : 32'h1fff}, //phyinit_io_write: 0x310a0, 0x3fff
                          '{ step_type : REG_WRITE, reg_addr : 32'h1008a, value : 32'h7ff}, //phyinit_io_write: 0x10089, 0x1fff
                          '{ step_type : REG_WRITE, reg_addr : 32'h11089, value : 32'h1fff}, //phyinit_io_write: 0x1008a, 0x7ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h1108a, value : 32'h7ff}, //phyinit_io_write: 0x11089, 0x1fff
                          '{ step_type : REG_WRITE, reg_addr : 32'h12089, value : 32'h1fff}, //phyinit_io_write: 0x1108a, 0x7ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h1208a, value : 32'h7ff}, //phyinit_io_write: 0x12089, 0x1fff
                          '{ step_type : REG_WRITE, reg_addr : 32'h13089, value : 32'h1fff}, //phyinit_io_write: 0x1208a, 0x7ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h1308a, value : 32'h7ff}, //phyinit_io_write: 0x13089, 0x1fff
                          '{ step_type : REG_WRITE, reg_addr : 32'h20006, value : 32'hf}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming LpDqPhaseDisable to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h2000c, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming PipeNetDis to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he000d, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE0 RxGainCtrl to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he100d, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE1 RxGainCtrl to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he200d, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE2 RxGainCtrl to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he300d, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE3 RxGainCtrl to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he400d, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE4 RxGainCtrl to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he500d, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE5 RxGainCtrl to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he600d, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE6 RxGainCtrl to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he700d, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming HMDBYTE7 RxGainCtrl to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h30027, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACDlyScaleGatingDisable AC0 to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC0 Instance0 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h103f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC1 Instance1 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h203f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC2 Instance2 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h303f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC3 Instance3 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h403f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC4 Instance4 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX0 HMAC5 Instance5 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h31027, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACDlyScaleGatingDisable AC1 to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h703f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC0 Instance7 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h803f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC1 Instance8 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h903f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC2 Instance9 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'ha03f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC3 Instance10 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'hb03f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC4 Instance11 to NeverGateACDlyScaleValClk 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'hc03f, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfig] Programming ACX1 HMAC5 Instance12 to NeverGateACDlyScaleValClk 0x1
//[dwc_ddrphy_phyinit_programDfiMode] Skip DfiMode Programming: Keeping the reset value of 0x3
//[phyinit_C_initPhyConfig] End of dwc_ddrphy_phyinit_C_initPhyConfig()
//[dwc_ddrphy_phyinit_sequence] initCtrl = 33
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0080, value : 32'h5}    },
   "D" : '{                 
// [dwc_ddrphy_phyinit_D_loadIMEM] Start of dwc_ddrphy_phyinit_D_loadIMEM
                          '{ step_type : REG_WRITE, reg_addr : 32'h50000, value : 32'h58c}, // [dwc_ddrphy_phyinit_WriteOutMem] STARTING. offset 0x50000 size 0x53a4, sparse_write=0
                          '{ step_type : REG_WRITE, reg_addr : 32'h50001, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50002, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50003, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50004, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50005, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50006, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50007, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50008, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50009, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5000a, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5000b, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5000c, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5000d, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5000e, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5000f, value : 32'h90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50010, value : 32'h50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50011, value : 32'h50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50012, value : 32'h50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50013, value : 32'h50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50014, value : 32'h7000264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50015, value : 32'h7000264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50016, value : 32'h7000264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50017, value : 32'h7000264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50018, value : 32'h402069},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50019, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5001a, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5001b, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5001c, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5001d, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5001e, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5001f, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50020, value : 32'hc0d1c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50021, value : 32'h7ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50022, value : 32'hc0d1c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50023, value : 32'h7ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50024, value : 32'hf80220a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50025, value : 32'h8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50026, value : 32'hf80230a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50027, value : 32'hdead1234},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50028, value : 32'hc01a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50029, value : 32'h23aa7444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5002a, value : 32'h1a000010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5002b, value : 32'h744400c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5002c, value : 32'hd023aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5002d, value : 32'hc01a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5002e, value : 32'h1a007444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5002f, value : 32'h74440000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50030, value : 32'h401a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50031, value : 32'h1a007444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50032, value : 32'h74440700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50033, value : 32'h6c01a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50034, value : 32'h230a7444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50035, value : 32'habcd0f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50036, value : 32'h1a00dead},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50037, value : 32'h206900c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50038, value : 32'h78e00040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50039, value : 32'h803c2242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5003a, value : 32'h42007ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5003b, value : 32'h18020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5003c, value : 32'h4831101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5003d, value : 32'hd21a01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5003e, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5003f, value : 32'h803c2242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50040, value : 32'h42007ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50041, value : 32'h10020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50042, value : 32'h521a01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50043, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50044, value : 32'hb6881cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50045, value : 32'hb6481cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50046, value : 32'hb6081cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50047, value : 32'hb5c81cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50048, value : 32'hb5881cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50049, value : 32'hb5481cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5004a, value : 32'hb5081cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5004b, value : 32'hb4c81cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5004c, value : 32'hb4881cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5004d, value : 32'hb4481cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5004e, value : 32'hb4081cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5004f, value : 32'hb3c81cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50050, value : 32'hb3881cfc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50051, value : 32'h1cfc7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50052, value : 32'h78e0b348},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50053, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50054, value : 32'hdd38748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50055, value : 32'h78e0f038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50056, value : 32'hdd34748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50057, value : 32'h78e0f036},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50058, value : 32'hdd30748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50059, value : 32'h78e0f034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5005a, value : 32'hdd2c748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5005b, value : 32'h78e0f032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5005c, value : 32'hdd28748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5005d, value : 32'h78e0f030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5005e, value : 32'hdd24748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5005f, value : 32'h78e0f02e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50060, value : 32'hdd20748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50061, value : 32'h78e0f02c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50062, value : 32'hdd1c748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50063, value : 32'h78e0f02a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50064, value : 32'hdd18748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50065, value : 32'h78e0f028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50066, value : 32'hdd14748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50067, value : 32'h78e0f026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50068, value : 32'hdd10748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50069, value : 32'h78e0f024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5006a, value : 32'hdd0c748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5006b, value : 32'h78e0f022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5006c, value : 32'hdd08748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5006d, value : 32'h78e0f01f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5006e, value : 32'h74ad748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5006f, value : 32'h78e0f01c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50070, value : 32'hf01c748d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50071, value : 32'h301a1434},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50072, value : 32'h30191430},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50073, value : 32'h3018142c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50074, value : 32'h30171428},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50075, value : 32'h30161424},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50076, value : 32'h30151420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50077, value : 32'h3014141c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50078, value : 32'h30131418},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50079, value : 32'h30121414},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5007a, value : 32'h30111410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5007b, value : 32'h3010140c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5007c, value : 32'hc601c702},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5007d, value : 32'h334d24b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5007e, value : 32'h331f24b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5007f, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50080, value : 32'h1cfcc4c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50081, value : 32'h1cfcb1c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50082, value : 32'h1cfcb188},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50083, value : 32'h1cfcb148},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50084, value : 32'hc3e1b108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50085, value : 32'hc1e1c2e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50086, value : 32'hc4e1c0e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50087, value : 32'hc0017fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50088, value : 32'ha11c2f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50089, value : 32'h42300032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5008a, value : 32'h81292f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5008b, value : 32'hf00369e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5008c, value : 32'h280070ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5008d, value : 32'h274e03d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5008e, value : 32'h2a011800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5008f, value : 32'h70f52000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50090, value : 32'h3d02a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50091, value : 32'h200921c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50092, value : 32'h240e2841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50093, value : 32'hab24022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50094, value : 32'h41c10020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50095, value : 32'h23c22a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50096, value : 32'h42d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50097, value : 32'h4508ffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50098, value : 32'hba307f50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50099, value : 32'h2408232f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5009a, value : 32'h20542240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5009b, value : 32'h23640a13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5009c, value : 32'h4002940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5009d, value : 32'h14c3251a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5009e, value : 32'h80f6058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5009f, value : 32'h61d900c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a0, value : 32'h852409ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a1, value : 32'h294077a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a2, value : 32'h251a2411},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a3, value : 32'h72221400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a4, value : 32'ha6e4a10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a5, value : 32'h41c10020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a6, value : 32'ha154300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a7, value : 32'h294020e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a8, value : 32'h231a0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500a9, value : 32'h60f804c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500aa, value : 32'h85080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ab, value : 32'h9ef61d9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ac, value : 32'h77648524},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ad, value : 32'h14002d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ae, value : 32'h2000bd30},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500af, value : 32'h254180c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b0, value : 32'hc6d09001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b1, value : 32'heb884408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b2, value : 32'ha5090d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b3, value : 32'h7554020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b4, value : 32'h4181ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b5, value : 32'h200071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b6, value : 32'h78e04081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b7, value : 32'h4548c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b8, value : 32'h44084220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500b9, value : 32'h41407034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ba, value : 32'h700cf646},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500bb, value : 32'h900c240e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500bc, value : 32'h80812003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500bd, value : 32'h330b11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500be, value : 32'h700c4668},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500bf, value : 32'h900d250e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c0, value : 32'h80ce2003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c1, value : 32'h7cf2b41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c2, value : 32'h7d02a41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c3, value : 32'h917ee8b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c4, value : 32'h40200365},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c5, value : 32'h42a14181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c6, value : 32'h2007ffc2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c7, value : 32'hf40ea3fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c8, value : 32'h4081c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500c9, value : 32'h82242a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ca, value : 32'h43c10020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500cb, value : 32'ha3fe2007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500cc, value : 32'h2505f3f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500cd, value : 32'hf3f693be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ce, value : 32'h200e704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500cf, value : 32'h22038080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d0, value : 32'hc6c88041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d1, value : 32'h200031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d2, value : 32'h78e0708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d3, value : 32'hc42107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d4, value : 32'hf040262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d5, value : 32'h1270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d6, value : 32'h242f0026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d7, value : 32'h200e0104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d8, value : 32'h25038140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500d9, value : 32'h70740041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500da, value : 32'h3000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500db, value : 32'h8142220e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500dc, value : 32'hc32503},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500dd, value : 32'h80852305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500de, value : 32'h10116},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500df, value : 32'h44484368},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e0, value : 32'h43204200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e1, value : 32'h82c0250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e2, value : 32'h1a704d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e3, value : 32'h22c00004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e4, value : 32'h25ca1821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e5, value : 32'h2f2f8301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e6, value : 32'h22c00141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e7, value : 32'h22c01063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e8, value : 32'h70ec11c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500e9, value : 32'h80c0250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ea, value : 32'h82127c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500eb, value : 32'h40014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ec, value : 32'h808125ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ed, value : 32'h141282f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ee, value : 32'h6327c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ef, value : 32'h327c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f0, value : 32'h8287270e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f1, value : 32'h2427ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f2, value : 32'h45e071e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f3, value : 32'h8800274c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f4, value : 32'h12702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f5, value : 32'h700c0024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f6, value : 32'h42604140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f7, value : 32'h2742706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f8, value : 32'h240a8807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500f9, value : 32'h2a7140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500fa, value : 32'h274e0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500fb, value : 32'h7c880a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500fc, value : 32'h29000001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500fd, value : 32'h29010280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500fe, value : 32'h2a0001c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h500ff, value : 32'h71a00285},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50100, value : 32'h1c22a01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50101, value : 32'h2852b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50102, value : 32'h1c32b01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50103, value : 32'h224c72a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50104, value : 32'h629800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50105, value : 32'h20a80009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50106, value : 32'h200005c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50107, value : 32'h21018000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50108, value : 32'h22018041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50109, value : 32'h23018082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5010a, value : 32'h220200c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5010b, value : 32'h23038302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5010c, value : 32'he82c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5010d, value : 32'h22000006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5010e, value : 32'h23018302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5010f, value : 32'h20c082c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50110, value : 32'h70940066},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50111, value : 32'h2270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50112, value : 32'he0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50113, value : 32'h220e000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50114, value : 32'h25038142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50115, value : 32'h242f00c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50116, value : 32'he8100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50117, value : 32'h200e0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50118, value : 32'h25038140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50119, value : 32'h7ee00041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5011a, value : 32'h41404020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5011b, value : 32'h706c4260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5011c, value : 32'h20a8f1cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5011d, value : 32'h20000380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5011e, value : 32'h21018000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5011f, value : 32'h22018041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50120, value : 32'h72918082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50121, value : 32'h30622c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50122, value : 32'h6620c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50123, value : 32'h704cf1db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50124, value : 32'h706c6a09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50125, value : 32'h2212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50126, value : 32'h78e0f1e7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50127, value : 32'h81422253},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50128, value : 32'h224e7ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50129, value : 32'h168803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5012a, value : 32'h2801000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5012b, value : 32'h290000cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5012c, value : 32'h28000081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5012d, value : 32'h7fe00080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5012e, value : 32'h234e7985},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5012f, value : 32'h28000003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50130, value : 32'h7fe000c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50131, value : 32'h78e07802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50132, value : 32'h81422253},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50133, value : 32'h224e7ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50134, value : 32'h168803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50135, value : 32'h2900000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50136, value : 32'h290100cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50137, value : 32'h28010081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50138, value : 32'h7fe00080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50139, value : 32'h234e7885},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5013a, value : 32'h29010003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5013b, value : 32'h7fe000c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5013c, value : 32'h78e07922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5013d, value : 32'h402069},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5013e, value : 32'hf1fe78e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5013f, value : 32'h20001d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50140, value : 32'h78e0700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50141, value : 32'h87c82941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50142, value : 32'h2221ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50143, value : 32'h87c32842},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50144, value : 32'h2220ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50145, value : 32'h10c82007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50146, value : 32'h8040220a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50147, value : 32'h210050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50148, value : 32'h700c4100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50149, value : 32'h2d2f6869},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5014a, value : 32'h25ca8041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5014b, value : 32'h2e2f00c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5014c, value : 32'h26ca8081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5014d, value : 32'h260200c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5014e, value : 32'h23ca8143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5014f, value : 32'h23400024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50150, value : 32'h2ac0007c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50151, value : 32'h20a800c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50152, value : 32'h210202c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50153, value : 32'h20cf8081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50154, value : 32'h21c00f06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50155, value : 32'h222f0085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50156, value : 32'h202f0082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50157, value : 32'h202f9202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50158, value : 32'h20ce0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50159, value : 32'h7fe00025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5015a, value : 32'h2221ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5015b, value : 32'hf802020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5015c, value : 32'h5740000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5015d, value : 32'hf000260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5015e, value : 32'hfbf208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5015f, value : 32'h6420ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50160, value : 32'h202f7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50161, value : 32'h7fe00003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50162, value : 32'h78e0770c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50163, value : 32'h704c702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50164, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50165, value : 32'h70cc70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50166, value : 32'h700d70ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50167, value : 32'h704d702d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50168, value : 32'h708d706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50169, value : 32'h70cd70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5016a, value : 32'h700e70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5016b, value : 32'h704e702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5016c, value : 32'h708e706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5016d, value : 32'h70ce70ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5016e, value : 32'h700f70ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5016f, value : 32'h706f702f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50170, value : 32'h3000254a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50171, value : 32'h3000264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50172, value : 32'h800144db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50173, value : 32'h42db8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50174, value : 32'h4008000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50175, value : 32'hffcf0ab6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50176, value : 32'h54009aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50177, value : 32'h719d830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50178, value : 32'hf1feffcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50179, value : 32'hc1ec0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5017a, value : 32'hc1a1ffcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5017b, value : 32'h7487e805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5017c, value : 32'h7fe0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5017d, value : 32'h40c3c0a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5017e, value : 32'h12298000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5017f, value : 32'h206f8840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50180, value : 32'ha84007c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50181, value : 32'h208c8803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50182, value : 32'hf20d8fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50183, value : 32'hc040c084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50184, value : 32'h9124020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50185, value : 32'hc1840960},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50186, value : 32'hd8ffd911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50187, value : 32'h26008ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50188, value : 32'hfbab911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50189, value : 32'hd8ff0920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5018a, value : 32'h20ab700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5018b, value : 32'h7fff00c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5018c, value : 32'h78e0f1ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5018d, value : 32'h47cbc2f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5018e, value : 32'h11e28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5018f, value : 32'h10951746},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50190, value : 32'h23784310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50191, value : 32'h40580000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50192, value : 32'h4130781b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50193, value : 32'h2040704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50194, value : 32'h23140057},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50195, value : 32'h19002556},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50196, value : 32'h252f0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50197, value : 32'hfaf1487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50198, value : 32'h72b52364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50199, value : 32'h2fc1208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5019a, value : 32'h20542244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5019b, value : 32'h352e089b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5019c, value : 32'h202620ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5019d, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5019e, value : 32'h1b8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5019f, value : 32'h800146cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a0, value : 32'h8214d6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a1, value : 32'h40c3009e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a2, value : 32'h4868000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a3, value : 32'he88a8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a4, value : 32'h20300b1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a5, value : 32'h88e7eb4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a6, value : 32'h961200e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a7, value : 32'hf00d961e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a8, value : 32'he00882},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501a9, value : 32'h134026f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501aa, value : 32'h96067eb4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ab, value : 32'h876f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ac, value : 32'h960c00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ad, value : 32'h87e9618},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ae, value : 32'h700c00c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501af, value : 32'ha00bfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b0, value : 32'h2c40712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b1, value : 32'h70ad20ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b2, value : 32'h23c02632},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b3, value : 32'h10250d3b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b4, value : 32'h21002d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b5, value : 32'h4c02016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b6, value : 32'he02460b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b7, value : 32'h294060e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b8, value : 32'h20050380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501b9, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ba, value : 32'h90000234},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501bb, value : 32'h260090e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501bc, value : 32'hb8c6b8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501bd, value : 32'h200771a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501be, value : 32'h40260401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501bf, value : 32'h782579d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c0, value : 32'h20001900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c1, value : 32'h7146f1e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c2, value : 32'hc6d8f1a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c3, value : 32'hc1b4c3f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c4, value : 32'h16004110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c5, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c6, value : 32'h4750000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c7, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c8, value : 32'h81b11e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501c9, value : 32'h4728003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ca, value : 32'hf483b8e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501cb, value : 32'h41e14022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501cc, value : 32'hf0642e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501cd, value : 32'h4380ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ce, value : 32'h1f00c7d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501cf, value : 32'hc0801001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d0, value : 32'h10951646},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d1, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d2, value : 32'hda4e0f1a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d3, value : 32'hffef099a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d4, value : 32'h700c708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d5, value : 32'h704c702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d6, value : 32'h4200f46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d7, value : 32'h42c3706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d8, value : 32'hffff0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501d9, value : 32'h722c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501da, value : 32'h44404340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501db, value : 32'h4200eaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501dc, value : 32'hc0804540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501dd, value : 32'h9a00b56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501de, value : 32'h2114d94e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501df, value : 32'h43d32552},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e0, value : 32'hf8049007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e1, value : 32'h21051b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e2, value : 32'h208a7296},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e3, value : 32'h24442fc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e4, value : 32'hf8b2056},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e5, value : 32'h20ca25ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e6, value : 32'h45cb2026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e7, value : 32'h4d6c8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e8, value : 32'h7400c06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501e9, value : 32'ha00f7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ea, value : 32'h150025f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501eb, value : 32'h15002514},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ec, value : 32'ha00f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ed, value : 32'h218a9006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ee, value : 32'h40c30fcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ef, value : 32'hc2ec9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f0, value : 32'h712cb020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f1, value : 32'h51800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f2, value : 32'haf2700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f3, value : 32'h70ad00a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f4, value : 32'h23802232},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f5, value : 32'h2e40e823},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f6, value : 32'h2d4020d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f7, value : 32'h20162100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f8, value : 32'h60b80440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501f9, value : 32'h60c9e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501fa, value : 32'h3802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501fb, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501fc, value : 32'h26fc9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501fd, value : 32'h208a9040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501fe, value : 32'h8020fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h501ff, value : 32'h78460260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50200, value : 32'h71a5b8c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50201, value : 32'h4002007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50202, value : 32'h5812800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50203, value : 32'h78258700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50204, value : 32'h2232a700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50205, value : 32'hdc72380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50206, value : 32'h71869004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50207, value : 32'ha1140c6d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50208, value : 32'h70051e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50209, value : 32'h4901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5020a, value : 32'h20051b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5020b, value : 32'h1f00c7d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5020c, value : 32'h708e1001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5020d, value : 32'h10931646},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5020e, value : 32'h24d22114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5020f, value : 32'h208a7296},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50210, value : 32'h24442fc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50211, value : 32'hf692055},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50212, value : 32'h20ca256e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50213, value : 32'h45cb2026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50214, value : 32'h4d6c8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50215, value : 32'h7400b52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50216, value : 32'ha00eca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50217, value : 32'h150025f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50218, value : 32'h150d2514},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50219, value : 32'ha00ece},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5021a, value : 32'h700c9506},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5021b, value : 32'ha00a4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5021c, value : 32'h2232712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5021d, value : 32'he81c2380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5021e, value : 32'h20d52d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5021f, value : 32'h2b4070ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50220, value : 32'h41222100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50221, value : 32'h4402016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50222, value : 32'he02460b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50223, value : 32'h7200a02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50224, value : 32'hb8c660c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50225, value : 32'h200771a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50226, value : 32'h28000400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50227, value : 32'h87000541},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50228, value : 32'ha7007825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50229, value : 32'h23802232},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5022a, value : 32'h90040dd7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5022b, value : 32'hc917186},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5022c, value : 32'hf144a114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5022d, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5022e, value : 32'h2494b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5022f, value : 32'h710c3923},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50230, value : 32'hfdf218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50231, value : 32'h5200c2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50232, value : 32'hc809704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50233, value : 32'h3643236f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50234, value : 32'h685270ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50235, value : 32'hf802205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50236, value : 32'h949004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50237, value : 32'hc0449000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50238, value : 32'h30801300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50239, value : 32'h80be2053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5023a, value : 32'hc004f20b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5023b, value : 32'hf812205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5023c, value : 32'hc0949007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5023d, value : 32'h80206c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5023e, value : 32'hc02045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5023f, value : 32'h2205b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50240, value : 32'h90080f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50241, value : 32'h9040002c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50242, value : 32'h2443276f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50243, value : 32'h17004040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50244, value : 32'h20842081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50245, value : 32'h217800cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50246, value : 32'h20b80103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50247, value : 32'h41c30084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50248, value : 32'h20192},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50249, value : 32'h40c37b04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5024a, value : 32'h12e28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5024b, value : 32'hddaa860},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5024c, value : 32'h740c0220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5024d, value : 32'hc08eda07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5024e, value : 32'hfc6ba09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5024f, value : 32'h702cffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50250, value : 32'ha08017f9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50251, value : 32'h19341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50252, value : 32'h20440000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50253, value : 32'h1c0c0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50254, value : 32'h20783344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50255, value : 32'hc5420000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50256, value : 32'hc540c541},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50257, value : 32'hffef0c8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50258, value : 32'h1713c54b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50259, value : 32'h47cb2081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5025a, value : 32'h4848000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5025b, value : 32'h1002941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5025c, value : 32'hdf0815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5025d, value : 32'h9f0819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5025e, value : 32'h7f081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5025f, value : 32'h1f00710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50260, value : 32'hf00d1043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50261, value : 32'h1f00d808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50262, value : 32'hf0091203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50263, value : 32'h1f00740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50264, value : 32'hf0051103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50265, value : 32'h1f00720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50266, value : 32'hb9e21083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50267, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50268, value : 32'h20ca0f14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50269, value : 32'h764c0062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5026a, value : 32'hf3eaf01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5026b, value : 32'hc08cffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5026c, value : 32'h712cc08c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5026d, value : 32'h7a00946},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5026e, value : 32'hb4e714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5026f, value : 32'hc08003a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50270, value : 32'h4c00d76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50271, value : 32'h46cb700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50272, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50273, value : 32'h30031c17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50274, value : 32'h408202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50275, value : 32'h2440c187},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50276, value : 32'h83a3ac2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50277, value : 32'h244003e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50278, value : 32'h8c535c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50279, value : 32'h40c30011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5027a, value : 32'h11408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5027b, value : 32'h431800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5027c, value : 32'h30801417},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5027d, value : 32'h2a00e92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5027e, value : 32'hb4a4210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5027f, value : 32'h142b0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50280, value : 32'h17133091},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50281, value : 32'hb8e22080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50282, value : 32'h1f024022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50283, value : 32'hf42b1003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50284, value : 32'hcca712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50285, value : 32'hc28e07e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50286, value : 32'hc18b8e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50287, value : 32'h3093141c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50288, value : 32'h19845cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50289, value : 32'h23140002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5028a, value : 32'h61792083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5028b, value : 32'ha9004362},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5028c, value : 32'hcd6740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5028d, value : 32'h41a10220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5028e, value : 32'hc3e4042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5028f, value : 32'hc18e0260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50290, value : 32'h702c4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50291, value : 32'h7e00c96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50292, value : 32'h8e40c28e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50293, value : 32'h1401254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50294, value : 32'hcb6740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50295, value : 32'h43620220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50296, value : 32'hc1e4042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50297, value : 32'hc18e0260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50298, value : 32'hc18ef022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50299, value : 32'h706c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5029a, value : 32'hfc1248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5029b, value : 32'h200c7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5029c, value : 32'h8e2070ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5029d, value : 32'h2514c527},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5029e, value : 32'hc18b1042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5029f, value : 32'ha9006159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a0, value : 32'hdf64022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a1, value : 32'hc18e0360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a2, value : 32'h740c8e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a3, value : 32'h19641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a4, value : 32'hc760002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a5, value : 32'h43a10220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a6, value : 32'hbde4042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a7, value : 32'hc18e0260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a8, value : 32'h10431f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502a9, value : 32'h202f7106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502aa, value : 32'h8290408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ab, value : 32'hc8098114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ac, value : 32'hdd07708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ad, value : 32'h20057885},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ae, value : 32'h30f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502af, value : 32'he72f0d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b0, value : 32'h702c0920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b1, value : 32'h258dc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b2, value : 32'h24561e3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b3, value : 32'hb802180c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b4, value : 32'h2005700f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b5, value : 32'h900f0f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b6, value : 32'hc1ec364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b7, value : 32'h180006e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b8, value : 32'h14170604},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502b9, value : 32'h44d33080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ba, value : 32'h1668000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502bb, value : 32'h30192440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502bc, value : 32'h1c00700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502bd, value : 32'h1cff2fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502be, value : 32'hc046afc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502bf, value : 32'h200cc006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c0, value : 32'h292a000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c1, value : 32'hd9d30026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c2, value : 32'h20801713},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c3, value : 32'hff0821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c4, value : 32'h876d840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c5, value : 32'h43000780},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c6, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c7, value : 32'h2019b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c8, value : 32'h2200be6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502c9, value : 32'h228a4202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ca, value : 32'hf00e2001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502cb, value : 32'h7a0085a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502cc, value : 32'h4300700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502cd, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ce, value : 32'h2019a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502cf, value : 32'h2200bca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d0, value : 32'h704e4202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d1, value : 32'h28152255},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d2, value : 32'h2480260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d3, value : 32'h203e2680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d4, value : 32'h7676706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d5, value : 32'h2d013a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d6, value : 32'h2fc3218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d7, value : 32'h70ad70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d8, value : 32'h708d706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502d9, value : 32'hc18e4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502da, value : 32'h1c209a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502db, value : 32'h61197ad0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502dc, value : 32'h22002b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502dd, value : 32'h60496038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502de, value : 32'h448202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502df, value : 32'h8fc3208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e0, value : 32'h7034f408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e1, value : 32'hd8ff41a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e2, value : 32'h41d170ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e3, value : 32'hf02bf429},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e4, value : 32'h228ce924},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e5, value : 32'h3e8042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e6, value : 32'h7ab00025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e7, value : 32'h9377970},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e8, value : 32'hfe60085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502e9, value : 32'h43000740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ea, value : 32'hfde6e09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502eb, value : 32'h78100760},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ec, value : 32'h8f014400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ed, value : 32'hfd260b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ee, value : 32'h78100760},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ef, value : 32'h740c4500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f0, value : 32'h19d41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f1, value : 32'hb420004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f2, value : 32'h42620220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f3, value : 32'h442a8f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f4, value : 32'h41a1651b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f5, value : 32'hf005d8ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f6, value : 32'h40228f21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f7, value : 32'h452861b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f8, value : 32'h8f014110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502f9, value : 32'h79d0661e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502fa, value : 32'h8004218c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502fb, value : 32'hffc50778},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502fc, value : 32'h262f7970},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502fd, value : 32'h2179f348},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502fe, value : 32'h651d0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h502ff, value : 32'h6121c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50300, value : 32'h3082120b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50301, value : 32'h80412144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50302, value : 32'h78b0757c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50303, value : 32'ha5081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50304, value : 32'h41c3d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50305, value : 32'h101a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50306, value : 32'h2000aee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50307, value : 32'h702c7bae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50308, value : 32'h832b44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50309, value : 32'hf01f710f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5030a, value : 32'h70347bae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5030b, value : 32'h832b44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5030c, value : 32'h144124ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5030d, value : 32'h23002600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5030e, value : 32'h262f6078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5030f, value : 32'h16f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50310, value : 32'h704c0024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50311, value : 32'hd137910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50312, value : 32'h25022065},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50313, value : 32'h42a22001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50314, value : 32'h4100f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50315, value : 32'h702cf003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50316, value : 32'hc0874200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50317, value : 32'h4c02014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50318, value : 32'h6179b040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50319, value : 32'h2048782e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5031a, value : 32'h8170000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5031b, value : 32'h780f2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5031c, value : 32'h20811400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5031d, value : 32'h402009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5031e, value : 32'h20021c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5031f, value : 32'h14fff007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50320, value : 32'h2009a081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50321, value : 32'h1cff0040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50322, value : 32'h7166a002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50323, value : 32'h2840f163},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50324, value : 32'h2440230d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50325, value : 32'hde073713},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50326, value : 32'h2640250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50327, value : 32'h25001302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50328, value : 32'h24831501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50329, value : 32'h7600ee2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5032a, value : 32'h44004610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5032b, value : 32'h7600eda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5032c, value : 32'h45004042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5032d, value : 32'h4202750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5032e, value : 32'h1a241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5032f, value : 32'ha4a0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50330, value : 32'h41700220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50331, value : 32'h22012940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50332, value : 32'h79a5c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50333, value : 32'h20057825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50334, value : 32'h30f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50335, value : 32'hc5a00d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50336, value : 32'h41c20920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50337, value : 32'h183f268d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50338, value : 32'h3b112440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50339, value : 32'h24112114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5033a, value : 32'h20c01100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5033b, value : 32'h20487042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5033c, value : 32'h7e100000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5033d, value : 32'h7600e92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5033e, value : 32'h430040c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5033f, value : 32'h7600e8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50340, value : 32'h44004042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50341, value : 32'h41c3750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50342, value : 32'h301a3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50343, value : 32'h22009fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50344, value : 32'hc8094202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50345, value : 32'h200578a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50346, value : 32'h30f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50347, value : 32'hc1208d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50348, value : 32'h41c10920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50349, value : 32'h20c01101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5034a, value : 32'h20487042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5034b, value : 32'h7e100000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5034c, value : 32'h7600e56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5034d, value : 32'h430040c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5034e, value : 32'h7600e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5034f, value : 32'h44004042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50350, value : 32'h41c3750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50351, value : 32'h301a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50352, value : 32'h22009be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50353, value : 32'hc8094202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50354, value : 32'h200578a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50355, value : 32'h30f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50356, value : 32'hbd609d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50357, value : 32'h41c10920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50358, value : 32'h7600e26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50359, value : 32'h43004042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5035a, value : 32'h41c3750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5035b, value : 32'h201a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5035c, value : 32'h2200996},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5035d, value : 32'hc8094202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5035e, value : 32'h200578a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5035f, value : 32'h30f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50360, value : 32'hbae00d9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50361, value : 32'h41420920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50362, value : 32'h31d92140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50363, value : 32'hffef0571},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50364, value : 32'h20787106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50365, value : 32'h8523000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50366, value : 32'hb911ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50367, value : 32'h6c0095a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50368, value : 32'h7000e06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50369, value : 32'h20801713},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5036a, value : 32'h3e0815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5036b, value : 32'hb88d700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5036c, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5036d, value : 32'h148000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5036e, value : 32'h5000a22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5036f, value : 32'h30801300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50370, value : 32'h80be2053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50371, value : 32'hde2f20b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50372, value : 32'hc8090700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50373, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50374, value : 32'h90070f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50375, value : 32'hc004c094},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50376, value : 32'hc08cb100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50377, value : 32'hd1e712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50378, value : 32'h704c0760},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50379, value : 32'h702c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5037a, value : 32'h4e00f0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5037b, value : 32'h2494704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5037c, value : 32'h1404371c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5037d, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5037e, value : 32'h47cbc2f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5037f, value : 32'h11e28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50380, value : 32'h10921746},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50381, value : 32'h46304550},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50382, value : 32'h7200d9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50383, value : 32'h40c24410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50384, value : 32'h428241a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50385, value : 32'h9600c7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50386, value : 32'h40c3706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50387, value : 32'h27100000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50388, value : 32'h5a00972},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50389, value : 32'h2453702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5038a, value : 32'h702e2040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5038b, value : 32'h902078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5038c, value : 32'h201470cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5038d, value : 32'h70ad2493},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5038e, value : 32'h23c02332},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5038f, value : 32'h10250d4b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50390, value : 32'h21002a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50391, value : 32'h4002016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50392, value : 32'he02460b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50393, value : 32'h160060e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50394, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50395, value : 32'h2053000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50396, value : 32'hf20780be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50397, value : 32'hc324020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50398, value : 32'h410206e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50399, value : 32'h2940f00b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5039a, value : 32'h20050380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5039b, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5039c, value : 32'h90000234},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5039d, value : 32'h2200986},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5039e, value : 32'h2053b8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5039f, value : 32'h71a581be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a0, value : 32'h106226c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a1, value : 32'hd22f1da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a2, value : 32'h40c20700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a3, value : 32'h428241a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a4, value : 32'h9600bfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a5, value : 32'h2332db7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a6, value : 32'h94d23c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a7, value : 32'h2a402025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a8, value : 32'h20162100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503a9, value : 32'h70220400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503aa, value : 32'h60e9e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ab, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ac, value : 32'hc8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ad, value : 32'h80be2053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ae, value : 32'h4020f206},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503af, value : 32'h6e00bd2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b0, value : 32'hf00c4102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b1, value : 32'h3802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b2, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b3, value : 32'h2349004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b4, value : 32'h92a9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b5, value : 32'hb8c80220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b6, value : 32'h7126b8c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b7, value : 32'hfc120b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b8, value : 32'hf1db7e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503b9, value : 32'hc6d478cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ba, value : 32'hc1a1c3fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503bb, value : 32'hd8404210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503bc, value : 32'h210ab89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503bd, value : 32'h250a3140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503be, value : 32'h47682100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503bf, value : 32'h901000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c0, value : 32'h10e54350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c1, value : 32'h46308097},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c2, value : 32'h800041d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c3, value : 32'hea081140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c4, value : 32'hb764042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c5, value : 32'h712c02a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c6, value : 32'h20031900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c7, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c8, value : 32'h1b8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503c9, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ca, value : 32'h8291228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503cb, value : 32'h708e007e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503cc, value : 32'h20300b21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503cd, value : 32'he524042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ce, value : 32'h8d400480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503cf, value : 32'h750c4410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d0, value : 32'h18941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d1, value : 32'h43420003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d2, value : 32'h1e00fbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d3, value : 32'h500240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d4, value : 32'h740c8d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d5, value : 32'h41c34342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d6, value : 32'h5018c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d7, value : 32'h4c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d8, value : 32'h260a45e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503d9, value : 32'hfa20540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503da, value : 32'h225301e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503db, value : 32'h46cb2058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503dc, value : 32'h4878000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503dd, value : 32'he8128e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503de, value : 32'h201f0f09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503df, value : 32'h201e080b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e0, value : 32'h4200aa6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e1, value : 32'hf0b710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e2, value : 32'h80d205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e3, value : 32'ha9a205e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e4, value : 32'h720c0420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e5, value : 32'h10031e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e6, value : 32'h41c37156},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e7, value : 32'h8d80003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e8, value : 32'h2078c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503e9, value : 32'h21d63097},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ea, value : 32'h78250822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503eb, value : 32'hb90c8d20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ec, value : 32'h97e7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ed, value : 32'hd9400920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ee, value : 32'h710e7076},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ef, value : 32'h24a220ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f0, value : 32'hd937ef0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f1, value : 32'h740c23a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f2, value : 32'h234a708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f3, value : 32'hc80911c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f4, value : 32'h3012005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f5, value : 32'hb80c8d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f6, value : 32'h20057825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f7, value : 32'h30f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f8, value : 32'h94e00d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503f9, value : 32'h41c10920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503fa, value : 32'h1cff238d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503fb, value : 32'h180c2456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503fc, value : 32'h6800f06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503fd, value : 32'hc18040e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503fe, value : 32'h716c734c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h503ff, value : 32'hffaf0f12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50400, value : 32'hc400718c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50401, value : 32'h71c0244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50402, value : 32'h20a8706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50403, value : 32'h2c0108c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50404, value : 32'h2b4012c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50405, value : 32'h20441202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50406, value : 32'h8d000043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50407, value : 32'h1c209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50408, value : 32'h605870c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50409, value : 32'h882060d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5040a, value : 32'ha8207965},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5040b, value : 32'h12002340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5040c, value : 32'h10002c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5040d, value : 32'h20447165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5040e, value : 32'h8d000041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5040f, value : 32'h1c209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50410, value : 32'h621a70c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50411, value : 32'h10806658},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50412, value : 32'h79450282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50413, value : 32'h7702a820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50414, value : 32'h8d40f1b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50415, value : 32'h41c34342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50416, value : 32'h3018e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50417, value : 32'h1e00eaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50418, value : 32'h4c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50419, value : 32'hdc0770ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5041a, value : 32'h78a5c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5041b, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5041c, value : 32'hf0d80003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5041d, value : 32'h92008ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5041e, value : 32'h248d702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5041f, value : 32'h25561e3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50420, value : 32'he76180d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50421, value : 32'h9170680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50422, value : 32'hb133010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50423, value : 32'h40422031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50424, value : 32'hc86702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50425, value : 32'h190002e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50426, value : 32'h40822043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50427, value : 32'h78e0c7da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50428, value : 32'h41c3c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50429, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5042a, value : 32'h89208941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5042b, value : 32'h2c1229f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5042c, value : 32'h582219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5042d, value : 32'h621a6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5042e, value : 32'hb8c38a02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5042f, value : 32'h2009d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50430, value : 32'h68d205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50431, value : 32'h802079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50432, value : 32'h186209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50433, value : 32'h2534651d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50434, value : 32'h80001f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50435, value : 32'hc6c20a84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50436, value : 32'h962c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50437, value : 32'h716c0100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50438, value : 32'hda62e89d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50439, value : 32'h800140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5043a, value : 32'hba9f4e7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5043b, value : 32'h8a208800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5043c, value : 32'h262f7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5043d, value : 32'h26f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5043e, value : 32'h12340004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5043f, value : 32'h208b0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50440, value : 32'hf40d8401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50441, value : 32'h10008ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50442, value : 32'h916e889},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50443, value : 32'he8870100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50444, value : 32'h801230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50445, value : 32'h4032044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50446, value : 32'hc0d1bb24},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50447, value : 32'h40607fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50448, value : 32'h4508c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50449, value : 32'hd8fa4110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5044a, value : 32'h46284748},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5044b, value : 32'h4e00e96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5044c, value : 32'h22c1219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5044d, value : 32'h20096a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5044e, value : 32'h40c34010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5044f, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50450, value : 32'h762c8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50451, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50452, value : 32'h244ada22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50453, value : 32'h70cc0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50454, value : 32'h20327022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50455, value : 32'h80010f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50456, value : 32'h710c4e8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50457, value : 32'hb80278b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50458, value : 32'h340200f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50459, value : 32'h7d0fbb86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5045a, value : 32'h97a700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5045b, value : 32'h45a10060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5045c, value : 32'h402202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5045d, value : 32'hf33e008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5045e, value : 32'h202f103e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5045f, value : 32'h700c2007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50460, value : 32'h724cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50461, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50462, value : 32'h95a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50463, value : 32'h260a0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50464, value : 32'h700c0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50465, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50466, value : 32'h244a43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50467, value : 32'h45a10380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50468, value : 32'h600942},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50469, value : 32'hf2f70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5046a, value : 32'h700c107e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5046b, value : 32'h724cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5046c, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5046d, value : 32'h92e70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5046e, value : 32'h260a0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5046f, value : 32'h700c0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50470, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50471, value : 32'h244a43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50472, value : 32'h45a103c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50473, value : 32'h600916},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50474, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50475, value : 32'h724cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50476, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50477, value : 32'h90670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50478, value : 32'h260a0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50479, value : 32'h700c0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5047a, value : 32'h724cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5047b, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5047c, value : 32'h8f270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5047d, value : 32'h264a0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5047e, value : 32'h700c0a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5047f, value : 32'h600896},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50480, value : 32'hc6ca712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50481, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50482, value : 32'h7fe0046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50483, value : 32'h51800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50484, value : 32'h1e00700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50485, value : 32'h901c7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50486, value : 32'h7ee00480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50487, value : 32'he08e4100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50488, value : 32'hf707710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50489, value : 32'h704e0e0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5048a, value : 32'h40410000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5048b, value : 32'he1a87ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5048c, value : 32'h7fe07ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5048d, value : 32'h78e0700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5048e, value : 32'h45cbc2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5048f, value : 32'h1a188000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50490, value : 32'he8049511},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50491, value : 32'h10451d28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50492, value : 32'h200872},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50493, value : 32'h460840a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50494, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50495, value : 32'hb0c0046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50496, value : 32'h702c40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50497, value : 32'hff6f0ea2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50498, value : 32'h700cda20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50499, value : 32'hb513b514},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5049a, value : 32'hb511b512},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5049b, value : 32'hc6c440c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5049c, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5049d, value : 32'h9103046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5049e, value : 32'h71109120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5049f, value : 32'h7ce0700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a0, value : 32'hffcf07b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a1, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a2, value : 32'h9000046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a3, value : 32'hb8227fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a4, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a5, value : 32'h7fe00476},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a6, value : 32'h78e08800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a7, value : 32'hc86c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a8, value : 32'h700c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504a9, value : 32'h600c8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504aa, value : 32'hada700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ab, value : 32'h700c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ac, value : 32'hffcf0f56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ad, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ae, value : 32'hc1a4c3f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504af, value : 32'h800043c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b0, value : 32'h8b28046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b1, value : 32'he90770cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b2, value : 32'h71c56949},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b3, value : 32'h80812104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b4, value : 32'h904ff5fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b5, value : 32'h100e8ba3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b6, value : 32'hb0b30115},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b7, value : 32'h1171004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b8, value : 32'h1161002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504b9, value : 32'h1028bd0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ba, value : 32'h1000010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504bb, value : 32'h10240109},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504bc, value : 32'h10120108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504bd, value : 32'h10140107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504be, value : 32'h2b400106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504bf, value : 32'h101012cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c0, value : 32'h90910104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c1, value : 32'h1051020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c2, value : 32'h11e100a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c3, value : 32'h11f1006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c4, value : 32'h1101008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c5, value : 32'h1131016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c6, value : 32'h111101a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c7, value : 32'h114100c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c8, value : 32'h1121018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504c9, value : 32'h226d902e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ca, value : 32'h1c0c0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504cb, value : 32'hb9c33004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504cc, value : 32'hda7f6a14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504cd, value : 32'h24537825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ce, value : 32'h1c0a20c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504cf, value : 32'h256d3004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d0, value : 32'h1c042300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d1, value : 32'h2d403004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d2, value : 32'h78252100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d3, value : 32'h1c02ba07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d4, value : 32'h2a403004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d5, value : 32'h235321c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d6, value : 32'h78442181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d7, value : 32'h29407905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d8, value : 32'h78252380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504d9, value : 32'h31812753},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504da, value : 32'h30041c08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504db, value : 32'h21c02840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504dc, value : 32'h93e37844},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504dd, value : 32'h2e407905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504de, value : 32'h78253380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504df, value : 32'h2012d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e0, value : 32'h30041c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e1, value : 32'h21846c17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e2, value : 32'h2004000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e3, value : 32'hf80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e4, value : 32'h78257c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e5, value : 32'h1012c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e6, value : 32'h4012144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e7, value : 32'h7905bc0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e8, value : 32'h1402f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504e9, value : 32'h8012084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ea, value : 32'h79058b4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504eb, value : 32'h1c02e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ec, value : 32'h7825780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ed, value : 32'h12012840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ee, value : 32'h30041c0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ef, value : 32'h1f802404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f0, value : 32'h70000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f1, value : 32'hc2184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f2, value : 32'h782578a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f3, value : 32'h1f812304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f4, value : 32'h8000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f5, value : 32'h29407825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f6, value : 32'h21441101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f7, value : 32'h79050401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f8, value : 32'h21402e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504f9, value : 32'h8012084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504fa, value : 32'h2f407905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504fb, value : 32'h780f21c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504fc, value : 32'h79fd7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504fd, value : 32'h30041c06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504fe, value : 32'ha6dea08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h504ff, value : 32'h7ccf0071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50500, value : 32'h641c8b09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50501, value : 32'h12140c57},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50502, value : 32'h244a6912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50503, value : 32'h20057100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50504, value : 32'h100f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50505, value : 32'hc0804000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50506, value : 32'h3c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50507, value : 32'h50b1002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50508, value : 32'hf8d2105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50509, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5050a, value : 32'h50c1002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5050b, value : 32'hbc107424},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5050c, value : 32'h12cc2405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5050d, value : 32'h4f98a580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5050e, value : 32'h907e2053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5050f, value : 32'hb323b9a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50510, value : 32'h710cf205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50511, value : 32'h2002006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50512, value : 32'h40c3ab0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50513, value : 32'h1a388000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50514, value : 32'h710a15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50515, value : 32'h51800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50516, value : 32'h60d88b09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50517, value : 32'h31b08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50518, value : 32'hab09b8c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50519, value : 32'hc7d67830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5051a, value : 32'h4350c2ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5051b, value : 32'h9d74130},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5051c, value : 32'h47080030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5051d, value : 32'h2fc3208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5051e, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5051f, value : 32'h70cd1a18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50520, value : 32'h2448222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50521, value : 32'h21140a1d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50522, value : 32'h20300b19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50523, value : 32'h90be2753},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50524, value : 32'h700cf219},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50525, value : 32'ha5077726},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50526, value : 32'ha505a506},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50527, value : 32'hf02ea504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50528, value : 32'h90be2753},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50529, value : 32'ha69f21f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5052a, value : 32'h74e52070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5052b, value : 32'ha5c6a5c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5052c, value : 32'hd8aa5c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5052d, value : 32'ha5c4ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5052e, value : 32'h20b00a49},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5052f, value : 32'h77264708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50530, value : 32'h40a1f1e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50531, value : 32'hc3a702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50532, value : 32'hda20ff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50533, value : 32'ha048228c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50534, value : 32'h250046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50535, value : 32'h1d22732c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50536, value : 32'h21801404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50537, value : 32'hb5322038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50538, value : 32'ha21f00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50539, value : 32'h40a12070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5053a, value : 32'hc16702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5053b, value : 32'hda20ff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5053c, value : 32'h20b00a3b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5053d, value : 32'h20912142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5053e, value : 32'hffcf0d42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5053f, value : 32'hf1c24708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50540, value : 32'h74e5a5c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50541, value : 32'ha5c1a5c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50542, value : 32'hf01da5c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50543, value : 32'ha5c6a5c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50544, value : 32'ha5c4a5c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50545, value : 32'h2104f017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50546, value : 32'h2f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50547, value : 32'h781dfffe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50548, value : 32'h203f090f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50549, value : 32'hb5327704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5054a, value : 32'he708b511},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5054b, value : 32'hb532f00b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5054c, value : 32'hffef0d0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5054d, value : 32'h702cb511},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5054e, value : 32'ha52068e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5054f, value : 32'ha522a521},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50550, value : 32'h78f0a523},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50551, value : 32'h78e0c6ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50552, value : 32'h4508c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50553, value : 32'h600836},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50554, value : 32'h80c208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50555, value : 32'h752cd809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50556, value : 32'hda0cb813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50557, value : 32'h8238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50558, value : 32'h45a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50559, value : 32'h200d7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5055a, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5055b, value : 32'h724c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5055c, value : 32'h244a736c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5055d, value : 32'h45a10680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5055e, value : 32'h200d6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5055f, value : 32'hb3270cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50560, value : 32'h700c03c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50561, value : 32'h724c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50562, value : 32'h244a716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50563, value : 32'h45a10680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50564, value : 32'h200d52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50565, value : 32'hb1a70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50566, value : 32'h700c03c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50567, value : 32'h724c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50568, value : 32'h244a706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50569, value : 32'h45a10680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5056a, value : 32'h200d3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5056b, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5056c, value : 32'h826d922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5056d, value : 32'h704c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5056e, value : 32'h752c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5056f, value : 32'h238a744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50570, value : 32'h708c000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50571, value : 32'hd1e45a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50572, value : 32'h70cc0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50573, value : 32'hd907d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50574, value : 32'h744cb893},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50575, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50576, value : 32'hd0a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50577, value : 32'h70cc0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50578, value : 32'hffcf0ca6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50579, value : 32'h78107704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5057a, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5057b, value : 32'h40c3c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5057c, value : 32'h61a80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5057d, value : 32'h80e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5057e, value : 32'hffcf0c1a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5057f, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50580, value : 32'h72081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50581, value : 32'h1600714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50582, value : 32'h901c7101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50583, value : 32'he9850484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50584, value : 32'h71447210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50585, value : 32'h2179f6b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50586, value : 32'hf0030000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50587, value : 32'hd90b700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50588, value : 32'hff6f07c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50589, value : 32'h78e0b912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5058a, value : 32'h82dc2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5058b, value : 32'h43200072},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5058c, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5058d, value : 32'h8d42046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5058e, value : 32'h28057810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5058f, value : 32'hb110081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50590, value : 32'h9500027f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50591, value : 32'hea848d4b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50592, value : 32'hf003714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50593, value : 32'he1e704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50594, value : 32'hb500ffcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50595, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50596, value : 32'h70adc0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50597, value : 32'hb0a2e2b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50598, value : 32'hb0a7b0a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50599, value : 32'h302b0a6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5059a, value : 32'hb0a0002d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5059b, value : 32'h24ad4468},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5059c, value : 32'h20241203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5059d, value : 32'hf50080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5059e, value : 32'h1090000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5059f, value : 32'h1310000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a0, value : 32'h15b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a1, value : 32'h1850000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a2, value : 32'h1a50000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a3, value : 32'h1b30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a4, value : 32'hb70000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a5, value : 32'hbb0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a6, value : 32'h2cf0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a7, value : 32'hbd0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a8, value : 32'h1ab0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505a9, value : 32'h1b30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505aa, value : 32'h2bf0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ab, value : 32'h1af0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ac, value : 32'h1c10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ad, value : 32'h1c70000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ae, value : 32'ha10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505af, value : 32'h2ab0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b0, value : 32'h2a70000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b1, value : 32'h2a30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b2, value : 32'h29f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b3, value : 32'h29b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b4, value : 32'h2970000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b5, value : 32'h2930000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b6, value : 32'h1ad0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b7, value : 32'h1bb0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b8, value : 32'h6f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505b9, value : 32'h1c10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ba, value : 32'h1e90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505bb, value : 32'h1e90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505bc, value : 32'h1eb0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505bd, value : 32'h6f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505be, value : 32'h17d0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505bf, value : 32'h1e90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c0, value : 32'h1e90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c1, value : 32'h1f10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c2, value : 32'h1f30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c3, value : 32'h570000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c4, value : 32'h370000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c5, value : 32'h1f30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c6, value : 32'h1f70000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c7, value : 32'h1f70000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c8, value : 32'h1f70000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505c9, value : 32'h1f90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ca, value : 32'h1f90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505cb, value : 32'h1fd0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505cc, value : 32'h20b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505cd, value : 32'h2210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ce, value : 32'hf0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505cf, value : 32'h21d0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d0, value : 32'h21d0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d1, value : 32'hb0a40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d2, value : 32'h20021f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d3, value : 32'hdb78b0a3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d4, value : 32'h2453b063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d5, value : 32'hf0a600c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d6, value : 32'hb063db38},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d7, value : 32'h832453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d8, value : 32'h203f0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505d9, value : 32'hbbc60020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505da, value : 32'h2f270d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505db, value : 32'h23530021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505dc, value : 32'hbb24018c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505dd, value : 32'he012384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505de, value : 32'h2345b084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505df, value : 32'hf0f400c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e0, value : 32'h2c406bf3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e1, value : 32'h2453008c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e2, value : 32'h274400c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e3, value : 32'h24841c0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e4, value : 32'h24051001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e5, value : 32'h24050384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e6, value : 32'h7b7d110c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e7, value : 32'h2344b084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e8, value : 32'h2744070c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505e9, value : 32'h7b851203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ea, value : 32'hf0debb80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505eb, value : 32'h2c406bd3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ec, value : 32'h2453008c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ed, value : 32'h264400c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ee, value : 32'h24841c0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ef, value : 32'h24051001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f0, value : 32'h240503c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f1, value : 32'h7b7d110c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f2, value : 32'h2644b084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f3, value : 32'h2344120c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f4, value : 32'h7b850603},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f5, value : 32'h1432345},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f6, value : 32'h6bd3f0c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f7, value : 32'h8c2c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f8, value : 32'hc42453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505f9, value : 32'h1c0f2644},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505fa, value : 32'h10012484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505fb, value : 32'h3c42405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505fc, value : 32'h110c2405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505fd, value : 32'hb0847b7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505fe, value : 32'h120c2644},
                          '{ step_type : REG_WRITE, reg_addr : 32'h505ff, value : 32'h6032344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50600, value : 32'h23457b85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50601, value : 32'hf0b00183},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50602, value : 32'hbb037c7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50603, value : 32'h160c2444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50604, value : 32'hc032344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50605, value : 32'hb083bc82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50606, value : 32'h8c2c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50607, value : 32'hc42453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50608, value : 32'h10012484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50609, value : 32'h1032305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5060a, value : 32'hf03c7b85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5060b, value : 32'h2453bb23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5060c, value : 32'h2384018c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5060d, value : 32'hb0840c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5060e, value : 32'h3032345},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5060f, value : 32'he25f094},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50610, value : 32'h2370011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50611, value : 32'h18080020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50612, value : 32'hbb050104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50613, value : 32'h2384dc68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50614, value : 32'hb0830801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50615, value : 32'hdb28f026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50616, value : 32'h70d4f060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50617, value : 32'h10218},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50618, value : 32'h18c2353},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50619, value : 32'h23847b7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5061a, value : 32'hb0840001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5061b, value : 32'hf07cbb83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5061c, value : 32'h1041808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5061d, value : 32'h6051806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5061e, value : 32'hdb38f077},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5061f, value : 32'h2453b063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50620, value : 32'hf00f0083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50621, value : 32'h18c2353},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50622, value : 32'h23847b7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50623, value : 32'hb0840001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50624, value : 32'hc032345},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50625, value : 32'hdb78f068},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50626, value : 32'h2453b063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50627, value : 32'hbb8600c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50628, value : 32'hf063b064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50629, value : 32'h2c406bd3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5062a, value : 32'h2453008c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5062b, value : 32'h264400c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5062c, value : 32'h24841c0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5062d, value : 32'h24051001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5062e, value : 32'h240503c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5062f, value : 32'h7b7d110c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50630, value : 32'h2644b084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50631, value : 32'h2344120c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50632, value : 32'h7b850703},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50633, value : 32'hf04cbb81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50634, value : 32'hf049db58},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50635, value : 32'hb083b084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50636, value : 32'h7b7df047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50637, value : 32'h12384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50638, value : 32'hf041bb83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50639, value : 32'hf041b084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5063a, value : 32'h2384bb23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5063b, value : 32'h23450c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5063c, value : 32'hf0390303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5063d, value : 32'h1832453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5063e, value : 32'h7b7df035},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5063f, value : 32'h12384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50640, value : 32'hc032345},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50641, value : 32'h70d4f02f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50642, value : 32'hdb40f51f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50643, value : 32'hdb60f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50644, value : 32'hdb20f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50645, value : 32'hdb50f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50646, value : 32'hf026b0a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50647, value : 32'hf023db38},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50648, value : 32'h832453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50649, value : 32'hf01fbb86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5064a, value : 32'hbb037c7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5064b, value : 32'h170c2444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5064c, value : 32'h2032344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5064d, value : 32'hbb807b85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5064e, value : 32'hbb03f015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5064f, value : 32'h8c2c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50650, value : 32'hc42453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50651, value : 32'hc032344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50652, value : 32'h10012484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50653, value : 32'h1032305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50654, value : 32'hf0097b85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50655, value : 32'hf007db40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50656, value : 32'hf005db68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50657, value : 32'h2384bb05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50658, value : 32'hb0640801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50659, value : 32'h91db063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5065a, value : 32'ha19041f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5065b, value : 32'h22780c70},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5065c, value : 32'h230b0a03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5065d, value : 32'hf4068180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5065e, value : 32'h432553},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5065f, value : 32'hf003b065},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50660, value : 32'h939b0a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50661, value : 32'hdb0d053f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50662, value : 32'h57f0937},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50663, value : 32'h939dbd0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50664, value : 32'hdb0d05bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50665, value : 32'h5ff0937},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50666, value : 32'h939db08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50667, value : 32'hdb80063f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50668, value : 32'h67f09b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50669, value : 32'h10238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5066a, value : 32'h6bf09d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5066b, value : 32'h4238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5066c, value : 32'h6ff09d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5066d, value : 32'hf010706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5066e, value : 32'h345180e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5066f, value : 32'hb067f00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50670, value : 32'hf00adbd0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50671, value : 32'hb067bb08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50672, value : 32'h180ef006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50673, value : 32'hf0040205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50674, value : 32'hdb80b067},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50675, value : 32'h909bb8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50676, value : 32'hb06704de},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50677, value : 32'h7550a13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50678, value : 32'h708f0e21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50679, value : 32'h181000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5067a, value : 32'hb21766c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5067b, value : 32'h2242008f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5067c, value : 32'hb190843},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5067d, value : 32'ha150094},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5067e, value : 32'he2a90af0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5067f, value : 32'hf414704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50680, value : 32'h180c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50681, value : 32'hf0100105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50682, value : 32'h832941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50683, value : 32'h7a66724c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50684, value : 32'h1032144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50685, value : 32'h21447074},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50686, value : 32'hb0d0303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50687, value : 32'h22cf0330},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50688, value : 32'hb0460021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50689, value : 32'h49e090b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5068a, value : 32'hc22245},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5068b, value : 32'h262fb046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5068c, value : 32'haf046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5068d, value : 32'h18040003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5068e, value : 32'h90b0045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5068f, value : 32'hba83033e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50690, value : 32'h90db046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50691, value : 32'hd09019f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50692, value : 32'hc4c6005f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50693, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50694, value : 32'hb067c4c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50695, value : 32'hbb0a756c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50696, value : 32'h2b41f1bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50697, value : 32'hbb2b01cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50698, value : 32'h1c012484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50699, value : 32'he012384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5069a, value : 32'h110e2405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5069b, value : 32'h1c32345},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5069c, value : 32'hf17ab0c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5069d, value : 32'hdb58b084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5069e, value : 32'hb067f176},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5069f, value : 32'hbb08db11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a0, value : 32'h238af1ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a1, value : 32'hb0670008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a2, value : 32'hbb09db09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a3, value : 32'h78e0f1a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a4, value : 32'hc1ac2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a5, value : 32'h45280020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a6, value : 32'h5200c6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a7, value : 32'hfea760c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a8, value : 32'h7704ff8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506a9, value : 32'h200c8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506aa, value : 32'hc6e7810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ab, value : 32'h70b50000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ac, value : 32'hffc20b3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ad, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ae, value : 32'hbf2c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506af, value : 32'h45280020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b0, value : 32'h5200c46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b1, value : 32'hc52760c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b2, value : 32'h70b50000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b3, value : 32'hffc20b20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b4, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b5, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b6, value : 32'h7fe00477},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b7, value : 32'h431800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b8, value : 32'h46cbc2f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506b9, value : 32'h46a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ba, value : 32'h8e4d4050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506bb, value : 32'h2180260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506bc, value : 32'h2140240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506bd, value : 32'h2100250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506be, value : 32'h43304270},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506bf, value : 32'h1b1092d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c0, value : 32'hea144110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c1, value : 32'h8e008ea2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c2, value : 32'h80be2053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c3, value : 32'h7dbbf402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c4, value : 32'h487212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c5, value : 32'ha8640a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c6, value : 32'h42820020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c7, value : 32'h23402002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c8, value : 32'hffef0b0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506c9, value : 32'hf0c94122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ca, value : 32'h81d8e0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506cb, value : 32'h40620071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506cc, value : 32'hffaf0eee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506cd, value : 32'h20788e68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ce, value : 32'hbb240000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506cf, value : 32'hb870b806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d0, value : 32'hae086078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d1, value : 32'h47cb7054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d2, value : 32'h1a188000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d3, value : 32'h223e090f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d4, value : 32'h206120c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d5, value : 32'hb8819710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d6, value : 32'h90db710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d7, value : 32'h9710235e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d8, value : 32'hb710b880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d9, value : 32'he699620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506da, value : 32'h21532030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506db, value : 32'h8190080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506dc, value : 32'h700c0131},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506dd, value : 32'ha706a707},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506de, value : 32'ha704a705},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506df, value : 32'hebe6904},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e0, value : 32'hb600ffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e1, value : 32'h42628e23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e2, value : 32'h43428e04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e3, value : 32'h41227825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e4, value : 32'h2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e5, value : 32'h540240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e6, value : 32'h40e1ae03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e7, value : 32'h500250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e8, value : 32'haba70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506e9, value : 32'h70adffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ea, value : 32'hffaf0e76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506eb, value : 32'h8c54062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ec, value : 32'h4fa80030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ed, value : 32'h41224020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ee, value : 32'h43424262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ef, value : 32'h540240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f0, value : 32'h500250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f1, value : 32'hffef0a96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f2, value : 32'hf05871cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f3, value : 32'h1110829},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f4, value : 32'h225f0911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f5, value : 32'h8e438e04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f6, value : 32'h10a09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f7, value : 32'he80c9712},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f8, value : 32'ha704700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506f9, value : 32'ha706a705},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506fa, value : 32'h6904a707},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506fb, value : 32'hffaf0e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506fc, value : 32'h9620b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506fd, value : 32'h9cbb9c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506fe, value : 32'h40620130},
                          '{ step_type : REG_WRITE, reg_addr : 32'h506ff, value : 32'h3109c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50700, value : 32'h8e23700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50701, value : 32'h8e044262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50702, value : 32'h78254342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50703, value : 32'h20794122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50704, value : 32'h240a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50705, value : 32'hae030540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50706, value : 32'h250a40e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50707, value : 32'ha3e0500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50708, value : 32'h70ccffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50709, value : 32'h96008e22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5070a, value : 32'h90f7404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5070b, value : 32'hb600227e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5070c, value : 32'hb8819712},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5070d, value : 32'h4062b712},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5070e, value : 32'hffaf0de6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5070f, value : 32'h204d2002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50710, value : 32'h4f28e813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50711, value : 32'h42624122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50712, value : 32'h240a4342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50713, value : 32'h250a0540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50714, value : 32'ha0a0500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50715, value : 32'h71ccffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50716, value : 32'h74049600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50717, value : 32'hffaf0e16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50718, value : 32'h8e02b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50719, value : 32'h40a17d02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5071a, value : 32'hffef09c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5071b, value : 32'hf0234122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5071c, value : 32'ha1a2a1a3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5071d, value : 32'ha1a0a1a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5071e, value : 32'h96008ea2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5071f, value : 32'hb600e008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50720, value : 32'h23402017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50721, value : 32'h72082b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50722, value : 32'h15841f22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50723, value : 32'h1f2460b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50724, value : 32'h77041085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50725, value : 32'hffaf0da6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50726, value : 32'h2f057f10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50727, value : 32'h96001341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50728, value : 32'hffaf0fca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50729, value : 32'hb600704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5072a, value : 32'h22d1214f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5072b, value : 32'h1f24f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5072c, value : 32'h8e0410c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5072d, value : 32'h8b6ae03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5072e, value : 32'h40220620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5072f, value : 32'hd62c6d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50730, value : 32'h4308ff8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50731, value : 32'h41224f28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50732, value : 32'h43424262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50733, value : 32'h540240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50734, value : 32'h500250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50735, value : 32'hffef0986},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50736, value : 32'h960070cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50737, value : 32'hb357404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50738, value : 32'hb6001030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50739, value : 32'hff8f0d56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5073a, value : 32'h40e18ea2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5073b, value : 32'h42624122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5073c, value : 32'h240a4342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5073d, value : 32'h250a0540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5073e, value : 32'h9620500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5073f, value : 32'h71ccffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50740, value : 32'h20029600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50741, value : 32'h74042341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50742, value : 32'h8e02b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50743, value : 32'hf10a4910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50744, value : 32'h20028e02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50745, value : 32'hd13200d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50746, value : 32'hd221052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50747, value : 32'h40a1ff8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50748, value : 32'hffef090a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50749, value : 32'h9934122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5074a, value : 32'h9712a2de},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5074b, value : 32'hb712b880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5074c, value : 32'h78e0f1c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5074d, value : 32'hc1abc3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5074e, value : 32'h45284748},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5074f, value : 32'hc0804608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50750, value : 32'hbbe702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50751, value : 32'hda2aff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50752, value : 32'h41838e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50753, value : 32'h8e01b103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50754, value : 32'h8e02b104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50755, value : 32'h8e03b10b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50756, value : 32'h103e0f0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50757, value : 32'h1c0ab10c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50758, value : 32'hf0b3344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50759, value : 32'h1c1a105e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5075a, value : 32'hd523344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5075b, value : 32'hc080ffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5075c, value : 32'h78e0c7c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5075d, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5075e, value : 32'h7fe0046e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5075f, value : 32'h31800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50760, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50761, value : 32'hb100046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50762, value : 32'hb1037fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50763, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50764, value : 32'h7fe0046e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50765, value : 32'h431800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50766, value : 32'h800043c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50767, value : 32'hb30419ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50768, value : 32'hb303d858},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50769, value : 32'h1802153},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5076a, value : 32'h2253b30c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5076b, value : 32'hb30d0040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5076c, value : 32'h800044cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5076d, value : 32'hb305046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5076e, value : 32'hb308781d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5076f, value : 32'h783db300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50770, value : 32'h140206c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50771, value : 32'hb8839440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50772, value : 32'hb30be208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50773, value : 32'h4ed4060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50774, value : 32'hb440ffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50775, value : 32'hc1a4c3e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50776, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50777, value : 32'h4748046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50778, value : 32'h45289640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50779, value : 32'h812253},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5077a, value : 32'h700c4010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5077b, value : 32'hc042c043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5077c, value : 32'h91fc041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5077d, value : 32'hc0400131},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5077e, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5077f, value : 32'ha1001a28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50780, value : 32'ha102a101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50781, value : 32'h6a04a103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50782, value : 32'hffaf0c32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50783, value : 32'h8e02b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50784, value : 32'h781b70f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50785, value : 32'h80f780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50786, value : 32'h20ca2031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50787, value : 32'hd090062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50788, value : 32'h45081005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50789, value : 32'h100e2d05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5078a, value : 32'h781078c9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5078b, value : 32'h26c27510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5078c, value : 32'h78d01061},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5078d, value : 32'h8004208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5078e, value : 32'hd908f792},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5078f, value : 32'hb80ad81f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50790, value : 32'hb2074283},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50791, value : 32'h8002059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50792, value : 32'hb4ab203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50793, value : 32'hc08008e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50794, value : 32'h107c2680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50795, value : 32'h208c78d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50796, value : 32'hf7328fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50797, value : 32'hf388262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50798, value : 32'h2e40f212},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50799, value : 32'h20041300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5079a, value : 32'hf80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5079b, value : 32'hb8887000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5079c, value : 32'hb88bb889},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5079d, value : 32'h30041c06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5079e, value : 32'h20046e17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5079f, value : 32'hf80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a0, value : 32'hf0057c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a1, value : 32'h1c06700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a2, value : 32'h1c0e3005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a3, value : 32'hc0803004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a4, value : 32'h8e00b02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a5, value : 32'hc7c8d908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a6, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a7, value : 32'h1902046a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a8, value : 32'h7fe00043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507a9, value : 32'h78e0a90c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507aa, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ab, value : 32'h49c901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ac, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ad, value : 32'hc1a8c3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ae, value : 32'h47284648},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507af, value : 32'h24404508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b0, value : 32'h702c3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b1, value : 32'hff2f0a3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b2, value : 32'h6e13da1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b3, value : 32'h2044be0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b4, value : 32'h42830400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b5, value : 32'hb203b20b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b6, value : 32'h1f802605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b7, value : 32'h2c580000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b8, value : 32'h2753b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507b9, value : 32'h68371180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ba, value : 32'hb20c7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507bb, value : 32'h11802553},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507bc, value : 32'h78256837},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507bd, value : 32'h78fdb204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507be, value : 32'h140206c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507bf, value : 32'h2605b883},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c0, value : 32'hb8071001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c1, value : 32'hc0807905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c2, value : 32'ha8ab228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c3, value : 32'hd91008e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c4, value : 32'h78e0c7c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c5, value : 32'h1e00710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c6, value : 32'h901c7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c7, value : 32'h7ee00480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c8, value : 32'hb9025021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507c9, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ca, value : 32'h488901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507cb, value : 32'hb1007fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507cc, value : 32'hb9025021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507cd, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ce, value : 32'h48c901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507cf, value : 32'hb1007fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d0, value : 32'h4708c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d1, value : 32'h20846a15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d2, value : 32'h204f0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d3, value : 32'h204f06d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d4, value : 32'h2148068e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d5, value : 32'h77040040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d6, value : 32'h68a17810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d7, value : 32'h400270f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d8, value : 32'h38120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507d9, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507da, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507db, value : 32'hb7670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507dc, value : 32'h70ccffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507dd, value : 32'h1d3f258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507de, value : 32'h78e0c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507df, value : 32'h1600c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e0, value : 32'h800070c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e1, value : 32'h6a21000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e2, value : 32'h792f4408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e3, value : 32'hf4099f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e4, value : 32'h2a44700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e5, value : 32'h4381008d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e6, value : 32'h842380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e7, value : 32'hb20a2b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e8, value : 32'h14828bc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507e9, value : 32'h6e21170b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ea, value : 32'h7040240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507eb, value : 32'h2c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ec, value : 32'h13812415},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ed, value : 32'ha459141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ee, value : 32'h912002c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ef, value : 32'h10440b3d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f0, value : 32'h702c77c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f1, value : 32'he6bff01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f2, value : 32'hf719702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f3, value : 32'h170b1482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f4, value : 32'h79c2d940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f5, value : 32'h7040240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f6, value : 32'h20a8702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f7, value : 32'h241503c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f8, value : 32'h92e11382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507f9, value : 32'h12c40f15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507fa, value : 32'hb119240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507fb, value : 32'he6bf10a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507fc, value : 32'h21ca71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507fd, value : 32'hf0030fe1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507fe, value : 32'h148241c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h507ff, value : 32'h61b91702},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50800, value : 32'h7b2fab20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50801, value : 32'hf74ae3c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50802, value : 32'h10c12415},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50803, value : 32'hc0d9181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50804, value : 32'h91201084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50805, value : 32'h450a17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50806, value : 32'h345242f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50807, value : 32'h22041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50808, value : 32'hee60003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50809, value : 32'hd8c80160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5080a, value : 32'hc6c6d807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5080b, value : 32'hc76c2f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5080c, value : 32'h461001a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5080d, value : 32'h2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5080e, value : 32'h2040708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5080f, value : 32'h46cb0055},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50810, value : 32'h1a448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50811, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50812, value : 32'hca1122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50813, value : 32'hd82520b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50814, value : 32'h8820b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50815, value : 32'h7825881b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50816, value : 32'h50e0889},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50817, value : 32'h10901700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50818, value : 32'h35021a0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50819, value : 32'h407212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5081a, value : 32'h8798f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5081b, value : 32'h40c30044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5081c, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5081d, value : 32'h8698800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5081e, value : 32'h40c2006e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5081f, value : 32'hf93211f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50820, value : 32'ha3c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50821, value : 32'h30581a0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50822, value : 32'h7200a9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50823, value : 32'h23932300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50824, value : 32'h702e4710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50825, value : 32'h22950949},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50826, value : 32'h246e0f3d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50827, value : 32'h704e456a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50828, value : 32'h34581a0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50829, value : 32'heda40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5082a, value : 32'h1a0effef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5082b, value : 32'h120d3498},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5082c, value : 32'h20783082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5082d, value : 32'h120c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5082e, value : 32'h41c33603},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5082f, value : 32'h3021f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50830, value : 32'hff2f0d26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50831, value : 32'h3604120d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50832, value : 32'h75c37146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50833, value : 32'h51e00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50834, value : 32'ha5440ad5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50835, value : 32'h21842380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50836, value : 32'hf1de7126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50837, value : 32'hf1c47106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50838, value : 32'h17942696},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50839, value : 32'hf1b37186},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5083a, value : 32'h78e0c6d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5083b, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5083c, value : 32'hc1a8b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5083d, value : 32'hd8254318},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5083e, value : 32'h1600b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5083f, value : 32'h80007091},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50840, value : 32'h44d3122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50841, value : 32'h489004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50842, value : 32'h24428820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50843, value : 32'h881b2210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50844, value : 32'h20787825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50845, value : 32'h204000c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50846, value : 32'h16000055},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50847, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50848, value : 32'h8e1122b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50849, value : 32'h40c30444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5084a, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5084b, value : 32'h8d18800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5084c, value : 32'h212f046e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5084d, value : 32'h9ee0447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5084e, value : 32'h40630720},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5084f, value : 32'h23182940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50850, value : 32'h706e4118},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50851, value : 32'h34ee09b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50852, value : 32'h22002b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50853, value : 32'h200570ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50854, value : 32'hc8090601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50855, value : 32'h69127905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50856, value : 32'h20054230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50857, value : 32'h90040f96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50858, value : 32'h215a0320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50859, value : 32'hc7802a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5085a, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5085b, value : 32'h7fb4c00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5085c, value : 32'h4c02015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5085d, value : 32'h603278b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5085e, value : 32'h11a06119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5085f, value : 32'h20340101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50860, value : 32'h80000f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50861, value : 32'hb740becc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50862, value : 32'h1c08b722},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50863, value : 32'h25053004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50864, value : 32'h68d21480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50865, value : 32'h15002605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50866, value : 32'he009d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50867, value : 32'hb7059000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50868, value : 32'h140e2605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50869, value : 32'he009ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5086a, value : 32'hb7079600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5086b, value : 32'h160071a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5086c, value : 32'hdb32100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5086d, value : 32'h1c129564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5086e, value : 32'h40a23004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5086f, value : 32'h5e00cbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50870, value : 32'h706cc180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50871, value : 32'h2305c485},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50872, value : 32'h14020480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50873, value : 32'hb8021501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50874, value : 32'h20057164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50875, value : 32'hb2200502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50876, value : 32'h4012005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50877, value : 32'hbeb9401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50878, value : 32'hb1008564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50879, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5087a, value : 32'hee8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5087b, value : 32'h141ce885},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5087c, value : 32'h1e003100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5087d, value : 32'h71662004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5087e, value : 32'ha2540b4d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5087f, value : 32'hf18f7126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50880, value : 32'h1404c0a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50881, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50882, value : 32'hc1a3c3f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50883, value : 32'hd8254018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50884, value : 32'h1600b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50885, value : 32'h8000708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50886, value : 32'h1600122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50887, value : 32'h80007092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50888, value : 32'h88200187},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50889, value : 32'h881b7056},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5088a, value : 32'h242122ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5088b, value : 32'h20787825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5088c, value : 32'h204000c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5088d, value : 32'h16000053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5088e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5088f, value : 32'h8db122b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50890, value : 32'h40c30344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50891, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50892, value : 32'h8cb8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50893, value : 32'h79af036e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50894, value : 32'h72008d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50895, value : 32'h2d404003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50896, value : 32'h47101316},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50897, value : 32'hfb1700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50898, value : 32'h2840242e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50899, value : 32'h702e2200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5089a, value : 32'h5812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5089b, value : 32'h2105c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5089c, value : 32'h25050015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5089d, value : 32'hc1812440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5089e, value : 32'h260568d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5089f, value : 32'h90041f8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a0, value : 32'ha860048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a1, value : 32'h97000260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a2, value : 32'h1f8e2605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a3, value : 32'h409004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a4, value : 32'ha769600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a5, value : 32'hc1820260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a6, value : 32'h30821409},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a7, value : 32'h30811405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a8, value : 32'h483223d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508a9, value : 32'h480213d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508aa, value : 32'hc022786b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ab, value : 32'he810f410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ac, value : 32'h8022254},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ad, value : 32'h2154c321},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ae, value : 32'h77040801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508af, value : 32'h1c097764},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b0, value : 32'hc0623082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b1, value : 32'h1c05c361},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b2, value : 32'hf0033042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b3, value : 32'h792fc321},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b4, value : 32'h7252f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b5, value : 32'h262fc140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b6, value : 32'h272f0087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b7, value : 32'h740c00c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b8, value : 32'h41c34222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508b9, value : 32'h7025a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ba, value : 32'hc1e43a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508bb, value : 32'h240a0160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508bc, value : 32'hcca0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508bd, value : 32'hc0810160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508be, value : 32'hcc2b700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508bf, value : 32'hc0820160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c0, value : 32'h2140b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c1, value : 32'h86f2040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c2, value : 32'h712e84e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c3, value : 32'h8537106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c4, value : 32'h71a5a254},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c5, value : 32'hc7d8f191},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c6, value : 32'h88606038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c7, value : 32'ha8607b44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c8, value : 32'h83104b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508c9, value : 32'h184b7b44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ca, value : 32'h109600c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508cb, value : 32'h7b440083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508cc, value : 32'hc21896},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508cd, value : 32'h8310e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ce, value : 32'h7fe07a64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508cf, value : 32'h8218e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d0, value : 32'h2482c3f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d1, value : 32'h250a3306},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d2, value : 32'h230a2180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d3, value : 32'h40702100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d4, value : 32'h45284650},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d5, value : 32'h248a4410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d6, value : 32'h24407001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d7, value : 32'h218a3011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d8, value : 32'hc0800fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508d9, value : 32'h14020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508da, value : 32'h1804b021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508db, value : 32'h18000015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508dc, value : 32'hd8ff0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508dd, value : 32'h301c1c82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508de, value : 32'h38002456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508df, value : 32'h42d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e0, value : 32'h47cb0a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e1, value : 32'h1a448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e2, value : 32'h300d87},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e3, value : 32'h7c31802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e4, value : 32'h1481251f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e5, value : 32'h184228a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e6, value : 32'h2f80241f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e7, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e8, value : 32'h2184209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508e9, value : 32'h70026038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ea, value : 32'hd3e60f9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508eb, value : 32'hc080feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ec, value : 32'h8400b1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ed, value : 32'h3008d9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ee, value : 32'h1600dd3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ef, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f0, value : 32'h80f0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f1, value : 32'h1600009f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f2, value : 32'h8000708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f3, value : 32'hb020120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f4, value : 32'h24560840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f5, value : 32'h24003843},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f6, value : 32'h3f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f7, value : 32'ha901010c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f8, value : 32'h712c40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508f9, value : 32'h2e00d36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508fa, value : 32'h148a704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508fb, value : 32'h248a370c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508fc, value : 32'h700c7001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508fd, value : 32'h20a8c380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508fe, value : 32'h93200300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h508ff, value : 32'ha0f9341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50900, value : 32'h4a310064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50901, value : 32'h798a7124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50902, value : 32'h74646038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50903, value : 32'h2180f050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50904, value : 32'hea12084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50905, value : 32'hb11a344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50906, value : 32'hb152090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50907, value : 32'hd0d2051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50908, value : 32'hf006101f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50909, value : 32'h101f0d09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5090a, value : 32'hf1f571a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5090b, value : 32'hefd70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5090c, value : 32'hd139405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5090d, value : 32'h25002031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5090e, value : 32'h10201680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5090f, value : 32'he4d0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50910, value : 32'ha8e1000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50911, value : 32'h251a0840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50912, value : 32'h70141482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50913, value : 32'h2f81241f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50914, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50915, value : 32'h40c3708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50916, value : 32'h1b468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50917, value : 32'h42c16159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50918, value : 32'h184229a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50919, value : 32'hf207623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5091a, value : 32'h91616059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5091b, value : 32'h37011482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5091c, value : 32'h62f94b34},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5091d, value : 32'h1100620a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5091e, value : 32'h242f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5091f, value : 32'h4a130306},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50920, value : 32'hf9ac080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50921, value : 32'hc2800060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50922, value : 32'hf1d371c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50923, value : 32'h7001248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50924, value : 32'hc380700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50925, value : 32'h30020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50926, value : 32'h5021302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50927, value : 32'h5011302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50928, value : 32'h61197150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50929, value : 32'h71247942},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5092a, value : 32'h4620ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5092b, value : 32'h78e0c7d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5092c, value : 32'h4308c0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5092d, value : 32'h7001248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5092e, value : 32'h700c70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5092f, value : 32'h7c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50930, value : 32'h44cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50931, value : 32'h7d9b28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50932, value : 32'h130f231f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50933, value : 32'hbc227d6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50934, value : 32'h67bf7c2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50935, value : 32'h4448679d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50936, value : 32'h1184249f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50937, value : 32'h44cb659d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50938, value : 32'h1a448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50939, value : 32'h71c57dd5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5093a, value : 32'h64bc6597},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5093b, value : 32'h74f19481},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5093c, value : 32'h7ce2641c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5093d, value : 32'h20ca7185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5093e, value : 32'hc4c60306},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5093f, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50940, value : 32'h70851e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50941, value : 32'h88900c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50942, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50943, value : 32'h921c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50944, value : 32'h271400a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50945, value : 32'haa6000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50946, value : 32'h40a00160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50947, value : 32'ha9eb40a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50948, value : 32'h40c00160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50949, value : 32'h2740b40c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5094a, value : 32'hf00c0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5094b, value : 32'h1600a8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5094c, value : 32'hb40a4060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5094d, value : 32'h1600a86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5094e, value : 32'hb40c4080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5094f, value : 32'h4802740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50950, value : 32'hc0d19000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50951, value : 32'h1f1c7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50952, value : 32'h78e00004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50953, value : 32'h8e9c3f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50954, value : 32'hc1a40071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50955, value : 32'h47cb712e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50956, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50957, value : 32'h20f509d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50958, value : 32'h447202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50959, value : 32'h900813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5095a, value : 32'h51081b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5095b, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5095c, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5095d, value : 32'h1600f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5095e, value : 32'h80007081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5095f, value : 32'h9af0040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50960, value : 32'hb0600d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50961, value : 32'h9c601c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50962, value : 32'h706e0600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50963, value : 32'h20b50b9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50964, value : 32'hdba4062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50965, value : 32'h702c00a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50966, value : 32'h20408fa0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50967, value : 32'h8f010a94},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50968, value : 32'h3440887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50969, value : 32'h13122d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5096a, value : 32'h2205c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5096b, value : 32'hc1802510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5096c, value : 32'h4002005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5096d, value : 32'h4c22116},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5096e, value : 32'h46cbb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5096f, value : 32'h9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50970, value : 32'h78c57ab4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50971, value : 32'hb5f9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50972, value : 32'hb2002071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50973, value : 32'h34021f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50974, value : 32'h422279b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50975, value : 32'h9124716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50976, value : 32'h603844a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50977, value : 32'h41e41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50978, value : 32'h78100006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50979, value : 32'h2252f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5097a, value : 32'h1d62841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5097b, value : 32'h1552553},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5097c, value : 32'h260a740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5097d, value : 32'h9120580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5097e, value : 32'h270a0160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5097f, value : 32'h2e400540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50980, value : 32'h20052180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50981, value : 32'hc8090541},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50982, value : 32'h4822005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50983, value : 32'h4002005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50984, value : 32'hb802ba02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50985, value : 32'h22057e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50986, value : 32'h90040f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50987, value : 32'hb22000a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50988, value : 32'h71a5b620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50989, value : 32'h7166f1bd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5098a, value : 32'h7126f1b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5098b, value : 32'ha5af198},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5098c, value : 32'h730c01e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5098d, value : 32'h78e0c7d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5098e, value : 32'h41c3c2f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5098f, value : 32'h1d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50990, value : 32'h16008c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50991, value : 32'h43d3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50992, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50993, value : 32'h208e1300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50994, value : 32'h800142d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50995, value : 32'h22164d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50996, value : 32'h1301238d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50997, value : 32'h76102080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50998, value : 32'h2d0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50999, value : 32'h23802216},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5099a, value : 32'hcc2390e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5099b, value : 32'h702ee819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5099c, value : 32'h40f144b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5099d, value : 32'h21041400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5099e, value : 32'h42c1740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5099f, value : 32'h1d241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a0, value : 32'h8860003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a1, value : 32'h43220160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a2, value : 32'h25001402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a3, value : 32'h20087126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a4, value : 32'h27092010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a5, value : 32'hcc23100f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a6, value : 32'ha00409dd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a7, value : 32'h40f1f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a8, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509a9, value : 32'h201d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509aa, value : 32'h85e42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ab, value : 32'h43020160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ac, value : 32'h740c7702},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ad, value : 32'h41c37ffd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ae, value : 32'h201d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509af, value : 32'h1310274e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b0, value : 32'h232f42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b1, value : 32'h8420408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b2, value : 32'h41700160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b3, value : 32'h2e406f14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b4, value : 32'h20051343},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b5, value : 32'h29402010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b6, value : 32'h20052100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b7, value : 32'hc80903df},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b8, value : 32'h2300718c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509b9, value : 32'hf8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ba, value : 32'h726d1000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509bb, value : 32'h903842c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509bc, value : 32'hc0f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509bd, value : 32'h208a0031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509be, value : 32'h208a1c15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509bf, value : 32'h20051415},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c0, value : 32'hb9021001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c1, value : 32'h1016218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c2, value : 32'hc0d7945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c3, value : 32'h91200031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c4, value : 32'h1815218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c5, value : 32'hc2184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c6, value : 32'h2105708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c7, value : 32'h210507cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c8, value : 32'hb9021001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509c9, value : 32'h794572ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ca, value : 32'h912070cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509cb, value : 32'hc2184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509cc, value : 32'h20472005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509cd, value : 32'h2012600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ce, value : 32'h1e2105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509cf, value : 32'h30c12605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d0, value : 32'h7945b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d1, value : 32'h2605b1e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d2, value : 32'hb9023301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d3, value : 32'hb1e07945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d4, value : 32'h2412600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d5, value : 32'h62105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d6, value : 32'hc12605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d7, value : 32'h7945b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d8, value : 32'h1c41900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509d9, value : 32'h3012605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509da, value : 32'h71ccb902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509db, value : 32'h258d7945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509dc, value : 32'h1900093f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509dd, value : 32'h238c01c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509de, value : 32'he5081ffe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509df, value : 32'hf16f71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e0, value : 32'h78e0c6d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e1, value : 32'h14422aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e2, value : 32'h10421aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e3, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e4, value : 32'ha0410458},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e5, value : 32'ha0207fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e6, value : 32'h700026f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e7, value : 32'hf688000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e8, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509e9, value : 32'h803c2042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ea, value : 32'h12220e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509eb, value : 32'h40212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ec, value : 32'h7fe06909},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ed, value : 32'h78e07810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ee, value : 32'h4010c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ef, value : 32'h4568730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f0, value : 32'h8c64648},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f1, value : 32'h472801e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f2, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f3, value : 32'h88001140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f4, value : 32'h1600e810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f5, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f6, value : 32'h8190001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f7, value : 32'hd80f00ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f8, value : 32'h42e14102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509f9, value : 32'h708c43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509fa, value : 32'h8600e8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509fb, value : 32'hc6c845a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509fc, value : 32'h4102d80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509fd, value : 32'h43c142e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509fe, value : 32'h8600cde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h509ff, value : 32'hc6c844a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a00, value : 32'hea06c0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a01, value : 32'h248a76ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a02, value : 32'hf005100f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a03, value : 32'h248add07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a04, value : 32'h2278100e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a05, value : 32'hba060002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a06, value : 32'h2204e23f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a07, value : 32'h7984004f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a08, value : 32'h7c0479b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a09, value : 32'h2c0169d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a0a, value : 32'h66fe1340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a0b, value : 32'he176836},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a0c, value : 32'h61581064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a0d, value : 32'h76107810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a0e, value : 32'h108d24c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a0f, value : 32'h6698f703},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a10, value : 32'hc8094834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a11, value : 32'hb8027865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a12, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a13, value : 32'h3c009004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a14, value : 32'hc4c6b080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a15, value : 32'h806c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a16, value : 32'h86602c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a17, value : 32'h450802e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a18, value : 32'h2a00c4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a19, value : 32'h609860bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a1a, value : 32'h412044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a1b, value : 32'h780f6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a1c, value : 32'h7012089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a1d, value : 32'h30021a04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a1e, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a1f, value : 32'h4008c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a20, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a21, value : 32'h8151229},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a22, value : 32'h88401071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a23, value : 32'h70831600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a24, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a25, value : 32'hf2957074},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a26, value : 32'h1030080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a27, value : 32'h100c2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a28, value : 32'hf0038865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a29, value : 32'hec848863},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a2a, value : 32'hf0038886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a2b, value : 32'hc8098884},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a2c, value : 32'hdd787034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a2d, value : 32'hc0f706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a2e, value : 32'h25ca10e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a2f, value : 32'h70cd1822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a30, value : 32'h2178f01f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a31, value : 32'h655d0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a32, value : 32'h70cdb903},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a33, value : 32'h462140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a34, value : 32'h3012b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a35, value : 32'h7180240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a36, value : 32'h702d61b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a37, value : 32'h69f27905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a38, value : 32'h30020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a39, value : 32'h13c12105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a3a, value : 32'h10102180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a3b, value : 32'hb99cb992},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a3c, value : 32'h9120b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a3d, value : 32'h38e2108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a3e, value : 32'h71647391},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a3f, value : 32'hb802f7aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a40, value : 32'h343236f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a41, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a42, value : 32'h209004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a43, value : 32'h730c9080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a44, value : 32'h5091302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a45, value : 32'h100c2479},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a46, value : 32'h210c8b20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a47, value : 32'h9f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a48, value : 32'h20ca0c7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a49, value : 32'h723400ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a4a, value : 32'h23ca7c9b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a4b, value : 32'h718510e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a4c, value : 32'h2300ddff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a4d, value : 32'h7c3d130b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a4e, value : 32'h2e01e407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a4f, value : 32'h7461130c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a50, value : 32'h208a641c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a51, value : 32'h20ca0fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a52, value : 32'h78c40341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a53, value : 32'h2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a54, value : 32'h2356641c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a55, value : 32'h10000940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a56, value : 32'h609800c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a57, value : 32'h2048780e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a58, value : 32'hca070003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a59, value : 32'h813e80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a5a, value : 32'h12220231},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a5b, value : 32'hc17370c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a5c, value : 32'h1f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a5d, value : 32'h8176815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a5e, value : 32'hc130251},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a5f, value : 32'h1f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a60, value : 32'h9177196},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a61, value : 32'hbb620111},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a62, value : 32'h210cf007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a63, value : 32'h9f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a64, value : 32'h23c22156},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a65, value : 32'h202f0066},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a66, value : 32'h242f0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a67, value : 32'h785500c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a68, value : 32'h7441c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a69, value : 32'h70c30003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a6a, value : 32'h4608000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a6b, value : 32'h6b09b060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a6c, value : 32'h43017810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a6d, value : 32'hfeef0c32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a6e, value : 32'h3c0207c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a6f, value : 32'h40c3c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a70, value : 32'h4608000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a71, value : 32'h90207855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a72, value : 32'hc6c6b021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a73, value : 32'hc80943e3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a74, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a75, value : 32'h90080f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a76, value : 32'h90000014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a77, value : 32'h2a00e5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a78, value : 32'h2044b8c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a79, value : 32'h781d0041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a7a, value : 32'h7b006038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a7b, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a7c, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a7d, value : 32'hd98e3905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a7e, value : 32'hb99f70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a7f, value : 32'hc652da80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a80, value : 32'h11f88900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a81, value : 32'hc653808d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a82, value : 32'h8908c048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a83, value : 32'hc654702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a84, value : 32'hc044c655},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a85, value : 32'hfeaf0eea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a86, value : 32'h3e402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a87, value : 32'h702cc099},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a88, value : 32'hededa80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a89, value : 32'hc658feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a8a, value : 32'h14002544},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a8b, value : 32'hc64e720e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a8c, value : 32'hc650c64f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a8d, value : 32'hc64ac651},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a8e, value : 32'hc64cc64b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a8f, value : 32'hc657c64d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a90, value : 32'hc008c047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a91, value : 32'h807e2053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a92, value : 32'h4ec8f212},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a93, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a94, value : 32'h79d6c192},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a95, value : 32'h5e00e8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a96, value : 32'h1600714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a97, value : 32'h8000708b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a98, value : 32'h1600122b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a99, value : 32'h80007082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a9a, value : 32'hf02d122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a9b, value : 32'h708b1600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a9c, value : 32'h122b8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a9d, value : 32'h70821600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a9e, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a9f, value : 32'h10a40b47},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa0, value : 32'h1f012654},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa1, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa2, value : 32'h68324448},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa3, value : 32'h13832c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa4, value : 32'h7200244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa5, value : 32'h70ad7b25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa6, value : 32'h48020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa7, value : 32'h24556e16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa8, value : 32'h671f3e4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aa9, value : 32'h671f6c14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aaa, value : 32'h12802d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aab, value : 32'h7fb47865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aac, value : 32'h71a5b892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aad, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aae, value : 32'hb7009000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aaf, value : 32'h71857471},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab0, value : 32'hb47f7a6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab1, value : 32'h6e3610a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab2, value : 32'h611b6a14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab3, value : 32'h1f412654},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab4, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab5, value : 32'h2a4068b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab6, value : 32'hc099038f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab7, value : 32'h244a7fa5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab8, value : 32'h60797200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ab9, value : 32'h20a8700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aba, value : 32'h27050340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50abb, value : 32'h2080100c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50abc, value : 32'hbc920010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50abd, value : 32'hbc9fbc9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50abe, value : 32'h19029480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50abf, value : 32'he3100314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac0, value : 32'h71447271},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac1, value : 32'hc007f7a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac2, value : 32'h4edae809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac3, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac4, value : 32'h79d6c18a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac5, value : 32'h5e00dce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac6, value : 32'hc004714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac7, value : 32'h13e0815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac8, value : 32'hc8094ed8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ac9, value : 32'hc18e7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aca, value : 32'hdba79d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50acb, value : 32'h714c05e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50acc, value : 32'h227e208d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50acd, value : 32'hc09971cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ace, value : 32'h2054702f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50acf, value : 32'hc0430800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad0, value : 32'h3e402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad1, value : 32'h8002054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad2, value : 32'h301b140c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad3, value : 32'hc08cc041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad4, value : 32'hc001c045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad5, value : 32'h140cc046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad6, value : 32'hc5973017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad7, value : 32'h30161404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad8, value : 32'h3c122454},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ad9, value : 32'h22147dd4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ada, value : 32'h24402392},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50adb, value : 32'h710e3c18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50adc, value : 32'ha380200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50add, value : 32'h1600f2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ade, value : 32'h8000709e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50adf, value : 32'h1600122b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae0, value : 32'h8000708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae1, value : 32'hc007122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae2, value : 32'h706de8bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae3, value : 32'h33240e65},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae4, value : 32'h1414700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae5, value : 32'hc7973009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae6, value : 32'h140f2714},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae7, value : 32'h33002602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae8, value : 32'h33072014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ae9, value : 32'h462040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aea, value : 32'h706d700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aeb, value : 32'h13092114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aec, value : 32'h15001102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aed, value : 32'hc32762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aee, value : 32'hda400120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aef, value : 32'hb5004408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af0, value : 32'h5001702},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af1, value : 32'hc22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af2, value : 32'hda400120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af3, value : 32'h222fb700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af4, value : 32'h9d2002c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af5, value : 32'hb700b580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af6, value : 32'h7902780e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af7, value : 32'h4b2208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af8, value : 32'h49109d20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50af9, value : 32'h206212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50afa, value : 32'h93f268d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50afb, value : 32'h82108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50afc, value : 32'h200c96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50afd, value : 32'h2c6202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50afe, value : 32'h202f4400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50aff, value : 32'hf0960206},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b00, value : 32'hc0066c34},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b01, value : 32'h482000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b02, value : 32'h2014c097},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b03, value : 32'hc0980411},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b04, value : 32'h4052014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b05, value : 32'h20442700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b06, value : 32'h30472300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b07, value : 32'h20462600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b08, value : 32'h706d702d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b09, value : 32'h33240ef9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b0a, value : 32'h11802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b0b, value : 32'h2053c008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b0c, value : 32'hf219807e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b0d, value : 32'h2016c092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b0e, value : 32'h20160381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b0f, value : 32'h21f40400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b10, value : 32'h20f40301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b11, value : 32'hb9260300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b12, value : 32'h1a00b826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b13, value : 32'h1d002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b14, value : 32'h12000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b15, value : 32'h4f11214f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b16, value : 32'h246202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b17, value : 32'h492008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b18, value : 32'h244af018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b19, value : 32'h43c07200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b1a, value : 32'h20a84201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b1b, value : 32'h12020500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b1c, value : 32'hb8260500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b1d, value : 32'h20041a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b1e, value : 32'h5001302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b1f, value : 32'h1d00b826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b20, value : 32'h12000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b21, value : 32'h4f11214f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b22, value : 32'h246202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b23, value : 32'h492008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b24, value : 32'h2200234a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b25, value : 32'h2100250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b26, value : 32'h21c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b27, value : 32'h25001402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b28, value : 32'hb46762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b29, value : 32'hda400120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b2a, value : 32'h762cb500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b2b, value : 32'h25001502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b2c, value : 32'h1200b36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b2d, value : 32'h1900da40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b2e, value : 32'h790e2004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b2f, value : 32'h78229d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b30, value : 32'h2c6212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b31, value : 32'h2b3f238d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b32, value : 32'hb2108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b33, value : 32'h83dc004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b34, value : 32'h2440013e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b35, value : 32'h762c3e13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b36, value : 32'h23802316},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b37, value : 32'hb0ada40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b38, value : 32'h20f40120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b39, value : 32'hb5000300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b3a, value : 32'h24002316},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b3b, value : 32'hda40762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b3c, value : 32'h1200af6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b3d, value : 32'h30020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b3e, value : 32'h20041900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b3f, value : 32'h4f10780e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b40, value : 32'h2c6212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b41, value : 32'hb2108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b42, value : 32'h4042440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b43, value : 32'h4072740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b44, value : 32'h4062640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b45, value : 32'h14082040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b46, value : 32'hf1867185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b47, value : 32'h200b6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b48, value : 32'h4400780e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b49, value : 32'h2c6202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b4a, value : 32'hb5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b4b, value : 32'h202f4110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b4c, value : 32'hc1890647},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b4d, value : 32'h38a47cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b4e, value : 32'h61190003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b4f, value : 32'h190042c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b50, value : 32'hc1960442},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b51, value : 32'h41e16038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b52, value : 32'h1021800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b53, value : 32'h9ba740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b54, value : 32'h43020120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b55, value : 32'h1401274f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b56, value : 32'h42c1740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b57, value : 32'h9aa4302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b58, value : 32'h240a0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b59, value : 32'h71270440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b5a, value : 32'h203f2780},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b5b, value : 32'h203f2680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b5c, value : 32'h32182042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b5d, value : 32'h5fc7016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b5e, value : 32'h7706ffe2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b5f, value : 32'h2380c006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b60, value : 32'h2080303f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b61, value : 32'h70d5003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b62, value : 32'h77c5c046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b63, value : 32'hb868c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b64, value : 32'hffe205c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b65, value : 32'hc136c045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b66, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b67, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b68, value : 32'hd841e803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b69, value : 32'hd826f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b6a, value : 32'h140cb89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b6b, value : 32'h700e3015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b6c, value : 32'h1801712e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b6d, value : 32'h14590052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b6e, value : 32'ha8203081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b6f, value : 32'ha829c129},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b70, value : 32'h30811425},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b71, value : 32'hc007a82a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b72, value : 32'h172079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b73, value : 32'h34001c08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b74, value : 32'h34001c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b75, value : 32'h3014140c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b76, value : 32'h3b982454},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b77, value : 32'h3c162454},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b78, value : 32'h34532014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b79, value : 32'h24562614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b7a, value : 32'h273971ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b7b, value : 32'h704e1440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b7c, value : 32'h5c02006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b7d, value : 32'hb8e070cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b7e, value : 32'h1600f4cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b7f, value : 32'h8000708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b80, value : 32'h1600122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b81, value : 32'h80007092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b82, value : 32'h2014122b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b83, value : 32'hc00133ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b84, value : 32'h700d70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b85, value : 32'h25006c34},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b86, value : 32'h24002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b87, value : 32'h20002049},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b88, value : 32'h74520046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b89, value : 32'h2d015a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b8a, value : 32'hc00878ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b8b, value : 32'h807e2053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b8c, value : 32'hc092f23f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b8d, value : 32'h2016762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b8e, value : 32'hda400440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b8f, value : 32'h12009aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b90, value : 32'h30020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b91, value : 32'h43cb4700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b92, value : 32'hffff0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b93, value : 32'h3000264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b94, value : 32'h200254a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b95, value : 32'h20041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b96, value : 32'hc1996f16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b97, value : 32'h6c146119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b98, value : 32'h762c6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b99, value : 32'h78020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b9a, value : 32'h120097e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b9b, value : 32'h212fda40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b9c, value : 32'h264002c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b9d, value : 32'h258d305e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b9e, value : 32'h21090cbf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50b9f, value : 32'hb600000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba0, value : 32'h81dc004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba1, value : 32'hc08e013e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba2, value : 32'h78f6762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba3, value : 32'h95ada40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba4, value : 32'h20f40120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba5, value : 32'h23090300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba6, value : 32'hb600100b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba7, value : 32'h2c6212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba8, value : 32'h1c6202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ba9, value : 32'h79ae7822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50baa, value : 32'hd2108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bab, value : 32'h274af020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bac, value : 32'h260a0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bad, value : 32'h250a3240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bae, value : 32'h15020180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50baf, value : 32'h762c0500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb0, value : 32'h1200926},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb1, value : 32'h4308da40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb2, value : 32'h35001602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb3, value : 32'h91a762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb4, value : 32'hda400120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb5, value : 32'h2c6222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb6, value : 32'h4a31790e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb7, value : 32'h278d7aae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb8, value : 32'h22080bff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bb9, value : 32'hb600004d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bba, value : 32'h22c41e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bbb, value : 32'h14600f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bbc, value : 32'h1200234a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bbd, value : 32'h240250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bbe, value : 32'h100270a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bbf, value : 32'h5001702},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc0, value : 32'h8e6762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc1, value : 32'hda400120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc2, value : 32'h20041b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc3, value : 32'h1502762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc4, value : 32'h8d60500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc5, value : 32'hda400120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc6, value : 32'h790eb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc7, value : 32'h21401300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc8, value : 32'h212f7822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bc9, value : 32'h238d0206},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bca, value : 32'h21081b3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bcb, value : 32'hc0040008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bcc, value : 32'h13e083f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bcd, value : 32'h3e0b2440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bce, value : 32'h2316762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bcf, value : 32'hda401440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd0, value : 32'h12008a6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd1, value : 32'h30020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd2, value : 32'h13cb2316},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd3, value : 32'h20041b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd4, value : 32'hda40762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd5, value : 32'h1200892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd6, value : 32'h130023f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd7, value : 32'h790eb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd8, value : 32'h21401300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bd9, value : 32'h212f7822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bda, value : 32'h21080206},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bdb, value : 32'h24400008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bdc, value : 32'h21400404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bdd, value : 32'h26401409},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bde, value : 32'h71850406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bdf, value : 32'h90af153},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be0, value : 32'h42100000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be1, value : 32'h200902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be2, value : 32'h206202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be3, value : 32'h202f4608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be4, value : 32'hc1800407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be5, value : 32'h45cb6119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be6, value : 32'h3038e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be7, value : 32'hc182a9c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be8, value : 32'h41a16038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50be9, value : 32'h4821800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bea, value : 32'h4222740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50beb, value : 32'hf5a43e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bec, value : 32'h240a00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bed, value : 32'h254f0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bee, value : 32'h740c1401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bef, value : 32'h43e14222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf0, value : 32'he00f46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf1, value : 32'h248044c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf2, value : 32'h7106203f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf3, value : 32'h77e570f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf4, value : 32'hc001f50d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf5, value : 32'h203f2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf6, value : 32'h3f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf7, value : 32'h77267036},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf8, value : 32'hffe205f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bf9, value : 32'hc222c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bfa, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bfb, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bfc, value : 32'hd943e803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bfd, value : 32'hd928f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bfe, value : 32'h1409b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50bff, value : 32'h19013080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c00, value : 32'h19010092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c01, value : 32'h140a0012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c02, value : 32'h19013080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c03, value : 32'h19010012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c04, value : 32'hc0200492},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c05, value : 32'h121901},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c06, value : 32'h30801401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c07, value : 32'h1402a900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c08, value : 32'ha9013080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c09, value : 32'h2480a9c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c0a, value : 32'h14043905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c0b, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c0c, value : 32'h40d3c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c0d, value : 32'hc0c902c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c0e, value : 32'h21111000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c0f, value : 32'h2d0d2040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c10, value : 32'h214f71ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c11, value : 32'hb5e02100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c12, value : 32'h180070cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c13, value : 32'h40c32004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c14, value : 32'ha48007bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c15, value : 32'h10151d04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c16, value : 32'h1df0702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c17, value : 32'h1df093c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c18, value : 32'hf329384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c19, value : 32'hb5e00460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c1a, value : 32'he8069502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c1b, value : 32'h4600e9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c1c, value : 32'hf1fcd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c1d, value : 32'hb5deb5c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c1e, value : 32'hb5deb5fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c1f, value : 32'h24441800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c20, value : 32'h78e0c6ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c21, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c22, value : 32'h88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c23, value : 32'h720813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c24, value : 32'h7810b907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c25, value : 32'h77046038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c26, value : 32'h412804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c27, value : 32'h7813f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c28, value : 32'h28057810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c29, value : 32'h79130040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c2a, value : 32'h782e7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c2b, value : 32'hd9ec2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c2c, value : 32'h450807e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c2d, value : 32'h16007014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c2e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c2f, value : 32'h74cd0160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c30, value : 32'h11e226ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c31, value : 32'hee2e805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c32, value : 32'h712cffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c33, value : 32'h1600f009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c34, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c35, value : 32'hb8e20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c36, value : 32'h20ca700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c37, value : 32'h7f1003e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c38, value : 32'h40e141c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c39, value : 32'h716c42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c3a, value : 32'ha9e708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c3b, value : 32'h70ac0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c3c, value : 32'h702c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c3d, value : 32'h716c42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c3e, value : 32'h8e008d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c3f, value : 32'h40e1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c40, value : 32'h42a141c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c41, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c42, value : 32'h600a7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c43, value : 32'h710c70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c44, value : 32'h42a1702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c45, value : 32'h8ba716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c46, value : 32'h708c08e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c47, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c48, value : 32'h40d3c2f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c49, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c4a, value : 32'h20911000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c4b, value : 32'h46304550},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c4c, value : 32'ha942040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c4d, value : 32'h23122940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c4e, value : 32'h20801001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c4f, value : 32'h46408af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c50, value : 32'h25132205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c51, value : 32'h2005c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c52, value : 32'h47cb04c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c53, value : 32'h9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c54, value : 32'h41c3b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c55, value : 32'h303e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c56, value : 32'h422278e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c57, value : 32'h740c90c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c58, value : 32'h265343c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c59, value : 32'hda21144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c5a, value : 32'h23ad00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c5b, value : 32'hd230982},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c5c, value : 32'h740c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c5d, value : 32'h3e941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c5e, value : 32'hd8e0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c5f, value : 32'h160000c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c60, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c61, value : 32'hb8060008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c62, value : 32'h100d2e09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c63, value : 32'he0df00b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c64, value : 32'h26402030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c65, value : 32'hf007180d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c66, value : 32'h18340e0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c67, value : 32'h264270ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c68, value : 32'h2553180d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c69, value : 32'h25ad114e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c6a, value : 32'hd111982},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c6b, value : 32'h740c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c6c, value : 32'h3ea41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c6d, value : 32'hf00b0002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c6e, value : 32'h20100e0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c6f, value : 32'h3eb41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c70, value : 32'hf0050002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c71, value : 32'h3ec41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c72, value : 32'h42a10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c73, value : 32'he00d3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c74, value : 32'h6d1643c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c75, value : 32'h20082296},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c76, value : 32'hc8097e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c77, value : 32'h4c02005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c78, value : 32'hb8027126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c79, value : 32'hb7c07f05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c7a, value : 32'hd62f1a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c7b, value : 32'hc6d40580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c7c, value : 32'h800140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c7d, value : 32'h88204e89},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c7e, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c7f, value : 32'h728000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c80, value : 32'h20447824},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c81, value : 32'h7fe00800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c82, value : 32'h2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c83, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c84, value : 32'h8a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c85, value : 32'h7fe0b8c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c86, value : 32'h402078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c87, value : 32'h800141c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c88, value : 32'h89204e91},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c89, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c8a, value : 32'h928000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c8b, value : 32'h20447825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c8c, value : 32'h7fe00800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c8d, value : 32'h78e0b825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c8e, value : 32'h800141c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c8f, value : 32'h89204e7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c90, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c91, value : 32'h628000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c92, value : 32'h20847825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c93, value : 32'h7fe00001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c94, value : 32'h78e0b826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c95, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c96, value : 32'h8e8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c97, value : 32'h7fe0b8c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c98, value : 32'h2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c99, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c9a, value : 32'h968000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c9b, value : 32'h4002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c9c, value : 32'hb8247fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c9d, value : 32'hb7c81cf4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c9e, value : 32'h87f4200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50c9f, value : 32'h1c040065},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca0, value : 32'h78523001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca1, value : 32'h6038700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca2, value : 32'hb8224340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca3, value : 32'h71044140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca4, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca5, value : 32'h20a84308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca6, value : 32'h810005c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca7, value : 32'hc0427104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca8, value : 32'hc001c402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ca9, value : 32'hc0416098},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50caa, value : 32'h236fa160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cab, value : 32'h8100003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cac, value : 32'h210b0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cad, value : 32'hc002718d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cae, value : 32'ha1004409},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50caf, value : 32'h74247464},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb0, value : 32'h240a4089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb1, value : 32'h20a872c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb2, value : 32'h82000340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb3, value : 32'hc102c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb4, value : 32'h7822c001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb5, value : 32'hc002c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb6, value : 32'h1a047704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb7, value : 32'hec0d0010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb8, value : 32'h30a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cb9, value : 32'hc220001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cba, value : 32'hd80a00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cbb, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cbc, value : 32'h30b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cbd, value : 32'hc001f00e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cbe, value : 32'hc201e810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cbf, value : 32'h30c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc0, value : 32'hc060001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc1, value : 32'hd80a00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc2, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc3, value : 32'h30d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc4, value : 32'hfe8f0ad6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc5, value : 32'hf009710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc6, value : 32'h30e41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc7, value : 32'hbea0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc8, value : 32'hd80a00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cc9, value : 32'h140c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cca, value : 32'h7ee0341f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ccb, value : 32'hb7c81cf4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ccc, value : 32'h87d4200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ccd, value : 32'h1c040065},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cce, value : 32'h78523001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ccf, value : 32'h6038700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd0, value : 32'hb8224340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd1, value : 32'h71044140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd2, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd3, value : 32'h20a84308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd4, value : 32'h810005c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd5, value : 32'hc0427104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd6, value : 32'hc001c402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd7, value : 32'hc0416098},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd8, value : 32'h236fa160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cd9, value : 32'h8100003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cda, value : 32'h210b0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cdb, value : 32'hc002718d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cdc, value : 32'ha1004409},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cdd, value : 32'h74247464},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cde, value : 32'h240a4089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cdf, value : 32'h20a872c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce0, value : 32'h82000340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce1, value : 32'hc102c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce2, value : 32'h7822c001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce3, value : 32'hc002c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce4, value : 32'h1a047704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce5, value : 32'hec0c0010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce6, value : 32'h30f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce7, value : 32'hb6a0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce8, value : 32'hd80a00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ce9, value : 32'h700cd931},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cea, value : 32'hf00fb914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ceb, value : 32'he811c001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cec, value : 32'h41c3c201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ced, value : 32'h10311},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cee, value : 32'he00b4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cef, value : 32'h700cd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf0, value : 32'h31241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf1, value : 32'ha220000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf2, value : 32'h710cfe8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf3, value : 32'h41c3f008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf4, value : 32'h313},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf5, value : 32'he00b32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf6, value : 32'h700cd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf7, value : 32'h341f140c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf8, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cf9, value : 32'he18f714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cfa, value : 32'hfc7238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cfb, value : 32'h22ca7a38},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cfc, value : 32'hb80e00c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cfd, value : 32'hf812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cfe, value : 32'h2ec9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50cff, value : 32'h240224f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d00, value : 32'h51900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d01, value : 32'hb100b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d02, value : 32'h7fe0b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d03, value : 32'h51900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d04, value : 32'h7fe0720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d05, value : 32'hc420ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d06, value : 32'h2482c3ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d07, value : 32'h41303204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d08, value : 32'h740c4210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d09, value : 32'h21341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d0a, value : 32'h45880000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d0b, value : 32'hada4668},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d0c, value : 32'h474800e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d0d, value : 32'h3605120d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d0e, value : 32'h120c740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d0f, value : 32'h41c33604},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d10, value : 32'h40214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d11, value : 32'h3603120e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d12, value : 32'he00abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d13, value : 32'h3082120d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d14, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d15, value : 32'ha8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d16, value : 32'h7e0815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d17, value : 32'h41c3d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d18, value : 32'h20215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d19, value : 32'haa242c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d1a, value : 32'h43a100e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d1b, value : 32'h24407752},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d1c, value : 32'h27cc3010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d1d, value : 32'hf2039442},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d1e, value : 32'ha5640f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d1f, value : 32'h701407c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d20, value : 32'h7ec0706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d21, value : 32'h1fc7208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d22, value : 32'h9fc0234c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d23, value : 32'h2d006c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d24, value : 32'he0bf78d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d25, value : 32'h2d0052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d26, value : 32'h22c12215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d27, value : 32'hec259181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d28, value : 32'h211578ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d29, value : 32'h90612000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d2a, value : 32'h9000eb1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d2b, value : 32'h994078a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d2c, value : 32'h2048780e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d2d, value : 32'h79100000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d2e, value : 32'h20157230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d2f, value : 32'h20ca22c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d30, value : 32'h4bb2008a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d31, value : 32'h7b8e7a4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d32, value : 32'hfc72289},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d33, value : 32'h2209b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d34, value : 32'h781000c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d35, value : 32'h7a50b141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d36, value : 32'ha4081b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d37, value : 32'h1902d8ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d38, value : 32'hb1000005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d39, value : 32'h2015f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d3a, value : 32'h180222c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d3b, value : 32'h18000005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d3c, value : 32'h71650204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d3d, value : 32'hf1ca71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d3e, value : 32'ha3c0200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d3f, value : 32'h7001248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d40, value : 32'h2a220e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d41, value : 32'h25001002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d42, value : 32'h10141f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d43, value : 32'h25001002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d44, value : 32'h10141f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d45, value : 32'hc7cc700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d46, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d47, value : 32'hc1a8b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d48, value : 32'h31401c04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d49, value : 32'h41c34520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d4a, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d4b, value : 32'h42504078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d4c, value : 32'h42201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d4d, value : 32'hc0177b3b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d4e, value : 32'h9b2d41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d4f, value : 32'h1c1c786c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d50, value : 32'h44c33100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d51, value : 32'h1a448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d52, value : 32'h962440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d53, value : 32'h31c01c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d54, value : 32'h31801c14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d55, value : 32'h972000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d56, value : 32'h30191460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d57, value : 32'h25802700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d58, value : 32'hc000c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d59, value : 32'hd8406849},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d5a, value : 32'h952801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d5b, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d5c, value : 32'h10b7122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d5d, value : 32'h43500081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d5e, value : 32'h861000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d5f, value : 32'h8821c143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d60, value : 32'h222fc144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d61, value : 32'hc0040187},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d62, value : 32'h1dc7210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d63, value : 32'hc003000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d64, value : 32'h80802011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d65, value : 32'h221ff2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d66, value : 32'hf90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d67, value : 32'h225f0a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d68, value : 32'hc0020281},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d69, value : 32'h29e265e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d6a, value : 32'h2700700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d6b, value : 32'h20002414},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d6c, value : 32'hc0012010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d6d, value : 32'h21112400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d6e, value : 32'hc0467834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d6f, value : 32'h9240204c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d70, value : 32'h2d01a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d71, value : 32'h3787272f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d72, value : 32'h702d700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d73, value : 32'h702c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d74, value : 32'h436870cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d75, value : 32'hf005262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d76, value : 32'h800043c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d77, value : 32'h44c44c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d78, value : 32'h44eb0024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d79, value : 32'h100e249f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d7a, value : 32'h92b641c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d7b, value : 32'h646b1030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d7c, value : 32'h68a9eb95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d7d, value : 32'h12c7242f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d7e, value : 32'h4b977baf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d7f, value : 32'h7bcf7c2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d80, value : 32'h7b7b7b82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d81, value : 32'h3e50b17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d82, value : 32'h706c702d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d83, value : 32'h46a94161},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d84, value : 32'heb05f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d85, value : 32'h4300712d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d86, value : 32'h4361f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d87, value : 32'hf1db7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d88, value : 32'h1030091f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d89, value : 32'h7ecf782f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d8a, value : 32'h12c7242f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d8b, value : 32'h7e02dd7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d8c, value : 32'h7edb7d82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d8d, value : 32'h20ca75d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d8e, value : 32'h21ca030d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d8f, value : 32'h70a202cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d90, value : 32'h8002208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d91, value : 32'h41a2f784},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d92, value : 32'hfc12187},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d93, value : 32'h7d2f4709},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d94, value : 32'h1184279a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d95, value : 32'h7d0ac000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d96, value : 32'h308021f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d97, value : 32'h7782702d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d98, value : 32'h3cc2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d99, value : 32'h1c8060b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d9a, value : 32'hc005101c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d9b, value : 32'h248ae824},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d9c, value : 32'h27007001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d9d, value : 32'h80001f8b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d9e, value : 32'h20a81b48},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50d9f, value : 32'h40e30740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da0, value : 32'h14cc2901},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da1, value : 32'he209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da2, value : 32'h7c8f643c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da3, value : 32'h609845a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da4, value : 32'hb8816068},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da5, value : 32'h700c7314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da6, value : 32'h40a0f203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da7, value : 32'h271570ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da8, value : 32'h7125124c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50da9, value : 32'h110e2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50daa, value : 32'hb60074c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dab, value : 32'h1b00b4a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dac, value : 32'hf05016c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dad, value : 32'h7001248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dae, value : 32'h400270a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50daf, value : 32'h1440230a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db0, value : 32'h20120a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db1, value : 32'h290145eb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db2, value : 32'h259f14c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db3, value : 32'h6038100e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db4, value : 32'h708d7f0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db5, value : 32'h606e65f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db6, value : 32'hee2540a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db7, value : 32'h1180275f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db8, value : 32'h40c3651d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50db9, value : 32'hc14c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dba, value : 32'h10b00e11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dbb, value : 32'he1760bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dbc, value : 32'h444a1071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dbd, value : 32'hf0176510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dbe, value : 32'h94816510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dbf, value : 32'h160c2402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc0, value : 32'h60bef011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc1, value : 32'h96816515},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc2, value : 32'h160c2402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc3, value : 32'h7f104cb0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc4, value : 32'h22029602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc5, value : 32'h7ed0200e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc6, value : 32'h20ca76f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc7, value : 32'h24ca034e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc8, value : 32'h7d90148d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dc9, value : 32'h10040d23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dca, value : 32'hed07c507},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dcb, value : 32'h25f4c506},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dcc, value : 32'h60b8120d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dcd, value : 32'h7e1064bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dce, value : 32'h7dc27d90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dcf, value : 32'hd0b71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd0, value : 32'h708d1155},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd1, value : 32'h1b0440a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd2, value : 32'h71251014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd3, value : 32'h3141f04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd4, value : 32'h21842180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd5, value : 32'h21842080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd6, value : 32'h26407105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd7, value : 32'hf130305e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd8, value : 32'hf11171c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dd9, value : 32'h1404c0a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dda, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ddb, value : 32'h4130c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ddc, value : 32'hffef0ae6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ddd, value : 32'hd154508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dde, value : 32'h401011f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ddf, value : 32'h203278ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de0, value : 32'h80000f89},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de1, value : 32'hf00a0d88},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de2, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de3, value : 32'h10086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de4, value : 32'hfe6f0e56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de5, value : 32'h702d42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de6, value : 32'h900446cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de7, value : 32'h6d0a02d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de8, value : 32'h1750821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50de9, value : 32'h294096e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dea, value : 32'h27041289},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50deb, value : 32'h1f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dec, value : 32'h2005c3ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ded, value : 32'h1e000240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dee, value : 32'h90077004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50def, value : 32'hc6cafed4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df0, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df1, value : 32'h10b7122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df2, value : 32'h21540086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df3, value : 32'h88612f08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df4, value : 32'h240b2140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df5, value : 32'h45cb8880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df6, value : 32'h9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df7, value : 32'h36071209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df8, value : 32'h83040bdf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50df9, value : 32'h32e0e59},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dfa, value : 32'h13042c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dfb, value : 32'h7240244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dfc, value : 32'h20a870ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dfd, value : 32'h25050980},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dfe, value : 32'h20050100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50dff, value : 32'h220501c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e00, value : 32'hb90202c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e01, value : 32'h912079a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e02, value : 32'h20300817},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e03, value : 32'h2205b927},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e04, value : 32'hba020202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e05, value : 32'h92407aa5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e06, value : 32'h182226d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e07, value : 32'hb9e06159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e08, value : 32'h21c74121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e09, value : 32'hb90a03e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e0a, value : 32'h1f8f2704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e0b, value : 32'hc3ffffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e0c, value : 32'h2556b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e0d, value : 32'h7f250805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e0e, value : 32'hb0e078c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e0f, value : 32'hf1d27185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e10, value : 32'h226fc2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e11, value : 32'h44cb0443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e12, value : 32'h4988000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e13, value : 32'h8a6084a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e14, value : 32'h7d6c8406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e15, value : 32'h1231c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e16, value : 32'h810212fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e17, value : 32'h231a61b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e18, value : 32'h219a000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e19, value : 32'h40a1041f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e1a, value : 32'h141f259a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e1b, value : 32'h41f209c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e1c, value : 32'h61197bbd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e1d, value : 32'h20798c10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e1e, value : 32'h2447004c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e1f, value : 32'h799817c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e20, value : 32'h2b01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e21, value : 32'h7905706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e22, value : 32'hfe6f0a3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e23, value : 32'h13002d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e24, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e25, value : 32'hc1a1c3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e26, value : 32'hf2315},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e27, value : 32'h260a4008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e28, value : 32'h97013080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e29, value : 32'h703070ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e2a, value : 32'h2e0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e2b, value : 32'h97204328},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e2c, value : 32'h21cc7171},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e2d, value : 32'h1148005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e2e, value : 32'h2b400026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e2f, value : 32'h258a1407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e30, value : 32'h27050fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e31, value : 32'h772d0207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e32, value : 32'h334e2616},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e33, value : 32'h9e609e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e34, value : 32'he2082b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e35, value : 32'h240260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e36, value : 32'h7a7079af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e37, value : 32'h40e07b10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e38, value : 32'he00b3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e39, value : 32'h30c42440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e3a, value : 32'h210c4600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e3b, value : 32'h14039000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e3c, value : 32'h26ca3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e3d, value : 32'h25090245},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e3e, value : 32'h9e030005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e3f, value : 32'h82d9e62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e40, value : 32'h210a00e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e41, value : 32'h79af1180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e42, value : 32'h7b107a70},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e43, value : 32'hb0e40e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e44, value : 32'h244000e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e45, value : 32'h410830c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e46, value : 32'h8000260c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e47, value : 32'h30801403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e48, value : 32'h118521ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e49, value : 32'h52509},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e4a, value : 32'he5c071a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e4b, value : 32'hffc5079c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e4c, value : 32'h45cb9720},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e4d, value : 32'hffff0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e4e, value : 32'h2c5091b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e4f, value : 32'hb179701},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e50, value : 32'h20021025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e51, value : 32'h7a1002c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e52, value : 32'h10402302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e53, value : 32'h20097810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e54, value : 32'hd840008d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e55, value : 32'h3703121f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e56, value : 32'h2002002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e57, value : 32'h201a780c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e58, value : 32'h204000c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e59, value : 32'h780a1040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e5a, value : 32'h2509786c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e5b, value : 32'h210c0203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e5c, value : 32'h20ca9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e5d, value : 32'h70300245},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e5e, value : 32'h521ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e5f, value : 32'h8208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e60, value : 32'h2c22002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e61, value : 32'h7a4ccc1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e62, value : 32'h71507a0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e63, value : 32'h4522ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e64, value : 32'h1fc1204e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e65, value : 32'h2309792f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e66, value : 32'h16000043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e67, value : 32'h80007081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e68, value : 32'hb9e0000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e69, value : 32'hf409705c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e6a, value : 32'h10412340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e6b, value : 32'h782c792c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e6c, value : 32'h20ca7210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e6d, value : 32'h41c30085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e6e, value : 32'hffff00ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e6f, value : 32'h657d7030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e70, value : 32'h521ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e71, value : 32'h7d25b908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e72, value : 32'hc7c640a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e73, value : 32'h1200c0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e74, value : 32'h70ad3087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e75, value : 32'h47cb706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e76, value : 32'h11428000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e77, value : 32'hb69710d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e78, value : 32'h2b4001e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e79, value : 32'h235a0386},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e7a, value : 32'h702d0a0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e7b, value : 32'h704c706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e7c, value : 32'hb0a167d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e7d, value : 32'ha47b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e7e, value : 32'h26050255},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e7f, value : 32'h21050241},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e80, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e81, value : 32'h91200200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e82, value : 32'ha157c2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e83, value : 32'h28000321},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e84, value : 32'h9020130c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e85, value : 32'h81210f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e86, value : 32'hf00db020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e87, value : 32'h71249021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e88, value : 32'hb902b021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e89, value : 32'hf0f2184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e8a, value : 32'h61f961d9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e8b, value : 32'h2c41902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e8c, value : 32'h7425b180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e8d, value : 32'h71447165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e8e, value : 32'h9020f1df},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e8f, value : 32'hb9897164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e90, value : 32'hf1cfb020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e91, value : 32'h78e0c4c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e92, value : 32'hc1a1c3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e93, value : 32'h16004608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e94, value : 32'h80007100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e95, value : 32'h4528000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e96, value : 32'h980206d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e97, value : 32'h817e808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e98, value : 32'h80d0050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e99, value : 32'h1a0000d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e9a, value : 32'hf00700c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e9b, value : 32'h831a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e9c, value : 32'h1a00f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e9d, value : 32'h24400043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e9e, value : 32'h244030c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50e9f, value : 32'hd263081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea0, value : 32'h42c101e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea1, value : 32'hc7c6e802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea2, value : 32'h30821402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea3, value : 32'h308c1403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea4, value : 32'h7b3d6459},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea5, value : 32'h10c12615},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea6, value : 32'h91e0ad60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea7, value : 32'h61f99121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea8, value : 32'hb521793d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ea9, value : 32'h7c3d6399},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eaa, value : 32'h13012615},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eab, value : 32'h91e0ad84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eac, value : 32'h61f99121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ead, value : 32'hb523793d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eae, value : 32'h793d6359},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eaf, value : 32'had287e35},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb0, value : 32'h96219640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb1, value : 32'h793d6159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb2, value : 32'hc7c6b525},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb3, value : 32'hc1a2c3e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb4, value : 32'h45084628},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb5, value : 32'h30011c04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb6, value : 32'hfeaf0fc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb7, value : 32'h30011c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb8, value : 32'hd907d841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eb9, value : 32'hda08b813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eba, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ebb, value : 32'hff670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ebc, value : 32'h70ccfeef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ebd, value : 32'h742c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ebe, value : 32'hff2f0ade},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ebf, value : 32'hc080714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec0, value : 32'ha3641a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec1, value : 32'h734cff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec2, value : 32'h700c4508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec3, value : 32'haca742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec4, value : 32'h714cff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec5, value : 32'hd907706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec6, value : 32'h744c4060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec7, value : 32'h708cb892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec8, value : 32'hfc270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ec9, value : 32'h70ccfeef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eca, value : 32'hd907d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ecb, value : 32'hda08b893},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ecc, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ecd, value : 32'hfae70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ece, value : 32'h70ccfeef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ecf, value : 32'hfe8f0f4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed0, value : 32'hb600b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed1, value : 32'hc7c440a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed2, value : 32'h2044781b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed3, value : 32'hd8e40181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed4, value : 32'h7fe07839},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed5, value : 32'h78e0b8c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed6, value : 32'h1422053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed7, value : 32'h206da941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed8, value : 32'h20ad0182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ed9, value : 32'h605801c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eda, value : 32'ha9007fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50edb, value : 32'h43e3c1a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50edc, value : 32'hffef0fea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50edd, value : 32'hc020c180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ede, value : 32'h30811401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50edf, value : 32'h6038b806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee0, value : 32'h74877b20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee1, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee2, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee3, value : 32'h1cc83a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee4, value : 32'h40383080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee5, value : 32'h30001cc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee6, value : 32'h1cc4700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee7, value : 32'h1cfc3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee8, value : 32'h1cf83000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ee9, value : 32'h1cf43000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eea, value : 32'h1cf03000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eeb, value : 32'h14c83000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eec, value : 32'h1ca03000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eed, value : 32'h20843000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eee, value : 32'h1ca00004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eef, value : 32'h14a03000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef0, value : 32'h1c8c3010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef1, value : 32'h148c30c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef2, value : 32'h1ce03001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef3, value : 32'h28413140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef4, value : 32'h1cac2200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef5, value : 32'h87e3100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef6, value : 32'h401000e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef7, value : 32'h70911600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef8, value : 32'hd8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ef9, value : 32'h30001ce8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50efa, value : 32'h2a00d8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50efb, value : 32'h46084003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50efc, value : 32'h702cc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50efd, value : 32'hb802da50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50efe, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50eff, value : 32'h89038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f00, value : 32'hcfe90e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f01, value : 32'h2456fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f02, value : 32'h148c3800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f03, value : 32'hb8a03000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f04, value : 32'h30001c98},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f05, value : 32'h22002144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f06, value : 32'hd2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f07, value : 32'h30001498},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f08, value : 32'h910811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f09, value : 32'hff8f0e42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f0a, value : 32'h30001cc4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f0b, value : 32'hf004710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f0c, value : 32'hc0085e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f0d, value : 32'h30001cbc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f0e, value : 32'h40037dc4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f0f, value : 32'h2a00d36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f10, value : 32'h33401cd4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f11, value : 32'h30011498},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f12, value : 32'hb1092d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f13, value : 32'h24012144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f14, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f15, value : 32'h148000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f16, value : 32'h4110819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f17, value : 32'h78009fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f18, value : 32'haa6e888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f19, value : 32'h70140780},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f1a, value : 32'h1ca4710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f1b, value : 32'hf40b3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f1c, value : 32'hf007700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f1d, value : 32'h2052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f1e, value : 32'h12178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f1f, value : 32'h1ca47824},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f20, value : 32'h148c3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f21, value : 32'hbfc13000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f22, value : 32'h2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f23, value : 32'h7a009ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f24, value : 32'h30001c9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f25, value : 32'h300214c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f26, value : 32'h24541c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f27, value : 32'h148c0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f28, value : 32'h240a3003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f29, value : 32'h1cd80600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f2a, value : 32'h740c3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f2b, value : 32'h300614ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f2c, value : 32'ha00a56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f2d, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f2e, value : 32'h300014d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f2f, value : 32'h102079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f30, value : 32'h30402042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f31, value : 32'h81b7d0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f32, value : 32'h1cb001f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f33, value : 32'h14b03000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f34, value : 32'hb8c63000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f35, value : 32'h50080b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f36, value : 32'h300014a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f37, value : 32'h1600e88a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f38, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f39, value : 32'hb8e00107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f3a, value : 32'h1c94700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f3b, value : 32'hf2073000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f3c, value : 32'h5400e72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f3d, value : 32'h1c94710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f3e, value : 32'h27793000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f3f, value : 32'hda7d1000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f40, value : 32'h30001cb4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f41, value : 32'h148c708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f42, value : 32'h41db3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f43, value : 32'hc14c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f44, value : 32'h80207c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f45, value : 32'h30001cb8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f46, value : 32'h20402040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f47, value : 32'h30001ccc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f48, value : 32'h3000149c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f49, value : 32'hf80201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f4a, value : 32'h51e00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f4b, value : 32'h30001cec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f4c, value : 32'h800070c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f4d, value : 32'h1cd01b44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f4e, value : 32'h14b03000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f4f, value : 32'hb8c63000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f50, value : 32'h12a01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f51, value : 32'h11c0257c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f52, value : 32'h1ce47824},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f53, value : 32'h2a013000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f54, value : 32'hb8c00340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f55, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f56, value : 32'h1cdc1229},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f57, value : 32'h14983000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f58, value : 32'h20783000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f59, value : 32'h1ca80080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f5a, value : 32'h72963000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f5b, value : 32'h2606de},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f5c, value : 32'hb89fd825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f5d, value : 32'h881b8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f5e, value : 32'h710c7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f5f, value : 32'h5002800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f60, value : 32'h200fb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f61, value : 32'h7e2b050e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f62, value : 32'h2106b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f63, value : 32'hafa730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f64, value : 32'h1d000120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f65, value : 32'h148c1502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f66, value : 32'h24553001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f67, value : 32'h14e03f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f68, value : 32'h24553004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f69, value : 32'h14a43f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f6a, value : 32'h202f3005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f6b, value : 32'h43180507},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f6c, value : 32'h1600bb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f6d, value : 32'h300614d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f6e, value : 32'h300014a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f6f, value : 32'h2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f70, value : 32'h100115bb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f71, value : 32'h30001c90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f72, value : 32'h14904063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f73, value : 32'h81a3002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f74, value : 32'h14900320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f75, value : 32'h14d83003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f76, value : 32'h7fcf3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f77, value : 32'h3003148c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f78, value : 32'h3f052455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f79, value : 32'h30061490},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f7a, value : 32'h14ccc182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f7b, value : 32'h42033007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f7c, value : 32'h91a44e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f7d, value : 32'h43f10060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f7e, value : 32'h300014ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f7f, value : 32'h14a870ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f80, value : 32'hc3823001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f81, value : 32'h300214e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f82, value : 32'h35441c0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f83, value : 32'h2200b0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f84, value : 32'h30431c0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f85, value : 32'h300014a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f86, value : 32'hc809e835},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f87, value : 32'h15b8700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f88, value : 32'h15021086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f89, value : 32'h8de11089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f8a, value : 32'h78ef68d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f8b, value : 32'h10040957},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f8c, value : 32'h2e0e4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f8d, value : 32'h38c2840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f8e, value : 32'h7240244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f8f, value : 32'h70ec7cc5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f90, value : 32'h20a8706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f91, value : 32'h205f0580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f92, value : 32'h24560501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f93, value : 32'h623a3ac2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f94, value : 32'h2812f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f95, value : 32'h22147985},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f96, value : 32'h210501cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f97, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f98, value : 32'h91200320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f99, value : 32'h633b71e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f9a, value : 32'h10441b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f9b, value : 32'h3a812456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f9c, value : 32'h2041a12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f9d, value : 32'h78707914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f9e, value : 32'h2402845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50f9f, value : 32'h71e5b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa0, value : 32'h14b0f1d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa1, value : 32'h8173000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa2, value : 32'h14a801d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa3, value : 32'h14dc3001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa4, value : 32'h20053000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa5, value : 32'hf207807e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa6, value : 32'h1498f00d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa7, value : 32'h8173000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa8, value : 32'h16000090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fa9, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50faa, value : 32'h2044000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fab, value : 32'h2d410815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fac, value : 32'hc972155},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fad, value : 32'hd932011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fae, value : 32'h70ed2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50faf, value : 32'h310b1412},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb0, value : 32'h3108140e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb1, value : 32'h12c02002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb2, value : 32'h31071410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb3, value : 32'h72700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb4, value : 32'h15b8c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb5, value : 32'h15021085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb6, value : 32'h8dc11084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb7, value : 32'h862840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb8, value : 32'hc677bcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fb9, value : 32'hd5f00c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fba, value : 32'h2b4000ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fbb, value : 32'h704c0389},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fbc, value : 32'h11892105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fbd, value : 32'h501235f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fbe, value : 32'h3ac02456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fbf, value : 32'h2750a45},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc0, value : 32'h20146038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc1, value : 32'h2a400081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc2, value : 32'h20050280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc3, value : 32'h20050240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc4, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc5, value : 32'h90000320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc6, value : 32'h2cc2000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc7, value : 32'h1325080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc8, value : 32'h1900b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fc9, value : 32'hf00c01c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fca, value : 32'h710c1600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fcb, value : 32'h13a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fcc, value : 32'h325080b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fcd, value : 32'hb1e07882},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fce, value : 32'hb100f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fcf, value : 32'hf1dc7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd0, value : 32'h71c5b0e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd1, value : 32'h14b8f1ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd2, value : 32'h14b43001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd3, value : 32'h790b3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd4, value : 32'h8de1f231},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd5, value : 32'h8d027eef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd6, value : 32'h384085b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd7, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd8, value : 32'h880012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fd9, value : 32'h3ae084b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fda, value : 32'hbba41c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fdb, value : 32'h14c80620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fdc, value : 32'h43083000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fdd, value : 32'h13002e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fde, value : 32'h244ac107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fdf, value : 32'h79057280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe0, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe1, value : 32'h6872702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe2, value : 32'h4c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe3, value : 32'h106e0b21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe4, value : 32'h38022456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe5, value : 32'h150c265f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe6, value : 32'h2940645c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe7, value : 32'h7a650282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe8, value : 32'hba927c34},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fe9, value : 32'hba9fba9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fea, value : 32'hb4409240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50feb, value : 32'h71e57124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fec, value : 32'hda23f1d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fed, value : 32'hba0a4023},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fee, value : 32'hfe2f0946},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fef, value : 32'h14d8702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff0, value : 32'he8093000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff1, value : 32'h40c3702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff2, value : 32'hbe2c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff3, value : 32'hfe2f0932},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff4, value : 32'h1412daa0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff5, value : 32'h14103112},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff6, value : 32'ha4d310e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff7, value : 32'h210a23a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff8, value : 32'h140d2500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ff9, value : 32'h70143080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ffa, value : 32'h102dc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ffb, value : 32'h108b15b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ffc, value : 32'h8d218d42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ffd, value : 32'h31031410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50ffe, value : 32'h7050782f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h50fff, value : 32'hd03b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51000, value : 32'h102e0b21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51001, value : 32'h7240244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51002, value : 32'hf80201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51003, value : 32'ha3c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51004, value : 32'h20020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51005, value : 32'h300c14d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51006, value : 32'h2080641c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51007, value : 32'hb4600184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51008, value : 32'hf1ec7124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51009, value : 32'h31171414},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5100a, value : 32'h20162479},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5100b, value : 32'h2e812185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5100c, value : 32'h2a162640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5100d, value : 32'h900740d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5100e, value : 32'h14acc29c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5100f, value : 32'h89d3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51010, value : 32'h14980010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51011, value : 32'h8133000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51012, value : 32'h79cf00b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51013, value : 32'h8d64063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51014, value : 32'h734cfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51015, value : 32'hc809f042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51016, value : 32'h108815b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51017, value : 32'h108b1502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51018, value : 32'h8d016852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51019, value : 32'hb51790f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5101a, value : 32'h8491044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5101b, value : 32'h2940106e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5101c, value : 32'hd37038c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5101d, value : 32'h7c452030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5101e, value : 32'h501215f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5101f, value : 32'h3ac32456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51020, value : 32'h7240244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51021, value : 32'h633b702d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51022, value : 32'h38020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51023, value : 32'h12812940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51024, value : 32'h24f23f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51025, value : 32'h67df7985},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51026, value : 32'h21057125},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51027, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51028, value : 32'hb1e00320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51029, value : 32'h2405f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5102a, value : 32'h90041f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5102b, value : 32'hb1c03f20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5102c, value : 32'hf1da7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5102d, value : 32'h440c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5102e, value : 32'heda93e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5102f, value : 32'h702c03e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51030, value : 32'h300114b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51031, value : 32'h300014b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51032, value : 32'hf208790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51033, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51034, value : 32'h1d8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51035, value : 32'hf4d0b8e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51036, value : 32'h1c0ac809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51037, value : 32'hb8023384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51038, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51039, value : 32'hc0049007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5103a, value : 32'h51800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5103b, value : 32'h7014c022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5103c, value : 32'hf217c082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5103d, value : 32'h3101140e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5103e, value : 32'h3f032455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5103f, value : 32'h30051490},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51040, value : 32'h3f842455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51041, value : 32'h300614a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51042, value : 32'hc1404263},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51043, value : 32'h3001148c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51044, value : 32'h4003c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51045, value : 32'h2200d46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51046, value : 32'h3007149c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51047, value : 32'h148cf012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51048, value : 32'h24553001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51049, value : 32'h14c03f05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5104a, value : 32'h704c3003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5104b, value : 32'h300414bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5104c, value : 32'h30061490},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5104d, value : 32'h30071494},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5104e, value : 32'h9b6c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5104f, value : 32'h40030060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51050, value : 32'h300014c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51051, value : 32'hf2917014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51052, value : 32'h30001494},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51053, value : 32'ha147014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51054, value : 32'h1c1c0561},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51055, value : 32'h710c3580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51056, value : 32'he00fda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51057, value : 32'h40034162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51058, value : 32'hfb24162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51059, value : 32'h704c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5105a, value : 32'h8c1c022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5105b, value : 32'hc0820030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5105c, value : 32'h24051800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5105d, value : 32'he81cca00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5105e, value : 32'h2940702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5105f, value : 32'h228a0380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51060, value : 32'h20050004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51061, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51062, value : 32'hb04002f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51063, value : 32'h7200244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51064, value : 32'h10228a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51065, value : 32'h20020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51066, value : 32'h832005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51067, value : 32'h102280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51068, value : 32'h51b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51069, value : 32'hca007124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5106a, value : 32'h800409d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5106b, value : 32'h3101140e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5106c, value : 32'h1490c082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5106d, value : 32'h24553005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5106e, value : 32'h14a83f03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5106f, value : 32'h24553006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51070, value : 32'h149c3f84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51071, value : 32'h42633007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51072, value : 32'h4003c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51073, value : 32'hc8ec140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51074, value : 32'h732c0220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51075, value : 32'h43c3702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51076, value : 32'h4fa88001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51077, value : 32'h945ca00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51078, value : 32'h29400025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51079, value : 32'h700d038b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5107a, value : 32'h833700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5107b, value : 32'h71ed0255},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5107c, value : 32'h30021494},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5107d, value : 32'h70547f18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5107e, value : 32'h900442c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5107f, value : 32'hf20702f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51080, value : 32'hbc0a630c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51081, value : 32'h12cc2405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51082, value : 32'h2305f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51083, value : 32'h7a85120c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51084, value : 32'h10102080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51085, value : 32'h7104b2e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51086, value : 32'he309f1e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51087, value : 32'hf1e07124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51088, value : 32'h1800d820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51089, value : 32'hf0102004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5108a, value : 32'h300314c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5108b, value : 32'h300414bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5108c, value : 32'h3f052455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5108d, value : 32'h4003c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5108e, value : 32'h704c732c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5108f, value : 32'h8b270cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51090, value : 32'h71ec0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51091, value : 32'h30001494},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51092, value : 32'hda47014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51093, value : 32'h14e80581},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51094, value : 32'h40033002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51095, value : 32'h200ebe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51096, value : 32'h700c4162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51097, value : 32'he00ed6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51098, value : 32'h1c1c4162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51099, value : 32'h76e23440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5109a, value : 32'h705278d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5109b, value : 32'hffce05ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5109c, value : 32'hffcf0573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5109d, value : 32'h108b15b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5109e, value : 32'h8d827fd0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5109f, value : 32'h796f8d61},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a0, value : 32'h6587191},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a1, value : 32'hb3dffcd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a2, value : 32'h2456106e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a3, value : 32'h20f43a80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a4, value : 32'h16000042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a5, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a6, value : 32'h6058011b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a7, value : 32'hd81170f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a8, value : 32'h1600f7ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510a9, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510aa, value : 32'h4a10011c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ab, value : 32'hd89170f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ac, value : 32'h6b20ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ad, value : 32'h2105b90e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ae, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510af, value : 32'hb1003ed4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b0, value : 32'hf1df7164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b1, value : 32'h8c1c022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b2, value : 32'h140e0030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b3, value : 32'h8de13113},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b4, value : 32'h8d0279ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b5, value : 32'h6408df},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b6, value : 32'h40c34030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b7, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b8, value : 32'h8a18800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510b9, value : 32'h70cd042e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ba, value : 32'h1291275e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510bb, value : 32'h447202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510bc, value : 32'h1a00d16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510bd, value : 32'h205f4210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510be, value : 32'h14cc2502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510bf, value : 32'hc182300c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c0, value : 32'h248a7c09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c1, value : 32'h623a7001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c2, value : 32'h923a7ad4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c3, value : 32'h41c3643c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c4, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c5, value : 32'h2043241a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c6, value : 32'h201fb922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c7, value : 32'h14ec2041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c8, value : 32'h627a3002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510c9, value : 32'h41c1623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ca, value : 32'h184219a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510cb, value : 32'h2300623b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510cc, value : 32'h80000f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510cd, value : 32'h43681b44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ce, value : 32'h708db180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510cf, value : 32'h78020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d0, value : 32'h300114d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d1, value : 32'h43627a8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d2, value : 32'h62197a39},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d3, value : 32'h218c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d4, value : 32'hf74c8002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d5, value : 32'h215a4242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d6, value : 32'h229f0181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d7, value : 32'h623a000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d8, value : 32'h6432234},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510d9, value : 32'h92417223},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510da, value : 32'h13012315},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510db, value : 32'h71c37185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510dc, value : 32'h1a448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510dd, value : 32'hb141b160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510de, value : 32'he7571c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510df, value : 32'h712692b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e0, value : 32'hf1a871e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e1, value : 32'h3f802455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e2, value : 32'h916a4183},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e3, value : 32'h24569149},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e4, value : 32'hc0413ac5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e5, value : 32'h149c4162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e6, value : 32'h240a3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e7, value : 32'h14cc0540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e8, value : 32'hc0403007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510e9, value : 32'h300014ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ea, value : 32'h62078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510eb, value : 32'hffaf096e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ec, value : 32'h149c4063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ed, value : 32'h40633001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ee, value : 32'h30021490},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ef, value : 32'h1a0093e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f0, value : 32'h300314c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f1, value : 32'h300114b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f2, value : 32'h300014b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f3, value : 32'hf232790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f4, value : 32'h7eef8de1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f5, value : 32'h85d8d02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f6, value : 32'h40c30384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f7, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f8, value : 32'h84d8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510f9, value : 32'h41c103ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510fa, value : 32'h5e00f3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510fb, value : 32'h300014c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510fc, value : 32'h2e404408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510fd, value : 32'hc1071300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510fe, value : 32'h7280244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h510ff, value : 32'hc8097905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51100, value : 32'h700c7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51101, value : 32'h20a86952},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51102, value : 32'hc230500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51103, value : 32'h2456102e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51104, value : 32'h265f3801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51105, value : 32'h61791503},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51106, value : 32'h321f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51107, value : 32'h2812840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51108, value : 32'hb9927945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51109, value : 32'hb99fb99c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5110a, value : 32'h7104b160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5110b, value : 32'hf1d371e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5110c, value : 32'ha9ec082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5110d, value : 32'h702c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5110e, value : 32'h300014d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5110f, value : 32'h20967186},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51110, value : 32'h12b0794},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51111, value : 32'h1cd0ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51112, value : 32'h14943000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51113, value : 32'h70143000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51114, value : 32'h5820b9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51115, value : 32'h3a062480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51116, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51117, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51118, value : 32'h4110c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51119, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5111a, value : 32'h88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5111b, value : 32'h8114548},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5111c, value : 32'h462800b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5111d, value : 32'h2280204a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5111e, value : 32'hf00574ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5111f, value : 32'h2240204a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51120, value : 32'h90272ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51121, value : 32'h208afeef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51122, value : 32'hec1080c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51123, value : 32'h208a1275},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51124, value : 32'h8b90144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51125, value : 32'h923038e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51126, value : 32'h706c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51127, value : 32'hfecf08f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51128, value : 32'hd907706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51129, value : 32'h724c4060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5112a, value : 32'h708cb88f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5112b, value : 32'he3670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5112c, value : 32'h70ccfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5112d, value : 32'hd907f00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5112e, value : 32'hda184060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5112f, value : 32'h708cb88f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51130, value : 32'he2270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51131, value : 32'h70ccfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51132, value : 32'hfecf08c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51133, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51134, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51135, value : 32'h45a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51136, value : 32'hfeaf0e0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51137, value : 32'h704c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51138, value : 32'h4648752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51139, value : 32'hbe94db80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5113a, value : 32'h40c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5113b, value : 32'hdf645a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5113c, value : 32'h70ccfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5113d, value : 32'hd9296e13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5113e, value : 32'h706c42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5113f, value : 32'h45a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51140, value : 32'hfeaf0de2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51141, value : 32'h1c0264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51142, value : 32'h30821204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51143, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51144, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51145, value : 32'hdce45a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51146, value : 32'h70ccfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51147, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51148, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51149, value : 32'h45a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5114a, value : 32'hfeaf0dba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5114b, value : 32'h78db70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5114c, value : 32'h704c752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5114d, value : 32'h4238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5114e, value : 32'h45a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5114f, value : 32'hfeaf0da6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51150, value : 32'hd84170cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51151, value : 32'hf03cd92a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51152, value : 32'h20300921},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51153, value : 32'h842706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51154, value : 32'h706cfecf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51155, value : 32'h4060d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51156, value : 32'hb88f724c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51157, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51158, value : 32'hfeaf0d82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51159, value : 32'hf00d70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5115a, value : 32'h4060d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5115b, value : 32'hb88fda28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5115c, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5115d, value : 32'hfeaf0d6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5115e, value : 32'h81670cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5115f, value : 32'h700cfecf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51160, value : 32'hda08d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51161, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51162, value : 32'hd5a45a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51163, value : 32'h70ccfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51164, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51165, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51166, value : 32'h45a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51167, value : 32'hfeaf0d46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51168, value : 32'h704c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51169, value : 32'h4040752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5116a, value : 32'h4238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5116b, value : 32'h708cb895},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5116c, value : 32'hd3245a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5116d, value : 32'h70ccfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5116e, value : 32'hd92bd841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5116f, value : 32'h42e1b812},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51170, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51171, value : 32'hd1e45a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51172, value : 32'h264afeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51173, value : 32'h700c01c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51174, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51175, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51176, value : 32'hd0a45a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51177, value : 32'h260afeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51178, value : 32'hf960400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51179, value : 32'h700cfe8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5117a, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5117b, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5117c, value : 32'hcf270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5117d, value : 32'h70ccfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5117e, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5117f, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51180, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51181, value : 32'hfeaf0cde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51182, value : 32'hc7e70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51183, value : 32'h7704fe4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51184, value : 32'h78e0c6ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51185, value : 32'h88a0c0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51186, value : 32'h900743c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51187, value : 32'hed07c2cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51188, value : 32'h51b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51189, value : 32'h51b04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5118a, value : 32'h248af005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5118b, value : 32'hb3801fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5118c, value : 32'h1600b382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5118d, value : 32'h80007083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5118e, value : 32'h23780008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5118f, value : 32'h6b920103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51190, value : 32'h900743c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51191, value : 32'hed16c2c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51192, value : 32'h1b04b380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51193, value : 32'h9130085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51194, value : 32'hdb1000f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51195, value : 32'h26f47b2d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51196, value : 32'h800070c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51197, value : 32'h908810c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51198, value : 32'h23cf7295},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51199, value : 32'h1e000361},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5119a, value : 32'h900770c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5119b, value : 32'hf007c29c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5119c, value : 32'h1c0c2445},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5119d, value : 32'h1b04b380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5119e, value : 32'h43c30045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5119f, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a0, value : 32'h8b13b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a1, value : 32'h8bc08be1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a2, value : 32'hf417bcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a3, value : 32'hb3910c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a4, value : 32'h201410ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a5, value : 32'h91300cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a6, value : 32'hdd0a0070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a7, value : 32'h1c24e988},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a8, value : 32'h75ad1285},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511a9, value : 32'h1c24f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511aa, value : 32'hf0051145},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ab, value : 32'h1c24dd0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ac, value : 32'h9151005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ad, value : 32'h221400b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ae, value : 32'h130000c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511af, value : 32'hb0900c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b0, value : 32'hb4b20013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b1, value : 32'hf1e271c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b2, value : 32'h78e0c4c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b3, value : 32'h702cc0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b4, value : 32'h900742c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b5, value : 32'h1e00c2c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b6, value : 32'h90077044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b7, value : 32'hb220fed4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b8, value : 32'h1e00b222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511b9, value : 32'h90087044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ba, value : 32'h800801e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511bb, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511bc, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511bd, value : 32'hb020c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511be, value : 32'h2009e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511bf, value : 32'h80441adc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c0, value : 32'h1800b6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c1, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c2, value : 32'h46c8c2f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c3, value : 32'h47084528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c4, value : 32'h416040c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c5, value : 32'h21c0250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c6, value : 32'h2140220a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c7, value : 32'h2100200a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c8, value : 32'hd324170},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511c9, value : 32'h43500060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ca, value : 32'h40e14410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511cb, value : 32'h704c41a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511cc, value : 32'h240a4322},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511cd, value : 32'h250a0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ce, value : 32'h46c10480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511cf, value : 32'h20085e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d0, value : 32'h540270a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d1, value : 32'hef0870cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d2, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d3, value : 32'hed2ffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d4, value : 32'h712c05a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d5, value : 32'h4102d840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d6, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d7, value : 32'h1e49008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d8, value : 32'h42828508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511d9, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511da, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511db, value : 32'h1800c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511dc, value : 32'h1e000045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511dd, value : 32'h90077384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511de, value : 32'h99ac29c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511df, value : 32'h40620020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e0, value : 32'h41628d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e1, value : 32'hffef0cde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e2, value : 32'ha5074202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e3, value : 32'h412240a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e4, value : 32'hffef0e86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e5, value : 32'hc6d24242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e6, value : 32'hc1a1c3f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e7, value : 32'hd8314608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e8, value : 32'h4528a108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511e9, value : 32'h210ac809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ea, value : 32'ha9c02180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511eb, value : 32'had24702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ec, value : 32'h2140230a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ed, value : 32'h200aa526},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ee, value : 32'hb8022100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ef, value : 32'h20054270},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f0, value : 32'h90380f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f1, value : 32'h90e00008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f2, value : 32'ha522b521},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f3, value : 32'h7200f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f4, value : 32'h11c41d10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f5, value : 32'h20f00a2b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f6, value : 32'ha31ad05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f7, value : 32'h204b2070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f8, value : 32'ha35a140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511f9, value : 32'h204b20b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511fa, value : 32'ha33a140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511fb, value : 32'h204b2031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511fc, value : 32'hf21da140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511fd, value : 32'h14811d18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511fe, value : 32'h14011d14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h511ff, value : 32'h204bf025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51200, value : 32'hf21aa140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51201, value : 32'hf020d828},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51202, value : 32'h1d18f218},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51203, value : 32'h1d141401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51204, value : 32'hf01b1481},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51205, value : 32'hd87af217},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51206, value : 32'h700cf016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51207, value : 32'h22541c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51208, value : 32'hdc60001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51209, value : 32'h4242fdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5120a, value : 32'h1d18f00f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5120b, value : 32'h1d1414c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5120c, value : 32'hf00b1441},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5120d, value : 32'hf008d829},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5120e, value : 32'h14411d18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5120f, value : 32'h14c11d14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51210, value : 32'hd87bf003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51211, value : 32'ha91a505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51212, value : 32'h275320b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51213, value : 32'hf244907e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51214, value : 32'h10310e85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51215, value : 32'h20112179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51216, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51217, value : 32'h8fc0122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51218, value : 32'h402202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51219, value : 32'h22112140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5121a, value : 32'h20522279},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5121b, value : 32'h542044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5121c, value : 32'h8658f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5121d, value : 32'h40c30384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5121e, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5121f, value : 32'h8558800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51220, value : 32'h7acf03ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51221, value : 32'h41424022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51222, value : 32'h1600dfa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51223, value : 32'hfde4382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51224, value : 32'hc1800160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51225, value : 32'h23802314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51226, value : 32'hc11000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51227, value : 32'hef2c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51228, value : 32'h21bf0320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51229, value : 32'hbea0fff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5122a, value : 32'he80d0040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5122b, value : 32'h30801401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5122c, value : 32'hf789e0c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5122d, value : 32'h3f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5122e, value : 32'h30021c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5122f, value : 32'h7104c020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51230, value : 32'hc080c060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51231, value : 32'h200ef6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51232, value : 32'h13902514},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51233, value : 32'h2004182c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51234, value : 32'hf1d071c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51235, value : 32'h78e0c7d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51236, value : 32'h42c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51237, value : 32'h901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51238, value : 32'h900741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51239, value : 32'hb200f800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5123a, value : 32'h151984},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5123b, value : 32'h41a44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5123c, value : 32'h80151980},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5123d, value : 32'h191cb202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5123e, value : 32'h19040015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5123f, value : 32'h19040015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51240, value : 32'h19080015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51241, value : 32'hb1000015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51242, value : 32'h7fe0b102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51243, value : 32'h78e0b104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51244, value : 32'h4050c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51245, value : 32'h82d4130},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51246, value : 32'h45080275},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51247, value : 32'h46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51248, value : 32'h2025ffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51249, value : 32'hf0310340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5124a, value : 32'hf008f015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5124b, value : 32'hf006f016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5124c, value : 32'hf01cf018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5124d, value : 32'hf026f01e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5124e, value : 32'h46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5124f, value : 32'hf025a536},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51250, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51251, value : 32'h10224},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51252, value : 32'hfdef0c9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51253, value : 32'h70cd42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51254, value : 32'hdefff01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51255, value : 32'hf019be08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51256, value : 32'h46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51257, value : 32'hf015aaaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51258, value : 32'h46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51259, value : 32'hf011b2b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5125a, value : 32'h46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5125b, value : 32'hf00d8241},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5125c, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5125d, value : 32'h88c10104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5125e, value : 32'hbe088820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5125f, value : 32'hf0057e25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51260, value : 32'h46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51261, value : 32'h70165a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51262, value : 32'hcc2dfaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51263, value : 32'h27ca0720},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51264, value : 32'he8061021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51265, value : 32'h708f1600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51266, value : 32'h1068000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51267, value : 32'h8e96d0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51268, value : 32'h26040155},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51269, value : 32'h1f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5126a, value : 32'hb928ff00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5126b, value : 32'h42e178cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5126c, value : 32'he2a43e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5126d, value : 32'h240a05a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5126e, value : 32'h16000440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5126f, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51270, value : 32'h72140008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51271, value : 32'h901c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51272, value : 32'h40c30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51273, value : 32'hf8009007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51274, value : 32'h1900f406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51275, value : 32'h18000005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51276, value : 32'hf0060005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51277, value : 32'h451900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51278, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51279, value : 32'h12300da7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5127a, value : 32'hd59d8ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5127b, value : 32'hd551110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5127c, value : 32'hdf111d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5127d, value : 32'hd9441031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5127e, value : 32'h901c40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5127f, value : 32'h45cb0044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51280, value : 32'hf8849007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51281, value : 32'h851800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51282, value : 32'h90951d80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51283, value : 32'h804418c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51284, value : 32'h94e4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51285, value : 32'h1d0005e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51286, value : 32'h700c1105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51287, value : 32'h901f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51288, value : 32'h7ad0c00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51289, value : 32'hb518b516},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5128a, value : 32'hb51a4340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5128b, value : 32'hb1004440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5128c, value : 32'hb1024540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5128d, value : 32'hb504712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5128e, value : 32'h2200bde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5128f, value : 32'hc6cab506},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51290, value : 32'h900745cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51291, value : 32'h1d04f830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51292, value : 32'h704c13d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51293, value : 32'hfc7208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51294, value : 32'h388242f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51295, value : 32'h722cb540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51296, value : 32'h700cb502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51297, value : 32'h250a706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51298, value : 32'hbb60100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51299, value : 32'h47480220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5129a, value : 32'h1c012542},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5129b, value : 32'h901f40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5129c, value : 32'h1900c00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5129d, value : 32'h1d500085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5129e, value : 32'hb0e013c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5129f, value : 32'hb1e4b0e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a0, value : 32'hc6cab1e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a1, value : 32'h90500d1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a2, value : 32'h45cbf199},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a3, value : 32'hf8209007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a4, value : 32'h13d41d04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a5, value : 32'h10151d04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a6, value : 32'h1d08700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a7, value : 32'h7ad01014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a8, value : 32'h13d41d04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512a9, value : 32'h901f47cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512aa, value : 32'h1d00c004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ab, value : 32'h25421404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ac, value : 32'hb5021c11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ad, value : 32'hb700d844},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ae, value : 32'h722c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512af, value : 32'h44404340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b0, value : 32'hb564540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b1, value : 32'h19000220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b2, value : 32'h1d502105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b3, value : 32'h1f081404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b4, value : 32'h1f0c1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b5, value : 32'h19081404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b6, value : 32'h190c2404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b7, value : 32'hc6ca2404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b8, value : 32'h70051e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512b9, value : 32'hf8049007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ba, value : 32'h78e0c6ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512bb, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512bc, value : 32'hc1bfb6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512bd, value : 32'h47084338},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512be, value : 32'hc08b70ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512bf, value : 32'hda50702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c0, value : 32'h31c01c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c1, value : 32'h2140200a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c2, value : 32'h31801c08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c3, value : 32'h31001c04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c4, value : 32'h1c28c348},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c5, value : 32'hdea3580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c6, value : 32'h1c24fdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c7, value : 32'hc8093580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c8, value : 32'h308d237c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512c9, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ca, value : 32'h90380f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512cb, value : 32'h90000008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512cc, value : 32'h2079b8c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512cd, value : 32'h6f0b000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ce, value : 32'h39c7514},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512cf, value : 32'h71f50026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d0, value : 32'h400962},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d1, value : 32'h25044610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d2, value : 32'hb0f1395},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d3, value : 32'h712f3070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d4, value : 32'h21ca70d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d5, value : 32'h47cb3541},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d6, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d7, value : 32'h25802504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d8, value : 32'h300e14b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512d9, value : 32'h71148f60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512da, value : 32'h202f8f41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512db, value : 32'h223c058a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512dc, value : 32'h25ca00c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512dd, value : 32'h78252021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512de, value : 32'h3f081b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512df, value : 32'h40614368},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e0, value : 32'h7104790f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e1, value : 32'h10412614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e2, value : 32'h51924},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e3, value : 32'haf5790f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e4, value : 32'h23788045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e5, value : 32'h737730c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e6, value : 32'h1618e009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e7, value : 32'hc0431017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e8, value : 32'hc044700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512e9, value : 32'h26120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ea, value : 32'h8605c044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512eb, value : 32'h9608c045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ec, value : 32'h30300969},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ed, value : 32'hc809c047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ee, value : 32'h12c0200a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ef, value : 32'h108717b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f0, value : 32'h5c02005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f1, value : 32'h10861701},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f2, value : 32'h212f6892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f3, value : 32'he4d0207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f4, value : 32'hf450044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f5, value : 32'h2940006e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f6, value : 32'h215f0383},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f7, value : 32'h7b850289},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f8, value : 32'hc203700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512f9, value : 32'h850831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512fa, value : 32'hea88c202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512fb, value : 32'h6822100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512fc, value : 32'h821220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512fd, value : 32'h80081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512fe, value : 32'h2422000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h512ff, value : 32'h7d54c58b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51300, value : 32'h2822840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51301, value : 32'hba927a65},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51302, value : 32'hba9fba9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51303, value : 32'hb5409240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51304, value : 32'hf1e97104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51305, value : 32'hf1db7105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51306, value : 32'h40cb7377},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51307, value : 32'hf000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51308, value : 32'h20002552},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51309, value : 32'h102120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5130a, value : 32'h800040db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5130b, value : 32'hc04612e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5130c, value : 32'h2c7222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5130d, value : 32'h8678f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5130e, value : 32'h10000084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5130f, value : 32'h85b3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51310, value : 32'h2a4000ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51311, value : 32'hc0050303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51312, value : 32'h2012305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51313, value : 32'h900444cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51314, value : 32'h79050000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51315, value : 32'h7905c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51316, value : 32'h208d20f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51317, value : 32'h7985b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51318, value : 32'hc106b1a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51319, value : 32'hb040210b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5131a, value : 32'h2305f20b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5131b, value : 32'h210505c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5131c, value : 32'h78250201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5131d, value : 32'h7c05b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5131e, value : 32'h208020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5131f, value : 32'hd1bb400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51320, value : 32'h26142030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51321, value : 32'h23051080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51322, value : 32'h903605c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51323, value : 32'h208020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51324, value : 32'hfeef0b72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51325, value : 32'h7165c201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51326, value : 32'hf0ef1cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51327, value : 32'h8f610500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51328, value : 32'hb458f20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51329, value : 32'h7a2f0044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5132a, value : 32'h2a407124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5132b, value : 32'h2614038b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5132c, value : 32'h2305108c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5132d, value : 32'h90041f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5132e, value : 32'h900002d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5132f, value : 32'h20849492},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51330, value : 32'hbc0a040e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51331, value : 32'h204f7885},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51332, value : 32'h2305000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51333, value : 32'h90041f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51334, value : 32'hb0803ed4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51335, value : 32'h7854c089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51336, value : 32'h208220f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51337, value : 32'h782fb040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51338, value : 32'h80050bc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51339, value : 32'hfeaf0a3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5133a, value : 32'ha4ad8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5133b, value : 32'h960efeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5133c, value : 32'h248a702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5133d, value : 32'hc0082002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5133e, value : 32'hfe6f0dc2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5133f, value : 32'h1700712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51340, value : 32'h8f211093},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51341, value : 32'h24c7202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51342, value : 32'ha040200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51343, value : 32'h2d0152},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51344, value : 32'hfcf228a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51345, value : 32'h30801000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51346, value : 32'h84002011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51347, value : 32'h2440f29f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51348, value : 32'hc507390b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51349, value : 32'h140123f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5134a, value : 32'h140b2314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5134b, value : 32'h30b50b37},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5134c, value : 32'hb9c6653d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5134d, value : 32'h6038c007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5134e, value : 32'h8002208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5134f, value : 32'h2555f796},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51350, value : 32'hd2d180d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51351, value : 32'h1b002030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51352, value : 32'h26141344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51353, value : 32'hc2011400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51354, value : 32'h23032840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51355, value : 32'h23059036},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51356, value : 32'haaa05c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51357, value : 32'h78b0feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51358, value : 32'h1b00f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51359, value : 32'hf0351344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5135a, value : 32'h13441b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5135b, value : 32'h119e0d63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5135c, value : 32'he82fc001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5135d, value : 32'h180d2554},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5135e, value : 32'h20300d1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5135f, value : 32'h13441b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51360, value : 32'h14002614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51361, value : 32'h23032840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51362, value : 32'h5c32305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51363, value : 32'h9036714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51364, value : 32'hfeef0a72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51365, value : 32'he3b78b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51366, value : 32'h28402031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51367, value : 32'hd90f238c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51368, value : 32'h1f802405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51369, value : 32'h2d49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5136a, value : 32'h26149060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5136b, value : 32'h90521400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5136c, value : 32'hb0327946},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5136d, value : 32'hf802304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5136e, value : 32'hc3ff0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5136f, value : 32'h7905b90a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51370, value : 32'h1f802405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51371, value : 32'h3ed49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51372, value : 32'h1300b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51373, value : 32'h2840110d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51374, value : 32'hc8092302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51375, value : 32'hc0057a05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51376, value : 32'h41c37845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51377, value : 32'h3c009004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51378, value : 32'h7825b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51379, value : 32'hc006b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5137a, value : 32'hb000210b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5137b, value : 32'h2205f208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5137c, value : 32'h6a1205c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5137d, value : 32'h13007825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5137e, value : 32'hb0201101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5137f, value : 32'h23802840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51380, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51381, value : 32'h26fc9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51382, value : 32'h1121000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51383, value : 32'hc002c504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51384, value : 32'he88e7aaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51385, value : 32'h2110a09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51386, value : 32'he89cc000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51387, value : 32'he888c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51388, value : 32'h26802000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51389, value : 32'h801020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5138a, value : 32'ha29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5138b, value : 32'he8098e04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5138c, value : 32'h11041602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5138d, value : 32'h447232f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5138e, value : 32'h4102c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5138f, value : 32'hc000f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51390, value : 32'h448242f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51391, value : 32'h706c4102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51392, value : 32'h4600f7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51393, value : 32'h480250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51394, value : 32'hc00371a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51395, value : 32'h9bb79af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51396, value : 32'h71668004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51397, value : 32'h40c3f153},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51398, value : 32'hc2ec9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51399, value : 32'hb0407126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5139a, value : 32'h21fd248d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5139b, value : 32'h51800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5139c, value : 32'h3010095d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5139d, value : 32'h108b17b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5139e, value : 32'h7c4f8f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5139f, value : 32'h3040951},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a0, value : 32'h132e0b49},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a1, value : 32'h13002c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a2, value : 32'h128d245f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a3, value : 32'h5c32005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a4, value : 32'h7865c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a5, value : 32'h68d2706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a6, value : 32'hb31c003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a7, value : 32'hc0020005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a8, value : 32'h2400e887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513a9, value : 32'h10201680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513aa, value : 32'hb1d0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ab, value : 32'h63bf0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ac, value : 32'h20f4c08b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ad, value : 32'h2b4003cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ae, value : 32'h78c50280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513af, value : 32'hb89cb892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b0, value : 32'hb0e0b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b1, value : 32'hf1ea7164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b2, value : 32'hf1d97144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b3, value : 32'h1404c0bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b4, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b5, value : 32'hffc1046c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b6, value : 32'hffcf046f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b7, value : 32'hf812032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b8, value : 32'hea48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513b9, value : 32'h2150809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ba, value : 32'hf0037933},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513bb, value : 32'h7fe0b9c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513bc, value : 32'h78e0782d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513bd, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513be, value : 32'h70c51e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513bf, value : 32'h88900c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c0, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c1, value : 32'hafec0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c2, value : 32'ha3afd8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c3, value : 32'h4608fd8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c4, value : 32'h4528ca09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c5, value : 32'heac7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c6, value : 32'hc1a10321},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c7, value : 32'hc040c086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c8, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513c9, value : 32'h128000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ca, value : 32'h10240e0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513cb, value : 32'hff640a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513cc, value : 32'hc10006e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513cd, value : 32'h7014ca09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ce, value : 32'h6c10cac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513cf, value : 32'hdc247487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d0, value : 32'hfd8f0273},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d1, value : 32'hc1a2c3e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d2, value : 32'h45284050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d3, value : 32'h41c34200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d4, value : 32'h1035e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d5, value : 32'hffef0fb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d6, value : 32'hed23750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d7, value : 32'h70cd704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d8, value : 32'h7100244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513d9, value : 32'h4040702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513da, value : 32'h24020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513db, value : 32'h20f4c380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513dc, value : 32'h7b34200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513dd, value : 32'h712460b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513de, value : 32'h1406b380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513df, value : 32'h750c3106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e0, value : 32'h31041402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e1, value : 32'h35f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e2, value : 32'h14040005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e3, value : 32'hf7a3105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e4, value : 32'h1400ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e5, value : 32'h71c53103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e6, value : 32'hac97ad0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e7, value : 32'hc7c88344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e8, value : 32'h2550a15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513e9, value : 32'h215fe808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ea, value : 32'h621a0240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513eb, value : 32'hf822232},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ec, value : 32'h4fa88001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ed, value : 32'h40407fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ee, value : 32'h88008821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ef, value : 32'h7fe0b807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f0, value : 32'h78e06038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f1, value : 32'h88008821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f2, value : 32'h7fe0b806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f3, value : 32'h78e06038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f4, value : 32'h216c791d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f5, value : 32'h20530142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f6, value : 32'h20840141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f7, value : 32'h60380001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f8, value : 32'h60587fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513f9, value : 32'h432801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513fa, value : 32'h2b007a69},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513fb, value : 32'h78220041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513fc, value : 32'h7fe0621a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513fd, value : 32'h78e07850},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513fe, value : 32'h215fc0e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h513ff, value : 32'h44cb0a03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51400, value : 32'h11428000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51401, value : 32'h647970cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51402, value : 32'h639291a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51403, value : 32'he257a04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51404, value : 32'h23151365},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51405, value : 32'h61990381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51406, value : 32'h790b9122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51407, value : 32'h79dbf208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51408, value : 32'h412314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51409, value : 32'h91236199},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5140a, value : 32'h42220f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5140b, value : 32'hf1f171c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5140c, value : 32'hc4c47850},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5140d, value : 32'hc1a4c3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5140e, value : 32'h1600d9b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5140f, value : 32'h80007093},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51410, value : 32'hb9120004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51411, value : 32'hffef0ec2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51412, value : 32'h45cb740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51413, value : 32'h4e7f8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51414, value : 32'h25546dcb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51415, value : 32'habe1915},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51416, value : 32'h40c10220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51417, value : 32'ha6640c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51418, value : 32'hd90b0560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51419, value : 32'ha5e40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5141a, value : 32'hd9110560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5141b, value : 32'hd91240c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5141c, value : 32'hfeaf0aaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5141d, value : 32'h40c1daef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5141e, value : 32'h5600a4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5141f, value : 32'h40c1d912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51420, value : 32'h5600a42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51421, value : 32'heead929},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51422, value : 32'h40c10520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51423, value : 32'h5200ee2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51424, value : 32'h40c340a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51425, value : 32'h4f128001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51426, value : 32'h5200ed6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51427, value : 32'h40c34210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51428, value : 32'h4f5d8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51429, value : 32'h5200eca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5142a, value : 32'h16034110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5142b, value : 32'h70ed10c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5142c, value : 32'h40d38e36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5142d, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5142e, value : 32'h18b88e4d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5142f, value : 32'h180023c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51430, value : 32'ha1323c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51431, value : 32'h18bc017e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51432, value : 32'h80b2380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51433, value : 32'h9350012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51434, value : 32'h7905011e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51435, value : 32'h1bf092d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51436, value : 32'had00b886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51437, value : 32'h1080154b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51438, value : 32'h1d4bb886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51439, value : 32'h15961002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5143a, value : 32'hb8861080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5143b, value : 32'h10021d96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5143c, value : 32'h108015e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5143d, value : 32'h1de1b886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5143e, value : 32'hb021002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5143f, value : 32'h710c06e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51440, value : 32'h6832c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51441, value : 32'h901c40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51442, value : 32'h79050504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51443, value : 32'h276fb1e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51444, value : 32'h18a410c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51445, value : 32'h41c38045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51446, value : 32'h94007735},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51447, value : 32'h20448f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51448, value : 32'h40c38082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51449, value : 32'h8480001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5144a, value : 32'h25ca4508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5144b, value : 32'h8f381041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5144c, value : 32'h41c3e908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5144d, value : 32'h2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5144e, value : 32'hffef0dce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5144f, value : 32'hf048d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51450, value : 32'h41c37054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51451, value : 32'hc2000beb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51452, value : 32'h4120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51453, value : 32'h3600e46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51454, value : 32'h1600702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51455, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51456, value : 32'h80d000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51457, value : 32'hd84000be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51458, value : 32'h6c00c7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51459, value : 32'hffcf0d96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5145a, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5145b, value : 32'h8820019b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5145c, value : 32'h808010ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5145d, value : 32'h807e2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5145e, value : 32'h782af219},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5145f, value : 32'hf80201a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51460, value : 32'h4240000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51461, value : 32'h3600e32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51462, value : 32'h4200702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51463, value : 32'h21aac80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51464, value : 32'h79120104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51465, value : 32'h850921},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51466, value : 32'h10423aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51467, value : 32'h80c408fd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51468, value : 32'h14420aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51469, value : 32'h7a225033},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5146a, value : 32'h40a1f008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5146b, value : 32'h3600de6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5146c, value : 32'hf00e702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5146d, value : 32'hc80b621a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5146e, value : 32'h10421aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5146f, value : 32'ha5090d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51470, value : 32'h14423aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51471, value : 32'h80c008f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51472, value : 32'h10420aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51473, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51474, value : 32'hd8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51475, value : 32'ha18b8e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51476, value : 32'hc1606c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51477, value : 32'h45cb0380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51478, value : 32'h11408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51479, value : 32'h88d8d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5147a, value : 32'h8f000010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5147b, value : 32'hdf0885},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5147c, value : 32'h800d0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5147d, value : 32'hfe0f08aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5147e, value : 32'h708e8d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5147f, value : 32'he807704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51480, value : 32'h20448f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51481, value : 32'h20780200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51482, value : 32'h700c0002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51483, value : 32'hfe6f0bca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51484, value : 32'h8d01d908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51485, value : 32'hb4081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51486, value : 32'h8d00704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51487, value : 32'h8f00e806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51488, value : 32'h2002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51489, value : 32'h22078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5148a, value : 32'hbae700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5148b, value : 32'h702cfe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5148c, value : 32'h704c8d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5148d, value : 32'h8f00e806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5148e, value : 32'h2002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5148f, value : 32'h22078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51490, value : 32'hb96700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51491, value : 32'hd90afe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51492, value : 32'he8078d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51493, value : 32'h20448f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51494, value : 32'h20780200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51495, value : 32'hd8080014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51496, value : 32'hb7e702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51497, value : 32'h4282fe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51498, value : 32'he80f8d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51499, value : 32'h20448f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5149a, value : 32'h20780200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5149b, value : 32'hf00a0002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5149c, value : 32'h1e40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5149d, value : 32'hd1e8480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5149e, value : 32'h702c0360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5149f, value : 32'h704cf00e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a0, value : 32'hb56700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a1, value : 32'hd996fe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a2, value : 32'h5400ee2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a3, value : 32'h806700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a4, value : 32'h712cfe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a5, value : 32'hc00bfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a6, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a7, value : 32'h2fe8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a8, value : 32'h3e0815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514a9, value : 32'h41c3d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514aa, value : 32'h2e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ab, value : 32'hffcf0c5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ac, value : 32'h7000e32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ad, value : 32'he82c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ae, value : 32'h23530560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514af, value : 32'hc08020d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b0, value : 32'h600ed2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b1, value : 32'h40c1d91c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b2, value : 32'hc280702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b3, value : 32'h708cdbff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b4, value : 32'h7200f0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b5, value : 32'ha5670ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b6, value : 32'he5e0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b7, value : 32'hc0800560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b8, value : 32'heb2c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514b9, value : 32'hd9100060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ba, value : 32'heaac080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514bb, value : 32'hd91c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514bc, value : 32'h712c40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514bd, value : 32'hdbffc280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514be, value : 32'h7200ee2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514bf, value : 32'h40c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c0, value : 32'h4e0094e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c1, value : 32'h40c1d90b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c2, value : 32'h4e00946},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c3, value : 32'h40c1d911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c4, value : 32'h4e0093e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c5, value : 32'h40c1d912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c6, value : 32'h4e00936},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c7, value : 32'hca0ed929},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c8, value : 32'h10050d2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514c9, value : 32'h2b02235f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ca, value : 32'h1f812532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514cb, value : 32'h4788000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514cc, value : 32'h7ab561cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514cd, value : 32'h720271a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ce, value : 32'h2132aa68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514cf, value : 32'haa6a0483},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d0, value : 32'h5432132},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d1, value : 32'h4412132},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d2, value : 32'haa2baa69},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d3, value : 32'hd0af1ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d4, value : 32'hda6efe8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d5, value : 32'h12c5ba9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d6, value : 32'h1a018480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d7, value : 32'h4afb0012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d8, value : 32'h6832240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514d9, value : 32'h4801101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514da, value : 32'h1101aa00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514db, value : 32'h1b010480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514dc, value : 32'h11050012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514dd, value : 32'hab000480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514de, value : 32'h4801101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514df, value : 32'h1101aa01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e0, value : 32'haa020480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e1, value : 32'h4801101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e2, value : 32'h1101ab01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e3, value : 32'hab020480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e4, value : 32'h4801176},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e5, value : 32'h8012198b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e6, value : 32'h4801101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e7, value : 32'h1a794220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e8, value : 32'h1101000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514e9, value : 32'h6a650480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ea, value : 32'h111dab00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514eb, value : 32'hab050480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ec, value : 32'h4801101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ed, value : 32'h21956},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ee, value : 32'h4801101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ef, value : 32'h1101aa01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f0, value : 32'hab010480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f1, value : 32'h4801111},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f2, value : 32'h1101ab06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f3, value : 32'h19430480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f4, value : 32'h89000002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f5, value : 32'h8901aa02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f6, value : 32'h8902ab02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f7, value : 32'hc7d2ab07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f8, value : 32'h40c3c5e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514f9, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514fa, value : 32'h706c88a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514fb, value : 32'h704c8880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514fc, value : 32'hca00702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514fd, value : 32'h50921},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514fe, value : 32'h3040909},
                          '{ step_type : REG_WRITE, reg_addr : 32'h514ff, value : 32'h10450d0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51500, value : 32'hf802205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51501, value : 32'h3ed49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51502, value : 32'h7124b060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51503, value : 32'h72c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51504, value : 32'hf1f14000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51505, value : 32'h78e0c4c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51506, value : 32'h1c00dc3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51507, value : 32'h7c0f0302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51508, value : 32'h80db830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51509, value : 32'h4c3100a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5150a, value : 32'hf00a4852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5150b, value : 32'h250b09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5150c, value : 32'hf0064872},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5150d, value : 32'h704c7831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5150e, value : 32'h21c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5150f, value : 32'hcc1f792c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51510, value : 32'h3211a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51511, value : 32'h221acc1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51512, value : 32'h782c0081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51513, value : 32'h60787fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51514, value : 32'h44cbc0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51515, value : 32'h1078000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51516, value : 32'h42008c60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51517, value : 32'h3f0b2d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51518, value : 32'hb29710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51519, value : 32'h700c007f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5151a, value : 32'h7234b9a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5151b, value : 32'hfec20dcc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5151c, value : 32'h40c3f40b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5151d, value : 32'h4e7f8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5151e, value : 32'h9081145b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5151f, value : 32'h78258800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51520, value : 32'h207a780d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51521, value : 32'h78440000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51522, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51523, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51524, value : 32'h68000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51525, value : 32'hf80203c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51526, value : 32'hc800000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51527, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51528, value : 32'h6c3216f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51529, value : 32'hb8e68900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5152a, value : 32'h7ce0700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5152b, value : 32'h20448907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5152c, value : 32'h7fe00200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5152d, value : 32'h78e0b823},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5152e, value : 32'h4528c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5152f, value : 32'hfdef0de2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51530, value : 32'hee1e4608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51531, value : 32'h5400cca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51532, value : 32'hd925700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51533, value : 32'hdb86704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51534, value : 32'h45a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51535, value : 32'hfe2f0e0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51536, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51537, value : 32'h704cd926},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51538, value : 32'h708cdb86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51539, value : 32'hdfe70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5153a, value : 32'h70ccfe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5153b, value : 32'hd910700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5153c, value : 32'hfe6f08e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5153d, value : 32'hc76714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5153e, value : 32'hf00c0540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5153f, value : 32'h10452553},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51540, value : 32'hd919d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51541, value : 32'hdb86744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51542, value : 32'hdda708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51543, value : 32'h70ccfe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51544, value : 32'hd82700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51545, value : 32'h712cfe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51546, value : 32'h40c3ee87},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51547, value : 32'h75300000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51548, value : 32'h3600a72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51549, value : 32'hc6c4d91e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5154a, value : 32'hb5ec0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5154b, value : 32'h730c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5154c, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5154d, value : 32'h88001140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5154e, value : 32'h1600e810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5154f, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51550, value : 32'h8190001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51551, value : 32'h9b600df},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51552, value : 32'h710c0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51553, value : 32'hffef0f6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51554, value : 32'h942d90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51555, value : 32'hf00600c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51556, value : 32'hf62700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51557, value : 32'hd90fffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51558, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51559, value : 32'h4430c2f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5155a, value : 32'hfeef0cd2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5155b, value : 32'h46cb4110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5155c, value : 32'h12e48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5155d, value : 32'h43108620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5155e, value : 32'h800140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5155f, value : 32'h88e04e7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51560, value : 32'h442202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51561, value : 32'h70901600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51562, value : 32'h628000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51563, value : 32'h704cb8c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51564, value : 32'h856706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51565, value : 32'h42100260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51566, value : 32'h900745cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51567, value : 32'he0ac17c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51568, value : 32'h1d0004e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51569, value : 32'hcfa1005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5156a, value : 32'h708cfdcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5156b, value : 32'h4080752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5156c, value : 32'hb895714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5156d, value : 32'h4238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5156e, value : 32'h440250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5156f, value : 32'hfe2f0d26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51570, value : 32'hd88070cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51571, value : 32'hb892d90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51572, value : 32'h706cda20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51573, value : 32'h500240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51574, value : 32'h440250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51575, value : 32'hfe2f0d0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51576, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51577, value : 32'hfe2f0cb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51578, value : 32'h2705712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51579, value : 32'h78ed140f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5157a, value : 32'h20310b0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5157b, value : 32'h10451d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5157c, value : 32'h120807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5157d, value : 32'h8620c6d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5157e, value : 32'h22084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5157f, value : 32'h1c32841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51580, value : 32'hfe64042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51581, value : 32'h42620220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51582, value : 32'h78e0c6d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51583, value : 32'hb7c81cf4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51584, value : 32'hc181c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51585, value : 32'h1c08714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51586, value : 32'haca3001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51587, value : 32'h1c0404a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51588, value : 32'hd96d3001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51589, value : 32'h8e2750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5158a, value : 32'hb913ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5158b, value : 32'h712c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5158c, value : 32'hffef0916},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5158d, value : 32'h140cc281},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5158e, value : 32'h7ee0341f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5158f, value : 32'hb7c81cf4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51590, value : 32'h70c3c181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51591, value : 32'h400100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51592, value : 32'h1c08714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51593, value : 32'ha963001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51594, value : 32'h1c0404a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51595, value : 32'h41c33001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51596, value : 32'h367},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51597, value : 32'hffef08aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51598, value : 32'h700c750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51599, value : 32'h8e2712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5159a, value : 32'hc281ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5159b, value : 32'h341f140c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5159c, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5159d, value : 32'h4130c2ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5159e, value : 32'h700e4210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5159f, value : 32'h21d508f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a0, value : 32'h203e0a75},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a1, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a2, value : 32'h100e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a3, value : 32'hffef087a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a4, value : 32'h702c4202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a5, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a6, value : 32'h88400485},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a7, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a8, value : 32'h88801228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515a9, value : 32'h7200244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515aa, value : 32'h706c706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ab, value : 32'h4c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ac, value : 32'h209f4081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ad, value : 32'h2100001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ae, value : 32'h2840200d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515af, value : 32'h60b82200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b0, value : 32'h6029615d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b1, value : 32'h11c0234e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b2, value : 32'h29007165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b3, value : 32'h41a10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b4, value : 32'h7a6f7b05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b5, value : 32'he241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b6, value : 32'h82e0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b7, value : 32'h740cffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b8, value : 32'h9004258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515b9, value : 32'hffe507b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ba, value : 32'hd9e341a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515bb, value : 32'h81a740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515bc, value : 32'hb910ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515bd, value : 32'h207e0a75},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515be, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515bf, value : 32'h100e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c0, value : 32'hffef0806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c1, value : 32'h702c4202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c2, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c3, value : 32'h88400485},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c4, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c5, value : 32'h88801228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c6, value : 32'h7200244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c7, value : 32'h706c706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c8, value : 32'h4c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515c9, value : 32'h209f4081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ca, value : 32'h2100001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515cb, value : 32'h2840200d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515cc, value : 32'h60b82200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515cd, value : 32'h6029615d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ce, value : 32'h11c0234e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515cf, value : 32'h29007165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d0, value : 32'h41a10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d1, value : 32'h7a6f7b05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d2, value : 32'he541c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d3, value : 32'hfba0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d4, value : 32'h740cffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d5, value : 32'h9004258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d6, value : 32'hffe507b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d7, value : 32'hd97341a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d8, value : 32'hfa6740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515d9, value : 32'hb911ffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515da, value : 32'hf18a7106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515db, value : 32'h78e0c6cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515dc, value : 32'hc1a2c3f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515dd, value : 32'h46504170},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515de, value : 32'hc1814730},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515df, value : 32'h30c22440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e0, value : 32'h1600af2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e1, value : 32'h30832440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e2, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e3, value : 32'h211a28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e4, value : 32'h14022011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e5, value : 32'h232f3094},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e6, value : 32'h46cb2000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e7, value : 32'h1b448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e8, value : 32'h308d1403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515e9, value : 32'h23640c9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ea, value : 32'hb7a79af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515eb, value : 32'h40e20560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ec, value : 32'h704e4510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ed, value : 32'h24ae0d85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ee, value : 32'h261f474a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ef, value : 32'h251a24c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f0, value : 32'h1f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f1, value : 32'h279a0a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f2, value : 32'h71221184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f3, value : 32'h671f6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f4, value : 32'h6a00efe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f5, value : 32'h13d02600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f6, value : 32'h20851002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f7, value : 32'h13842734},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f8, value : 32'h21061004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515f9, value : 32'h2d41e808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515fa, value : 32'h740c0085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515fb, value : 32'ha641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515fc, value : 32'hf0060005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515fd, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515fe, value : 32'h500a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h515ff, value : 32'hf0a42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51600, value : 32'h4342ffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51601, value : 32'h18002659},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51602, value : 32'h1600671f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51603, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51604, value : 32'h819000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51605, value : 32'h40e1007f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51606, value : 32'h200bca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51607, value : 32'h40e1712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51608, value : 32'h200bc2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51609, value : 32'hf00a702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5160a, value : 32'h90240e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5160b, value : 32'h712c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5160c, value : 32'h8fa40e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5160d, value : 32'h702c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5160e, value : 32'ha7d7146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5160f, value : 32'h71a5a294},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51610, value : 32'hc7d6f1b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51611, value : 32'hc1bfc3ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51612, value : 32'h47084548},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51613, value : 32'h702cc08b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51614, value : 32'h8aeda50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51615, value : 32'h4668fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51616, value : 32'h10b10f29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51617, value : 32'h41c3750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51618, value : 32'h10362},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51619, value : 32'hffaf0ea2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5161a, value : 32'hc08b42c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5161b, value : 32'ha8a702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5161c, value : 32'h704c04a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5161d, value : 32'hd909700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5161e, value : 32'hffaf0ece},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5161f, value : 32'hc7cac28b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51620, value : 32'hc046700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51621, value : 32'hc044c045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51622, value : 32'h30041c28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51623, value : 32'h750cc049},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51624, value : 32'h41c3ef12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51625, value : 32'h10365},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51626, value : 32'hffaf0e6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51627, value : 32'h255442c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51628, value : 32'h25001f42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51629, value : 32'h1001f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5162a, value : 32'h25400020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5162b, value : 32'h4d5a1a03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5162c, value : 32'hf00f712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5162d, value : 32'h36341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5162e, value : 32'he4e0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5162f, value : 32'h42c1ffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51630, value : 32'h148c2540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51631, value : 32'h14022540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51632, value : 32'hd9094d48},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51633, value : 32'hc040dbc8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51634, value : 32'h940c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51635, value : 32'h70ad0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51636, value : 32'h37102440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51637, value : 32'h30112440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51638, value : 32'hc047c241},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51639, value : 32'h4083c442},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5163a, value : 32'hc343b030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5163b, value : 32'hc08bb031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5163c, value : 32'h80e702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5163d, value : 32'hda50fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5163e, value : 32'h24011104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5163f, value : 32'h1002c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51640, value : 32'h7825250e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51641, value : 32'hfdec18b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51642, value : 32'h42c10460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51643, value : 32'h41c140a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51644, value : 32'hffaf0e36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51645, value : 32'h71a5c28b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51646, value : 32'h91140dd7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51647, value : 32'h90110f63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51648, value : 32'hcf2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51649, value : 32'h78e0c7ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5164a, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5164b, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5164c, value : 32'h20143f05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5164d, value : 32'h22550042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5164e, value : 32'h922a0800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5164f, value : 32'h30401ce8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51650, value : 32'h1cec9228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51651, value : 32'h92263040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51652, value : 32'h30401cf0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51653, value : 32'h1cf49224},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51654, value : 32'h92223040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51655, value : 32'h30401cf8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51656, value : 32'h1cfc9220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51657, value : 32'h922c3040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51658, value : 32'h30581c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51659, value : 32'h1c41922e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5165a, value : 32'h92303058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5165b, value : 32'h30581c42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5165c, value : 32'h1c439232},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5165d, value : 32'h92343058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5165e, value : 32'h30581c44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5165f, value : 32'h1c459236},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51660, value : 32'h92383058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51661, value : 32'h30581c46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51662, value : 32'h1c47923a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51663, value : 32'h923c3058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51664, value : 32'h30581c48},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51665, value : 32'h1c49923e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51666, value : 32'h12403058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51667, value : 32'h1c4a0101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51668, value : 32'h12443058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51669, value : 32'h1c4b0101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5166a, value : 32'h12483058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5166b, value : 32'h1c4c0101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5166c, value : 32'h124c3058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5166d, value : 32'h1c4d0101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5166e, value : 32'h12503058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5166f, value : 32'h1c4e0101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51670, value : 32'h12543058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51671, value : 32'h1c4f0101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51672, value : 32'h12583058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51673, value : 32'h1c500101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51674, value : 32'h125c3058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51675, value : 32'h1c510101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51676, value : 32'h12603058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51677, value : 32'h1c520101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51678, value : 32'h12643058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51679, value : 32'h1c530101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5167a, value : 32'h12683058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5167b, value : 32'h1c540101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5167c, value : 32'h126c3058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5167d, value : 32'h1c550101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5167e, value : 32'h12703058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5167f, value : 32'h1c560101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51680, value : 32'h12743058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51681, value : 32'h1c570101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51682, value : 32'h12783058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51683, value : 32'h1c580101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51684, value : 32'h127c3058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51685, value : 32'h1c590101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51686, value : 32'h90203058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51687, value : 32'h30581c5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51688, value : 32'h1c5b9022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51689, value : 32'h90243058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5168a, value : 32'h30581c5c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5168b, value : 32'h1c5d9026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5168c, value : 32'h90283058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5168d, value : 32'h30581c5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5168e, value : 32'h1061014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5168f, value : 32'h1091018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51690, value : 32'h108101c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51691, value : 32'h10b1020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51692, value : 32'h90f490d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51693, value : 32'h909890b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51694, value : 32'h905c907a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51695, value : 32'h1040903e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51696, value : 32'h10440119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51697, value : 32'h10480118},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51698, value : 32'h104c0117},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51699, value : 32'h10500116},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5169a, value : 32'h10540115},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5169b, value : 32'h10580114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5169c, value : 32'h105c0113},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5169d, value : 32'h10600112},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5169e, value : 32'h10640111},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5169f, value : 32'h10680110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a0, value : 32'h106c011f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a1, value : 32'h1070011e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a2, value : 32'h10740105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a3, value : 32'h10780104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a4, value : 32'h107c0107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a5, value : 32'h2455011b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a6, value : 32'h18643800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a7, value : 32'h186006c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a8, value : 32'h185c01c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516a9, value : 32'h18580100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516aa, value : 32'h18540140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ab, value : 32'h18500780},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ac, value : 32'h184c07c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ad, value : 32'h18480400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ae, value : 32'h18440440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516af, value : 32'h18400480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b0, value : 32'h183c04c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b1, value : 32'h18380500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b2, value : 32'h18340540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b3, value : 32'h18300580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b4, value : 32'h182c05c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b5, value : 32'h18280600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b6, value : 32'ha0290640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b7, value : 32'ha441c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b8, value : 32'ha0480040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516b9, value : 32'ha086a067},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ba, value : 32'ha0e4a0a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516bb, value : 32'h1808a0c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516bc, value : 32'h180402c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516bd, value : 32'h18000200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516be, value : 32'h145e0240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516bf, value : 32'h1c7c3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c0, value : 32'h14fc3180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c1, value : 32'hc05e3002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c2, value : 32'h3600145d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c3, value : 32'h300314f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c4, value : 32'h300414f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c5, value : 32'h145cc05d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c6, value : 32'h14ec3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c7, value : 32'h14f03006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c8, value : 32'hc05c3005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516c9, value : 32'h3600145b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ca, value : 32'h300714e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516cb, value : 32'h145ac05b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516cc, value : 32'hc05a3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516cd, value : 32'h36001459},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ce, value : 32'h1458c059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516cf, value : 32'hc0583600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d0, value : 32'h36001457},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d1, value : 32'h1456c057},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d2, value : 32'hc0563600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d3, value : 32'h36001455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d4, value : 32'h1454c055},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d5, value : 32'hc0543600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d6, value : 32'h36001453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d7, value : 32'h1452c053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d8, value : 32'hc0523600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516d9, value : 32'h36001451},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516da, value : 32'h1450c051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516db, value : 32'hc0503600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516dc, value : 32'h3600144f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516dd, value : 32'h144ec04f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516de, value : 32'hc04e3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516df, value : 32'h3600144d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e0, value : 32'h144cc04d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e1, value : 32'hc04c3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e2, value : 32'h3600144b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e3, value : 32'h144ac04b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e4, value : 32'hc04a3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e5, value : 32'h36001449},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e6, value : 32'h1448c049},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e7, value : 32'hc0483600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e8, value : 32'h36001447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516e9, value : 32'h1446c047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ea, value : 32'hc0463600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516eb, value : 32'h36001445},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ec, value : 32'h1444c045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ed, value : 32'hc0443600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ee, value : 32'h36001443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ef, value : 32'h1442c043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f0, value : 32'hc0423600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f1, value : 32'h36001441},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f2, value : 32'h1440c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f3, value : 32'hc0403600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f4, value : 32'hffaf0b36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f5, value : 32'h2480740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f6, value : 32'h14043f05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f7, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f8, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516f9, value : 32'hc1bcb6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516fa, value : 32'h20557834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516fb, value : 32'h90580801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516fc, value : 32'h1051158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516fd, value : 32'h1071160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516fe, value : 32'h9054c259},
                          '{ step_type : REG_WRITE, reg_addr : 32'h516ff, value : 32'h1061168},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51700, value : 32'h1041018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51701, value : 32'h9050c25a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51702, value : 32'h1161010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51703, value : 32'h1171008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51704, value : 32'h1038c25b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51705, value : 32'h10400108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51706, value : 32'h10480119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51707, value : 32'h10500118},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51708, value : 32'h10580115},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51709, value : 32'h10600114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5170a, value : 32'h10680113},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5170b, value : 32'h10700112},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5170c, value : 32'h10780111},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5170d, value : 32'h1100011b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5170e, value : 32'h9164010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5170f, value : 32'h91ec9148},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51710, value : 32'h91b491d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51711, value : 32'h911c9198},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51712, value : 32'h1101140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51713, value : 32'h11f1148},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51714, value : 32'h11e1150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51715, value : 32'h1091170},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51716, value : 32'h1011178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51717, value : 32'h31801c58},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51718, value : 32'h31c01c54},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51719, value : 32'h31401c50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5171a, value : 32'h3005146c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5171b, value : 32'h30061468},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5171c, value : 32'h30071464},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5171d, value : 32'h41c3c158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5171e, value : 32'h1f00a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5171f, value : 32'h740cc050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51720, value : 32'h42e2c24b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51721, value : 32'h43c2c34a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51722, value : 32'h32401c5c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51723, value : 32'h37801c4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51724, value : 32'h37c01c48},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51725, value : 32'h34001c44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51726, value : 32'hc54ec44f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51727, value : 32'hc74cc64d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51728, value : 32'h32c01c24},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51729, value : 32'h36c01c20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5172a, value : 32'h34401c1c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5172b, value : 32'h34801c18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5172c, value : 32'h34c01c14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5172d, value : 32'h35001c10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5172e, value : 32'h35401c0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5172f, value : 32'h36001c08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51730, value : 32'h36401c04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51731, value : 32'hffaf0a42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51732, value : 32'h32001c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51733, value : 32'h1404c0bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51734, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51735, value : 32'hc1a2c2f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51736, value : 32'h70901600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51737, value : 32'h48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51738, value : 32'h20d02053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51739, value : 32'h710c702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5173a, value : 32'h70ae724e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5173b, value : 32'h1600e807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5173c, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5173d, value : 32'he8890025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5173e, value : 32'h1600f040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5173f, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51740, value : 32'h8810040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51741, value : 32'h251f0010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51742, value : 32'h2f8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51743, value : 32'h706e7000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51744, value : 32'h23002b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51745, value : 32'h60be70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51746, value : 32'hc809728e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51747, value : 32'h3812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51748, value : 32'h300255f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51749, value : 32'hf802030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5174a, value : 32'h5c08000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5174b, value : 32'hb8027825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5174c, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5174d, value : 32'h20539000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5174e, value : 32'h205300c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5174f, value : 32'h274c0107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51750, value : 32'h26ce8400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51751, value : 32'hb8250026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51752, value : 32'hc12053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51753, value : 32'h2340909},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51754, value : 32'h7813b8c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51755, value : 32'h41c3c141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51756, value : 32'h80069},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51757, value : 32'h750cc040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51758, value : 32'h43a24202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51759, value : 32'hffaf09a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5175a, value : 32'h4c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5175b, value : 32'h25ff248d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5175c, value : 32'h716671ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5175d, value : 32'ha1940b9d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5175e, value : 32'h228d700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5175f, value : 32'h71ae2ebe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51760, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51761, value : 32'h880012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51762, value : 32'h46e087d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51763, value : 32'h724e708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51764, value : 32'h2414710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51765, value : 32'h2800244e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51766, value : 32'hbe0c050f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51767, value : 32'h45cb706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51768, value : 32'h5d88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51769, value : 32'h7f0b8d04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5176a, value : 32'hc809f227},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5176b, value : 32'h3812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5176c, value : 32'h78258500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5176d, value : 32'hb89cb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5176e, value : 32'h9000b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5176f, value : 32'hc62053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51770, value : 32'h1072053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51771, value : 32'h8400274c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51772, value : 32'h2626ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51773, value : 32'h2053b825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51774, value : 32'h90b00c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51775, value : 32'hb8c20234},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51776, value : 32'hc1417813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51777, value : 32'h6a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51778, value : 32'hc0400008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51779, value : 32'h4202750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5177a, value : 32'h240a4322},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5177b, value : 32'h91a0500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5177c, value : 32'h250affaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5177d, value : 32'h716604c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5177e, value : 32'ha1b40bad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5177f, value : 32'h228de50c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51780, value : 32'h718e22bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51781, value : 32'h97d7126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51782, value : 32'hc0a2a114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51783, value : 32'h78e0c6d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51784, value : 32'hc1b7c3ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51785, value : 32'h41c3d840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51786, value : 32'h36a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51787, value : 32'h88a0b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51788, value : 32'h809110e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51789, value : 32'hffaf08e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5178a, value : 32'h2105750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5178b, value : 32'h700e2351},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5178c, value : 32'he58770ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5178d, value : 32'h260162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5178e, value : 32'h20c02178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5178f, value : 32'h10b50d0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51790, value : 32'h1209704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51791, value : 32'hf009360e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51792, value : 32'hd0f704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51793, value : 32'h70cd10b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51794, value : 32'h360e1209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51795, value : 32'hc083744e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51796, value : 32'haa6702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51797, value : 32'hda50fd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51798, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51799, value : 32'h8901122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5179a, value : 32'h8e38980},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5179b, value : 32'h742c0324},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5179c, value : 32'h29007882},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5179d, value : 32'h732c048f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5179e, value : 32'h49f2900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5179f, value : 32'h2900722c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a0, value : 32'h712c049e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a1, value : 32'h4852900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a2, value : 32'h40c36821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a3, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a4, value : 32'h841000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a5, value : 32'h7040240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a6, value : 32'h903843c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a7, value : 32'h20a80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a8, value : 32'hca905c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517a9, value : 32'h2c40032e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517aa, value : 32'h26f01347},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ab, value : 32'h8000734b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ac, value : 32'h27051100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ad, value : 32'hc2830387},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ae, value : 32'h11c02305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517af, value : 32'h3012215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b0, value : 32'h2300b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b1, value : 32'h78651146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b2, value : 32'h17892300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b3, value : 32'h23009000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b4, value : 32'hb10017c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b5, value : 32'h1c02605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b6, value : 32'h7865b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b7, value : 32'hb1089000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b8, value : 32'h11c02105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517b9, value : 32'h7865b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ba, value : 32'hb1109000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517bb, value : 32'h11c02005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517bc, value : 32'h7865b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517bd, value : 32'hb1189000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517be, value : 32'h7894710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517bf, value : 32'h12214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c0, value : 32'h2005b80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c1, value : 32'h23050382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c2, value : 32'h23001080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c3, value : 32'hb80213cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c4, value : 32'h90007865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c5, value : 32'h2605b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c6, value : 32'hb8020080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c7, value : 32'h90007865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c8, value : 32'h2105b108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517c9, value : 32'hb8021080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ca, value : 32'h90007865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517cb, value : 32'h2005b110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517cc, value : 32'hb8021080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517cd, value : 32'h2c22205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ce, value : 32'h90007865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517cf, value : 32'h6a12b118},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d0, value : 32'h90007865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d1, value : 32'h41940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d2, value : 32'h750c7185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d3, value : 32'h36b41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d4, value : 32'h42a10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d5, value : 32'hff6f0fb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d6, value : 32'h6e3470cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d7, value : 32'h6038c083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d8, value : 32'h1071008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517d9, value : 32'h1061006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517da, value : 32'h1041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517db, value : 32'h1051004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517dc, value : 32'h90459060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517dd, value : 32'h90079026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517de, value : 32'h42c1c240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517df, value : 32'h41c3c141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e0, value : 32'h9036c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e1, value : 32'hf82c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e2, value : 32'h750cff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e3, value : 32'hecf71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e4, value : 32'h71a59154},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e5, value : 32'h68c1f14f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e6, value : 32'h41c3750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e7, value : 32'h1036d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e8, value : 32'hff6f0f66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517e9, value : 32'h70ad4202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ea, value : 32'h209f4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517eb, value : 32'h20140401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ec, value : 32'h40c30341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ed, value : 32'hbf6c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ee, value : 32'h6113603a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ef, value : 32'h123c750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f0, value : 32'h41c30106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f1, value : 32'h5036e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f2, value : 32'h1051228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f3, value : 32'h1041214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f4, value : 32'hff6f0f36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f5, value : 32'h71a542a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f6, value : 32'h92540dd1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f7, value : 32'h20402040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f8, value : 32'h83a408b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517f9, value : 32'hc7cc710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517fa, value : 32'hb62c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517fb, value : 32'h702cfeef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517fc, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517fd, value : 32'h8ee0122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517fe, value : 32'h9418e21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h517ff, value : 32'h204003e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51800, value : 32'hc8090a8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51801, value : 32'h78a57aef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51802, value : 32'h2a406832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51803, value : 32'h78250380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51804, value : 32'h3ed41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51805, value : 32'hb8920004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51806, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51807, value : 32'h750c9060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51808, value : 32'h23534460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51809, value : 32'hee20145},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5180a, value : 32'h24adff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5180b, value : 32'h71e50982},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5180c, value : 32'h79ef8e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5180d, value : 32'h804508cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5180e, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5180f, value : 32'hc1b4c3e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51810, value : 32'h360d1209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51811, value : 32'h702cc080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51812, value : 32'hfd2f08b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51813, value : 32'h41c3da50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51814, value : 32'h369},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51815, value : 32'hff6f0eb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51816, value : 32'h2585750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51817, value : 32'hc1801203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51818, value : 32'h88240a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51819, value : 32'hda090460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5181a, value : 32'hd909700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5181b, value : 32'hff6f0eda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5181c, value : 32'hc7c2c280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5181d, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5181e, value : 32'ha023702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5181f, value : 32'ha021a022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51820, value : 32'ha0207fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51821, value : 32'h4200c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51822, value : 32'h780f7704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51823, value : 32'h4c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51824, value : 32'h207c0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51825, value : 32'hd5200c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51826, value : 32'h4050fd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51827, value : 32'h901c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51828, value : 32'h42c301c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51829, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5182a, value : 32'h20b00821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5182b, value : 32'hdc25706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5182c, value : 32'h831bc9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5182d, value : 32'h8c002071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5182e, value : 32'hb162b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5182f, value : 32'h9201b178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51830, value : 32'hd83fb200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51831, value : 32'hf00cb806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51832, value : 32'h1600b160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51833, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51834, value : 32'hb1020040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51835, value : 32'h9202b178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51836, value : 32'hd83fb200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51837, value : 32'hf011b110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51838, value : 32'h8c1bb100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51839, value : 32'hb178b102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5183a, value : 32'h20049110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5183b, value : 32'hf80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5183c, value : 32'hb110ffbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5183d, value : 32'haa008a02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5183e, value : 32'haa018a05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5183f, value : 32'hba2b170},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51840, value : 32'h400204e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51841, value : 32'h78e0c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51842, value : 32'h40c37014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51843, value : 32'h48a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51844, value : 32'h1600f207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51845, value : 32'h90387101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51846, value : 32'hb9800030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51847, value : 32'h9020f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51848, value : 32'h1e00b9a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51849, value : 32'h903b7044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5184a, value : 32'h7fe0c030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5184b, value : 32'h78e0b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5184c, value : 32'h4528c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5184d, value : 32'hfdaf096a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5184e, value : 32'hee154608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5184f, value : 32'h762cc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51850, value : 32'h746cda22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51851, value : 32'hb80244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51852, value : 32'h70cc45a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51853, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51854, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51855, value : 32'h1800c004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51856, value : 32'h98a0045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51857, value : 32'h700cfdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51858, value : 32'h700cf013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51859, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5185a, value : 32'h244a706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5185b, value : 32'h45a10b80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5185c, value : 32'hfdef0972},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5185d, value : 32'hc80970cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5185e, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5185f, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51860, value : 32'h1800c004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51861, value : 32'h700c0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51862, value : 32'hfdef090a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51863, value : 32'hc6c4712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51864, value : 32'h4628c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51865, value : 32'h21534508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51866, value : 32'h710c0142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51867, value : 32'hfd2f0b02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51868, value : 32'hbe23702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51869, value : 32'h16022644},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5186a, value : 32'h8540655d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5186b, value : 32'h85017a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5186c, value : 32'ha5407826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5186d, value : 32'hc6c4a501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5186e, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5186f, value : 32'h18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51870, value : 32'h7ce0b8e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51871, value : 32'h900f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51872, value : 32'h704cc068},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51873, value : 32'h4c02150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51874, value : 32'hb040b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51875, value : 32'h900840c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51876, value : 32'hb0400068},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51877, value : 32'h804519d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51878, value : 32'h804518a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51879, value : 32'h18007fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5187a, value : 32'h78e000c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5187b, value : 32'h3c32841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5187c, value : 32'h3c12840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5187d, value : 32'h28417b25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5187e, value : 32'h21440341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5187f, value : 32'h28410081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51880, value : 32'h7b2500c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51881, value : 32'h2c12841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51882, value : 32'h1012144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51883, value : 32'h12284},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51884, value : 32'h28417b25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51885, value : 32'h21440241},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51886, value : 32'h7b250201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51887, value : 32'h1c12841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51888, value : 32'h4012144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51889, value : 32'h28417b25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5188a, value : 32'h21440141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5188b, value : 32'h79650801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5188c, value : 32'h79456875},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5188d, value : 32'h22847a1d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5188e, value : 32'h23840002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5188f, value : 32'h79450010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51890, value : 32'h22847a1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51891, value : 32'h79450004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51892, value : 32'h22846853},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51893, value : 32'h79450008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51894, value : 32'h7b25704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51895, value : 32'hba8b6837},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51896, value : 32'h23057944},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51897, value : 32'h2840004c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51898, value : 32'h795b0243},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51899, value : 32'h28407964},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5189a, value : 32'h7c2502c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5189b, value : 32'h79646a32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5189c, value : 32'h10432405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5189d, value : 32'h3412840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5189e, value : 32'h78246a13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5189f, value : 32'h7fe07b05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a0, value : 32'h78e07870},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a1, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a2, value : 32'hc1a9b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a3, value : 32'h800041db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a4, value : 32'h43101228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a5, value : 32'h308f1100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a6, value : 32'h4338b8c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a7, value : 32'h207841e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a8, value : 32'h219f0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518a9, value : 32'h40100582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518aa, value : 32'h2c1209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ab, value : 32'h800141d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ac, value : 32'h60384e7c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ad, value : 32'hef047022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ae, value : 32'hf003d94d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518af, value : 32'h880cd932},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b0, value : 32'h42c3b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b1, value : 32'h504901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b2, value : 32'h8920710f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b3, value : 32'h2014c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b4, value : 32'hc80923ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b5, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b6, value : 32'h214411e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b7, value : 32'h704e0054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b8, value : 32'h2fc7268a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518b9, value : 32'h900447d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ba, value : 32'hb8020224},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518bb, value : 32'h832005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518bc, value : 32'h6041b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518bd, value : 32'h86041aa4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518be, value : 32'hf822005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518bf, value : 32'hc0909007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c0, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c1, value : 32'h909004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c2, value : 32'hb8889000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c3, value : 32'h66a8b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c4, value : 32'h20250a3d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c5, value : 32'h20166f14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c6, value : 32'h70420400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c7, value : 32'h60a8e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c8, value : 32'h3952840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518c9, value : 32'h25c02505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ca, value : 32'h5841800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518cb, value : 32'h2e00c3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518cc, value : 32'h2740740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518cd, value : 32'h71462201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ce, value : 32'h20402505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518cf, value : 32'h5841800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d0, value : 32'h20056904},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d1, value : 32'h18000540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d2, value : 32'hf1e30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d3, value : 32'h20802b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d4, value : 32'h20057077},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d5, value : 32'hf2ca04d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d6, value : 32'hd9104022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d7, value : 32'h4a00f66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d8, value : 32'h20132452},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518d9, value : 32'hd9104022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518da, value : 32'h2600e9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518db, value : 32'h4022da41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518dc, value : 32'hfaad910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518dd, value : 32'hdaf3fdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518de, value : 32'hf4a4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518df, value : 32'hd90b04a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e0, value : 32'hd90b4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e1, value : 32'hfdef0f96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e2, value : 32'h4022daf0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e3, value : 32'h4a00f36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e4, value : 32'h4022d912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e5, value : 32'he72d912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e6, value : 32'hda080260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e7, value : 32'hd9124022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e8, value : 32'hfdef0f7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518e9, value : 32'h9dedaf8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ea, value : 32'h208afdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518eb, value : 32'hd1a0c12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ec, value : 32'h700c0160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ed, value : 32'hfd4f0ed2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ee, value : 32'h40c36829},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ef, value : 32'h4888000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f0, value : 32'h4e00dda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f1, value : 32'h40c3b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f2, value : 32'h13880000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f3, value : 32'h2e00bc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f4, value : 32'he02d90c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f5, value : 32'h402204c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f6, value : 32'he2ed90d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f7, value : 32'hda400260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f8, value : 32'h4e00d56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518f9, value : 32'hc081c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518fa, value : 32'hffef0daa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518fb, value : 32'hc081d90d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518fc, value : 32'hffef0da2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518fd, value : 32'hc081732c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518fe, value : 32'hffef0d9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h518ff, value : 32'hc081d90b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51900, value : 32'hffef0d92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51901, value : 32'hc081d911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51902, value : 32'hffef0d8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51903, value : 32'h1600d912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51904, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51905, value : 32'h80f0131},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51906, value : 32'hc0810071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51907, value : 32'hffef0d76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51908, value : 32'hb89d913},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51909, value : 32'h40222421},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5190a, value : 32'h4a00e9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5190b, value : 32'h4022d911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5190c, value : 32'hdd6d911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5190d, value : 32'hda080260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5190e, value : 32'hd9114022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5190f, value : 32'hfdef0ede},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51910, value : 32'h4022daef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51911, value : 32'hdc2d911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51912, value : 32'hda200260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51913, value : 32'h4e00cea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51914, value : 32'hc085c085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51915, value : 32'hffef0d3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51916, value : 32'h4102d911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51917, value : 32'h30801100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51918, value : 32'h2c1219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51919, value : 32'h209f704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5191a, value : 32'hc3850582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5191b, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5191c, value : 32'h710c6119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5191d, value : 32'h4002800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5191e, value : 32'hb8027122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5191f, value : 32'h400200f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51920, value : 32'h6a009f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51921, value : 32'h208a780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51922, value : 32'hb0a041f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51923, value : 32'h702c02e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51924, value : 32'hfbe4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51925, value : 32'hd9110420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51926, value : 32'hcaac081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51927, value : 32'hd90b04e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51928, value : 32'hca2c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51929, value : 32'hd91104e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5192a, value : 32'h40e14102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5192b, value : 32'h2c1219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5192c, value : 32'h209f704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5192d, value : 32'hc3810582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5192e, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5192f, value : 32'h202f6119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51930, value : 32'h9b20487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51931, value : 32'h712206a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51932, value : 32'hd9104022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51933, value : 32'hfdef0e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51934, value : 32'h4022daf3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51935, value : 32'hd32d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51936, value : 32'hda610260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51937, value : 32'hd9104022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51938, value : 32'hfdef0e3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51939, value : 32'hf011da7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5193a, value : 32'hd9104022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5193b, value : 32'hfdef0e2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5193c, value : 32'h4022daf3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5193d, value : 32'hd12d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5193e, value : 32'hda610260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5193f, value : 32'hd9104022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51940, value : 32'h2600d06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51941, value : 32'h4002da80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51942, value : 32'h70451e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51943, value : 32'h4c4901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51944, value : 32'h24210c21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51945, value : 32'h2c1209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51946, value : 32'hda1041e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51947, value : 32'h582219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51948, value : 32'h6119716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51949, value : 32'h487202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5194a, value : 32'h6a00b16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5194b, value : 32'hf0447122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5194c, value : 32'h35012800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5194d, value : 32'h210fb902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5194e, value : 32'h11000514},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5194f, value : 32'h219f3081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51950, value : 32'h60380582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51951, value : 32'hd5a7022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51952, value : 32'h1010fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51953, value : 32'h9ae0093},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51954, value : 32'hc3e0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51955, value : 32'h222f04c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51956, value : 32'hd8100487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51957, value : 32'hfdef095a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51958, value : 32'h700c4162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51959, value : 32'h872742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5195a, value : 32'h714cfdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5195b, value : 32'h22822384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5195c, value : 32'h507222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5195d, value : 32'h21412385},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5195e, value : 32'h93ed810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5195f, value : 32'h4162fdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51960, value : 32'hd920700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51961, value : 32'hfdef0852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51962, value : 32'h700c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51963, value : 32'hfdaf0d06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51964, value : 32'hd0e712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51965, value : 32'hb32fd4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51966, value : 32'h700c0160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51967, value : 32'h4c00bce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51968, value : 32'hcf2700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51969, value : 32'h702cfdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5196a, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5196b, value : 32'h9e61388},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5196c, value : 32'hd91402e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5196d, value : 32'he81866a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5196e, value : 32'h6f14706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5196f, value : 32'h4002016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51970, value : 32'he0247062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51971, value : 32'hd88060a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51972, value : 32'h4e00d5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51973, value : 32'h2a404230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51974, value : 32'h71662392},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51975, value : 32'h2f812205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51976, value : 32'h2309004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51977, value : 32'h66a8b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51978, value : 32'ha0040bdb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51979, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5197a, value : 32'h9aa1388},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5197b, value : 32'hd90c02e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5197c, value : 32'h4008a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5197d, value : 32'h4c00bde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5197e, value : 32'h340c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5197f, value : 32'h996d090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51980, value : 32'h702c02e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51981, value : 32'h30151400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51982, value : 32'h4e00b92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51983, value : 32'h21d5254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51984, value : 32'he81866a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51985, value : 32'h6f14706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51986, value : 32'h4002016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51987, value : 32'he0247062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51988, value : 32'h40a260a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51989, value : 32'h4e00cfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5198a, value : 32'h2a404230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5198b, value : 32'h71662392},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5198c, value : 32'h2f812205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5198d, value : 32'h2309004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5198e, value : 32'h66a8b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5198f, value : 32'ha0040bdb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51990, value : 32'h40c3d90c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51991, value : 32'h13880000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51992, value : 32'h2e0094a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51993, value : 32'h66a84410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51994, value : 32'h254fe819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51995, value : 32'h706e2215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51996, value : 32'h20166f14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51997, value : 32'h70620400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51998, value : 32'h60a9e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51999, value : 32'hcbe40a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5199a, value : 32'h423004e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5199b, value : 32'h23922a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5199c, value : 32'h22057166},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5199d, value : 32'h90042f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5199e, value : 32'hb1000230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5199f, value : 32'hbdd66a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a0, value : 32'h4082a004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a1, value : 32'h2e0090e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a2, value : 32'h66a8d90c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a3, value : 32'h704ee825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a4, value : 32'h20166f14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a5, value : 32'h70420400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a6, value : 32'h60a9e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a7, value : 32'h6208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a8, value : 32'h4e00c82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519a9, value : 32'h2b404330},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519aa, value : 32'h24052394},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ab, value : 32'h90042f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ac, value : 32'hb1000224},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ad, value : 32'h2e008b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ae, value : 32'h208a740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519af, value : 32'hc660006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b0, value : 32'h416204e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b1, value : 32'h2f812405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b2, value : 32'h22c9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b3, value : 32'h7146b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b4, value : 32'hac166a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b5, value : 32'h40c3a004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b6, value : 32'hd0900003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b7, value : 32'h2e008b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b8, value : 32'h4022702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519b9, value : 32'h4200d6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ba, value : 32'haead910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519bb, value : 32'hc0a904c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519bc, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519bd, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519be, value : 32'h40d3c2f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519bf, value : 32'h1e8901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c0, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c1, value : 32'h10000fff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c2, value : 32'h10102112},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c3, value : 32'h18102111},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c4, value : 32'h18002005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c5, value : 32'hc8092004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c6, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c7, value : 32'h900c0f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c8, value : 32'h90400020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519c9, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ca, value : 32'h88001226},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519cb, value : 32'h201204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519cc, value : 32'h1e006058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519cd, value : 32'h901c7044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ce, value : 32'h20420508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519cf, value : 32'h160000d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d0, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d1, value : 32'h70140114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d2, value : 32'hd93df281},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d3, value : 32'hb910750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d4, value : 32'hff2f0fb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d5, value : 32'h47cb70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d6, value : 32'h1188000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d7, value : 32'h45cb8f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d8, value : 32'h1003e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519d9, value : 32'hfa2750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519da, value : 32'h41a1ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519db, value : 32'h10562740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519dc, value : 32'h1401254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519dd, value : 32'h20821600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519de, value : 32'hff2f0f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519df, value : 32'h2640750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e0, value : 32'h71ad2057},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e1, value : 32'h20821700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e2, value : 32'h750cbd96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e3, value : 32'hff2f0f7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e4, value : 32'h274241a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e5, value : 32'h254f10d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e6, value : 32'h14001401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e7, value : 32'hf6a2082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e8, value : 32'h750cff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519e9, value : 32'h20532440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ea, value : 32'h1441254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519eb, value : 32'h20821300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ec, value : 32'hf56750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ed, value : 32'h4038ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ee, value : 32'h204f6fa9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ef, value : 32'h8d403401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f0, value : 32'hff2f0f46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f1, value : 32'h710c750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f2, value : 32'he808722d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f3, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f4, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f5, value : 32'hf037e887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f6, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f7, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f8, value : 32'hc809e835},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519f9, value : 32'h13812e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519fa, value : 32'h7180244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519fb, value : 32'h8b2840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519fc, value : 32'ha4020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519fd, value : 32'h3de208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519fe, value : 32'h201143e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h519ff, value : 32'h40a18380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a00, value : 32'h4062f40f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a01, value : 32'h11300e1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a02, value : 32'he1343c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a03, value : 32'h40621330},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a04, value : 32'h12f00e0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a05, value : 32'he2743c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a06, value : 32'h40821151},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a07, value : 32'h210543e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a08, value : 32'h884002c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a09, value : 32'h20058b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a0a, value : 32'h90001f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a0b, value : 32'hb40001c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a0c, value : 32'h1f802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a0d, value : 32'h1b49000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a0e, value : 32'h71c5b040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a0f, value : 32'h71c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a10, value : 32'hde074000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a11, value : 32'h10ff218d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a12, value : 32'h45cb700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a13, value : 32'h11408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a14, value : 32'h108015e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a15, value : 32'h27c12d42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a16, value : 32'h7824b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a17, value : 32'h1e0070a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a18, value : 32'h901c7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a19, value : 32'h40c30510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a1a, value : 32'h2af80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a1b, value : 32'h2a00f26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a1c, value : 32'h1800702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a1d, value : 32'h18102484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a1e, value : 32'h15e62444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a1f, value : 32'h781d1080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a20, value : 32'h7704b8a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a21, value : 32'hc6d8ad01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a22, value : 32'he36c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a23, value : 32'h40100600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a24, value : 32'h700c71ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a25, value : 32'h900f45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a26, value : 32'hd940c298},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a27, value : 32'h73c41e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a28, value : 32'hc028900f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a29, value : 32'h2a00eee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a2a, value : 32'h1e00b5e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a2b, value : 32'h902f73c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a2c, value : 32'he3ecc40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a2d, value : 32'h700c0360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a2e, value : 32'h2a00e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a2f, value : 32'h1d00d810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a30, value : 32'h16001005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a31, value : 32'h9018710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a32, value : 32'h8150018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a33, value : 32'h26842030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a34, value : 32'h1e001c07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a35, value : 32'h901b73c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a36, value : 32'hf02ec000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a37, value : 32'h901b45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a38, value : 32'h264fc018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a39, value : 32'h702c1280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a3a, value : 32'heaab500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a3b, value : 32'h208a02a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a3c, value : 32'h702c0a0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a3d, value : 32'hf40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a3e, value : 32'he9a4240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a3f, value : 32'h1dec02a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a40, value : 32'h160093c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a41, value : 32'h90187101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a42, value : 32'h1de8004c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a43, value : 32'hb9c493c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a44, value : 32'h90051dec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a45, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a46, value : 32'h48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a47, value : 32'h8002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a48, value : 32'h78c5b804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a49, value : 32'hc809b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a4a, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a4b, value : 32'h90180f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a4c, value : 32'hb0200024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a4d, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a4e, value : 32'h89001228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a4f, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a50, value : 32'h111bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a51, value : 32'h88216038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a52, value : 32'hdf090d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a53, value : 32'h21538834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a54, value : 32'hf20480fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a55, value : 32'h4c0098a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a56, value : 32'h70451e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a57, value : 32'hc0b49027},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a58, value : 32'h78e0c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a59, value : 32'hc1a3c3f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a5a, value : 32'h2140250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a5b, value : 32'h3100200a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a5c, value : 32'h47504670},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a5d, value : 32'h71344430},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a5e, value : 32'h2d012e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a5f, value : 32'hc8094210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a60, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a61, value : 32'hb802122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a62, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a63, value : 32'h1909038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a64, value : 32'h8159000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a65, value : 32'h1600025e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a66, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a67, value : 32'h701400f3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a68, value : 32'h10246},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a69, value : 32'h208a70d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a6a, value : 32'h218a003e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a6b, value : 32'hf2e2001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a6c, value : 32'h21cafd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a6d, value : 32'h8fa02002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a6e, value : 32'h132079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a6f, value : 32'h22132340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a70, value : 32'h75308f21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a71, value : 32'hd019e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a72, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a73, value : 32'h880012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a74, value : 32'h36e08c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a75, value : 32'hd137aaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a76, value : 32'h40622030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a77, value : 32'hca64182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a78, value : 32'h43420060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a79, value : 32'ha86f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a7a, value : 32'h40400020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a7b, value : 32'h234e2614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a7c, value : 32'h20700a25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a7d, value : 32'ha4fb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a7e, value : 32'h212f2031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a7f, value : 32'hf2138348},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a80, value : 32'h500997},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a81, value : 32'h90099b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a82, value : 32'hd1093b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a83, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a84, value : 32'hf01c014a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a85, value : 32'h8348222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a86, value : 32'h41c3f209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a87, value : 32'h14c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a88, value : 32'h41c3f008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a89, value : 32'h1478000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a8a, value : 32'h41c3f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a8b, value : 32'h14b8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a8c, value : 32'h83227c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a8d, value : 32'h21ca7074},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a8e, value : 32'h80000f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a8f, value : 32'ha0d014d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a90, value : 32'h41c300d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a91, value : 32'h14e8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a92, value : 32'h901100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a93, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a94, value : 32'hd8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a95, value : 32'h17e092f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a96, value : 32'he12c182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a97, value : 32'h94a0040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a98, value : 32'h140904a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a99, value : 32'hc2223080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a9a, value : 32'h8740813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a9b, value : 32'h16812500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a9c, value : 32'h1e0a0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a9d, value : 32'h43191c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a9e, value : 32'hafdf005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51a9f, value : 32'h191c801e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa0, value : 32'h96200003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa1, value : 32'h24402000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa2, value : 32'h2108780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa3, value : 32'h49100001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa4, value : 32'h71a5b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa5, value : 32'h41c3f196},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa6, value : 32'h1488000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa7, value : 32'h41c3f1d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa8, value : 32'h1498000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aa9, value : 32'h2450f1d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aaa, value : 32'h8bf2000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aab, value : 32'h708d00b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aac, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aad, value : 32'hdc3122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aae, value : 32'h73962030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aaf, value : 32'h20c82478},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab0, value : 32'h126124ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab1, value : 32'h12482040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab2, value : 32'hfd2f0e12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab3, value : 32'h12892c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab4, value : 32'h108615b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab5, value : 32'h15014700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab6, value : 32'h8d60108b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab7, value : 32'h1887371},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab8, value : 32'he7f000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ab9, value : 32'h2b4000ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aba, value : 32'hc8090301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51abb, value : 32'h47cb7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51abc, value : 32'hffff0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51abd, value : 32'h4812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51abe, value : 32'h69b270cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51abf, value : 32'h42814021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac0, value : 32'h2050a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac1, value : 32'h310f11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac2, value : 32'h6812300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac3, value : 32'h811120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac4, value : 32'h400a2b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac5, value : 32'h20b10c13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac6, value : 32'h3412005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac7, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac8, value : 32'h1e89004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ac9, value : 32'h2505f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aca, value : 32'h90041f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51acb, value : 32'h912000a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51acc, value : 32'h210871f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51acd, value : 32'h27ca038e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ace, value : 32'h20801045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51acf, value : 32'h71440010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad0, value : 32'h66fef1e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad1, value : 32'h20c22614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad2, value : 32'h268c79dd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad3, value : 32'h21809002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad4, value : 32'h21ca003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad5, value : 32'hb2200025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad6, value : 32'h20c22714},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad7, value : 32'h7164b220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad8, value : 32'h8fa0f1be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ad9, value : 32'h700cf07e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ada, value : 32'h39f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51adb, value : 32'ha7a0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51adc, value : 32'h4282fcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51add, value : 32'h4042f078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ade, value : 32'h714cc180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51adf, value : 32'hc441716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae0, value : 32'ha009d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae1, value : 32'h4042c440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae2, value : 32'h714cc180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae3, value : 32'ha009c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae4, value : 32'h8d01706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae5, value : 32'h8d18d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae6, value : 32'h784200a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae7, value : 32'h2a922240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae8, value : 32'hc8096821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ae9, value : 32'h7040240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aea, value : 32'h78020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aeb, value : 32'h3012a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aec, value : 32'h79057142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aed, value : 32'hb992b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aee, value : 32'hb99fb99c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aef, value : 32'hc1809180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af0, value : 32'h8321f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af1, value : 32'h6479bcc5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af2, value : 32'h8032142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af3, value : 32'h7930e120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af4, value : 32'h2614e1c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af5, value : 32'h23ca2081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af6, value : 32'hb1600025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af7, value : 32'h20812714},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af8, value : 32'hb1607144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51af9, value : 32'h8f21f040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51afa, value : 32'h9798fa0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51afb, value : 32'h49b00364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51afc, value : 32'h40c36841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51afd, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51afe, value : 32'h240a8880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51aff, value : 32'h40a17080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b00, value : 32'h20a8dac1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b01, value : 32'hc0d0240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b02, value : 32'h2614102e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b03, value : 32'hb3402003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b04, value : 32'hf0287104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b05, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b06, value : 32'h880012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b07, value : 32'h34e0843},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b08, value : 32'h234026f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b09, value : 32'h600c46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b0a, value : 32'hca05c182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b0b, value : 32'hc082e805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b0c, value : 32'h2200b5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b0d, value : 32'h16004103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b0e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b0f, value : 32'h815000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b10, value : 32'h2500017e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b11, value : 32'h101c1680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b12, value : 32'hb460081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b13, value : 32'hc0820220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b14, value : 32'hb6ac082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b15, value : 32'h2714ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b16, value : 32'h8f21234e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b17, value : 32'h71a5b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b18, value : 32'h834509b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b19, value : 32'h78e0c7d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b1a, value : 32'h2840c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b1b, value : 32'h4200038c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b1c, value : 32'h1f812405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b1d, value : 32'hab09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b1e, value : 32'h70ec9100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b1f, value : 32'h3204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b20, value : 32'hb8a0b160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b21, value : 32'h2a40b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b22, value : 32'hc8090301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b23, value : 32'h69127905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b24, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b25, value : 32'hab49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b26, value : 32'hb1d9060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b27, value : 32'h46600175},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b28, value : 32'h208040c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b29, value : 32'h7825080a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b2a, value : 32'hb892b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b2b, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b2c, value : 32'h1071000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b2d, value : 32'h1f802405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b2e, value : 32'h3549004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b2f, value : 32'h16009000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b30, value : 32'h80007101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b31, value : 32'h90d0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b32, value : 32'hf84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b33, value : 32'h781d0a6b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b34, value : 32'h211f7910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b35, value : 32'h20020180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b36, value : 32'hb80601c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b37, value : 32'h402805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b38, value : 32'h804218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b39, value : 32'h8252f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b3a, value : 32'h7d104910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b3b, value : 32'h1442053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b3c, value : 32'h11832d41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b3d, value : 32'h39941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b3e, value : 32'ha0e0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b3f, value : 32'h740cff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b40, value : 32'hc6c240a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b41, value : 32'h1822053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b42, value : 32'h1c120ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b43, value : 32'h7fe0a941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b44, value : 32'h78e0a900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b45, value : 32'hc1a4c3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b46, value : 32'h40c34410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b47, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b48, value : 32'h202f8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b49, value : 32'h20440502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b4a, value : 32'h43300052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b4b, value : 32'hd84de903},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b4c, value : 32'hd832f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b4d, value : 32'h8800b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b4e, value : 32'ha0db8c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b4f, value : 32'h712c2020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b50, value : 32'h4800cb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b51, value : 32'hffcf09b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b52, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b53, value : 32'ha46c350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b54, value : 32'h732c02a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b55, value : 32'h40c3d90b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b56, value : 32'h4e7c8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b57, value : 32'h3e00ef2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b58, value : 32'h40224110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b59, value : 32'h3e00eea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b5a, value : 32'h4022d911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b5b, value : 32'h3e00ee2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b5c, value : 32'h46cbd912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b5d, value : 32'h11e28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b5e, value : 32'h4a00c22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b5f, value : 32'h24cf2214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b60, value : 32'he81a67c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b61, value : 32'h21152b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b62, value : 32'h251670ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b63, value : 32'h60b82480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b64, value : 32'h60c9e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b65, value : 32'h4208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b66, value : 32'h4a00d8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b67, value : 32'h28404030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b68, value : 32'h71a52390},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b69, value : 32'h2f812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b6a, value : 32'h2309004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b6b, value : 32'h67c8b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b6c, value : 32'h90040ddb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b6d, value : 32'h40c3d90c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b6e, value : 32'h13880000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b6f, value : 32'h2a009d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b70, value : 32'hc124010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b71, value : 32'hc8090480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b72, value : 32'h70ad702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b73, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b74, value : 32'h901c0f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b75, value : 32'h18000504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b76, value : 32'h9ba0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b77, value : 32'h400202a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b78, value : 32'hce24022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b79, value : 32'hd9100460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b7a, value : 32'hd9104022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b7b, value : 32'hfdaf0d2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b7c, value : 32'h4022dacf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b7d, value : 32'hd26d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b7e, value : 32'hdafffdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b7f, value : 32'h4a00b3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b80, value : 32'hc080c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b81, value : 32'hffaf0b8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b82, value : 32'h4142d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b83, value : 32'h219f4062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b84, value : 32'h704c02c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b85, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b86, value : 32'h718cc380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b87, value : 32'h611970ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b88, value : 32'h8524082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b89, value : 32'h71220660},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b8a, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b8b, value : 32'h96636b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b8c, value : 32'hd90a02a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b8d, value : 32'he81567c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b8e, value : 32'h21002b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b8f, value : 32'h4802016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b90, value : 32'h71a560b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b91, value : 32'h60c8e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b92, value : 32'h2005b80e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b93, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b94, value : 32'h700c0230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b95, value : 32'hb100b88c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b96, value : 32'hde167c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b97, value : 32'h40229004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b98, value : 32'h3e00dee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b99, value : 32'hc809d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b9a, value : 32'h21056832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b9b, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b9c, value : 32'h2105c090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b9d, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b9e, value : 32'h91200090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51b9f, value : 32'hf812104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba0, value : 32'hfeff0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba1, value : 32'h882b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba2, value : 32'hd81402a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba3, value : 32'h78e0c7d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba4, value : 32'h46cbc2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba5, value : 32'h1e8901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba6, value : 32'h96a89620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba7, value : 32'h25464030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba8, value : 32'hb6081c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ba9, value : 32'hf802105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51baa, value : 32'hc300000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bab, value : 32'h1600b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bac, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bad, value : 32'he8360114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bae, value : 32'h750cd945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51baf, value : 32'hff2f084a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb0, value : 32'hc809b910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb1, value : 32'h726d702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb2, value : 32'h710c68f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb3, value : 32'h1600e807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb4, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb5, value : 32'he8880025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb6, value : 32'h1600f020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb7, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb8, value : 32'he8200040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bb9, value : 32'h7180244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bba, value : 32'h60020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bbb, value : 32'h3802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bbc, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bbd, value : 32'h78e519b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bbe, value : 32'h4c22f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bbf, value : 32'hf832005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc0, value : 32'h1c09000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc1, value : 32'he21cb380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc2, value : 32'hf832005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc3, value : 32'h1b49000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc4, value : 32'h4022f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc5, value : 32'hb3007124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc6, value : 32'h238dd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc7, value : 32'h700c16bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc8, value : 32'h901c40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bc9, value : 32'h18000508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bca, value : 32'h18080005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bcb, value : 32'h40c30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bcc, value : 32'h2af80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bcd, value : 32'h2a0085e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bce, value : 32'h1e00702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bcf, value : 32'hb6a81404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd0, value : 32'h78e0c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd1, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd2, value : 32'hc1a7b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd3, value : 32'hd9114528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd4, value : 32'h4608b913},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd5, value : 32'hc344d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd6, value : 32'hfeef0fae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd7, value : 32'hd8c8c243},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd8, value : 32'hd945ed04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bd9, value : 32'hf004b911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bda, value : 32'hb910d989},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bdb, value : 32'hfecf0f9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bdc, value : 32'hc18640a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bdd, value : 32'h35c22440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bde, value : 32'ha00afa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bdf, value : 32'h35832440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be0, value : 32'hee05d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be1, value : 32'hb912d923},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be2, value : 32'hd98bf003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be3, value : 32'hf7ab910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be4, value : 32'hc006fecf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be5, value : 32'h8d41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be6, value : 32'hc0410001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be7, value : 32'hf6ad8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be8, value : 32'hc201feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51be9, value : 32'h30801417},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bea, value : 32'h8e45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51beb, value : 32'h41a10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bec, value : 32'hd8c8c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bed, value : 32'hfeef0f52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bee, value : 32'h1416c200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bef, value : 32'h254f3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf0, value : 32'hc0421401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf1, value : 32'hf42d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf2, value : 32'hc202feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf3, value : 32'h46cbc203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf4, value : 32'h10090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf5, value : 32'hf32d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf6, value : 32'h41c1feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf7, value : 32'h264fdd20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf8, value : 32'hbd9f1401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bf9, value : 32'hf22d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bfa, value : 32'h1501feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bfb, value : 32'h8d401482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bfc, value : 32'h144f264f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bfd, value : 32'hf12d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bfe, value : 32'h41e1feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51bff, value : 32'h908215f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c00, value : 32'h1401274f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c01, value : 32'hfeef0f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c02, value : 32'h15f7d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c03, value : 32'h264f9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c04, value : 32'hd8c8148f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c05, value : 32'hfeef0ef2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c06, value : 32'h8d4441e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c07, value : 32'h1401274f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c08, value : 32'hfeef0ee6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c09, value : 32'h8d5fd8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c0a, value : 32'hd8c8bf91},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c0b, value : 32'hfeef0eda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c0c, value : 32'h274f41e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c0d, value : 32'hd8c81401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c0e, value : 32'hfeef0ece},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c0f, value : 32'h264fda0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c10, value : 32'hd8c814c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c11, value : 32'hfeef0ec2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c12, value : 32'hd999744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c13, value : 32'hebad8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c14, value : 32'hb910feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c15, value : 32'h7014c001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c16, value : 32'h2c013e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c17, value : 32'hc000704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c18, value : 32'h47d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c19, value : 32'h201f0a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c1a, value : 32'h2f4005c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c1b, value : 32'hc00420c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c1c, value : 32'h800046d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c1d, value : 32'h201f1a44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c1e, value : 32'h26400059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c1f, value : 32'h72232090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c20, value : 32'h5952200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c21, value : 32'h20902000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c22, value : 32'hc002c100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c23, value : 32'h6408f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c24, value : 32'h2540230a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c25, value : 32'h240ac600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c26, value : 32'hc0032400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c27, value : 32'h4a00a86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c28, value : 32'h431879cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c29, value : 32'hbc1702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c2a, value : 32'hd8c8346e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c2b, value : 32'h4342c204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c2c, value : 32'h9a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c2d, value : 32'h44c10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c2e, value : 32'hfeef0e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c2f, value : 32'h440250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c30, value : 32'hd8c8d99b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c31, value : 32'hfeef0e42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c32, value : 32'h70adb910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c33, value : 32'h34c0200a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c34, value : 32'h1704478a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c35, value : 32'hd8c81503},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c36, value : 32'h35021004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c37, value : 32'h9c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c38, value : 32'he260003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c39, value : 32'h44a1feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c3a, value : 32'he5c071a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c3b, value : 32'hd99df7b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c3c, value : 32'he16d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c3d, value : 32'hb910feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c3e, value : 32'hd8c8dd4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c3f, value : 32'he0abd11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c40, value : 32'h41a1feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c41, value : 32'h1401254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c42, value : 32'hfeef0dfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c43, value : 32'h221ad8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c44, value : 32'h2f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c45, value : 32'h261a28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c46, value : 32'h452a15c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c47, value : 32'h1184259a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c48, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c49, value : 32'h71231b46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c4a, value : 32'hda66038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c4b, value : 32'h651d05e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c4c, value : 32'h260065eb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c4d, value : 32'h65fd2341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c4e, value : 32'h7021180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c4f, value : 32'h11041502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c50, value : 32'hbb22e807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c51, value : 32'h41c3d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c52, value : 32'h300a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c53, value : 32'hd8c8f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c54, value : 32'ha141c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c55, value : 32'hdb20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c56, value : 32'hd951fecf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c57, value : 32'hdaad8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c58, value : 32'hb911feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c59, value : 32'h23807126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c5a, value : 32'h93f2184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c5b, value : 32'h2480a2b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c5c, value : 32'hc0022184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c5d, value : 32'h7267610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c5e, value : 32'h71c5ffe5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c5f, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c60, value : 32'h250028f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c61, value : 32'h20002015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c62, value : 32'h71462010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c63, value : 32'h220cc001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c64, value : 32'h6f8a000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c65, value : 32'hd9a3ffcb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c66, value : 32'hd6ed8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c67, value : 32'hb910feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c68, value : 32'h1404c0a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c69, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c6a, value : 32'hc1a2c3f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c6b, value : 32'h40c34310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c6c, value : 32'h122d8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c6d, value : 32'h800041d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c6e, value : 32'h88000025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c6f, value : 32'h11004748},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c70, value : 32'h4628208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c71, value : 32'h30021c03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c72, value : 32'hc181710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c73, value : 32'h30c22440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c74, value : 32'ha008a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c75, value : 32'h30c32440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c76, value : 32'h30121404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c77, value : 32'h10c02478},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c78, value : 32'h20087104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c79, value : 32'h84f0490},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c7a, value : 32'h44102072},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c7b, value : 32'hb1170ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c7c, value : 32'h740c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c7d, value : 32'ha941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c7e, value : 32'hf0050003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c7f, value : 32'ha841c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c80, value : 32'h42a10003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c81, value : 32'hd0243a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c82, value : 32'h44c1feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c83, value : 32'h15250d11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c84, value : 32'h41c1700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c85, value : 32'hd5e42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c86, value : 32'h43a1ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c87, value : 32'h14a30d11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c88, value : 32'h41c1710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c89, value : 32'hd4e42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c8a, value : 32'h43a1ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c8b, value : 32'hdc371a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c8c, value : 32'h11e59404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c8d, value : 32'h81fa080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c8e, value : 32'h4062003e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c8f, value : 32'h42c1702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c90, value : 32'hffef0d06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c91, value : 32'h406243e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c92, value : 32'h42c1712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c93, value : 32'hffef0cfa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c94, value : 32'hc7d043e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c95, value : 32'h2482c3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c96, value : 32'h42203608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c97, value : 32'h740c4210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c98, value : 32'h21841c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c99, value : 32'hca20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c9a, value : 32'h4450feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c9b, value : 32'hc1804042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c9c, value : 32'hfe2f0fda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c9d, value : 32'h35c22440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c9e, value : 32'h3108b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51c9f, value : 32'hc0864708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca0, value : 32'h200902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca1, value : 32'hc0204142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca2, value : 32'hc2864182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca3, value : 32'he0a4342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca4, value : 32'h4110fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca5, value : 32'h70cd4510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca6, value : 32'h70ed454a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca7, value : 32'h200a706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca8, value : 32'he7c02440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ca9, value : 32'h9500f755},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51caa, value : 32'h505081f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cab, value : 32'hc1b9501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cac, value : 32'h78cf2025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cad, value : 32'hc2864182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cae, value : 32'hfe2f0dde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51caf, value : 32'hb0b4342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb0, value : 32'h43102005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb1, value : 32'he60840d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb2, value : 32'he708e520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb3, value : 32'h74edf1eb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb4, value : 32'h2000740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb5, value : 32'h4508200e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb6, value : 32'he0bf78cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb7, value : 32'h4182f70a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb8, value : 32'hdb6c286},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cb9, value : 32'h4342fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cba, value : 32'h20050b09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cbb, value : 32'h40d14310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cbc, value : 32'h234e2002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cbd, value : 32'he0bf78cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cbe, value : 32'h4182f70a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cbf, value : 32'hd9ac286},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc0, value : 32'h4342fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc1, value : 32'h20050b09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc2, value : 32'h40d14310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc3, value : 32'h91350dc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc4, value : 32'hb1d78bd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc5, value : 32'h230c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc6, value : 32'h1a82a540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc7, value : 32'h21ca251c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc8, value : 32'h22802402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cc9, value : 32'h70ed2084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cca, value : 32'h24421a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ccb, value : 32'hc7d240e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ccc, value : 32'h4708c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ccd, value : 32'hb8226901},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cce, value : 32'h20494528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ccf, value : 32'h740c0fce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd0, value : 32'h41c342a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd1, value : 32'h20219},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd2, value : 32'hfeef0bbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd3, value : 32'h271543c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd4, value : 32'h90601380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd5, value : 32'ha179041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd6, value : 32'h740c00e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd7, value : 32'h21a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd8, value : 32'hba60002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cd9, value : 32'h74adfeef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cda, value : 32'h40e1f00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cdb, value : 32'h2080627a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cdc, value : 32'ha8a00084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cdd, value : 32'h70ad785d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cde, value : 32'h101c1f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cdf, value : 32'hc6c640a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce0, value : 32'h2155c0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce1, value : 32'h248a0f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce2, value : 32'h708d7001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce3, value : 32'h238a704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce4, value : 32'h20a80fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce5, value : 32'h20160280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce6, value : 32'h7144008f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce7, value : 32'hb762b783},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce8, value : 32'hb760b781},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ce9, value : 32'h2115716d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cea, value : 32'h234002cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ceb, value : 32'h94401048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cec, value : 32'hd3794a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ced, value : 32'h211510a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cee, value : 32'h93a00203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cef, value : 32'ha119341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf0, value : 32'h20160364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf1, value : 32'hb2a002c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf2, value : 32'hb2619361},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf3, value : 32'h910214fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf4, value : 32'h910314fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf5, value : 32'ha40b65},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf6, value : 32'h2c32016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf7, value : 32'h14feb340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf8, value : 32'hb3419102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cf9, value : 32'h2016f02a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cfa, value : 32'h774402cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cfb, value : 32'h9340b541},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cfc, value : 32'h232f7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cfd, value : 32'h14fc1088},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cfe, value : 32'h71449102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51cff, value : 32'h22097a50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d00, value : 32'hb54002c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d01, value : 32'h1086232f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d02, value : 32'h23099c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d03, value : 32'h77441082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d04, value : 32'h9441b540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d05, value : 32'hb5427144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d06, value : 32'h77449341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d07, value : 32'h14fe7b50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d08, value : 32'h77449102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d09, value : 32'h22087a50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d0a, value : 32'hb54300c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d0b, value : 32'h9c417b4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d0c, value : 32'h822308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d0d, value : 32'hb5437144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d0e, value : 32'h9ff4086f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d0f, value : 32'h1200230a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d10, value : 32'h91619140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d11, value : 32'ha50b17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d12, value : 32'h91427744},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d13, value : 32'hb3b9163},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d14, value : 32'hb0400084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d15, value : 32'hb0419143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d16, value : 32'hb041f017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d17, value : 32'h71449142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d18, value : 32'h7b4eb040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d19, value : 32'h23099940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d1a, value : 32'h77440082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d1b, value : 32'h9141b040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d1c, value : 32'hb0427144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d1d, value : 32'h77449143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d1e, value : 32'h7b4eb043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d1f, value : 32'h23089941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d20, value : 32'h71440082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d21, value : 32'h9642b043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d22, value : 32'h10311fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d23, value : 32'ha50b1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d24, value : 32'h96407744},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d25, value : 32'h10311fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d26, value : 32'h840b41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d27, value : 32'h11fab740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d28, value : 32'hb7210101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d29, value : 32'hb741f01a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d2a, value : 32'h71449640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d2b, value : 32'h7b4eb740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d2c, value : 32'h23099e42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d2d, value : 32'h77440082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d2e, value : 32'h11feb740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d2f, value : 32'h71440102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d30, value : 32'h11fab742},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d31, value : 32'h77440102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d32, value : 32'h7a4eb743},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d33, value : 32'h14111fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d34, value : 32'h412208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d35, value : 32'hb7237124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d36, value : 32'h7f80244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d37, value : 32'h34020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d38, value : 32'h9159024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d39, value : 32'hf81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d3a, value : 32'h218affff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d3b, value : 32'h180a0fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d3c, value : 32'hb0240005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d3d, value : 32'hc4c6e008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d3e, value : 32'h1600c2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d3f, value : 32'h8000708f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d40, value : 32'h46cb122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d41, value : 32'h1a468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d42, value : 32'h40584770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d43, value : 32'h46104138},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d44, value : 32'h10912642},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d45, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d46, value : 32'h122b8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d47, value : 32'h1627710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d48, value : 32'h40c3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d49, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d4a, value : 32'h20118800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d4b, value : 32'hf2a783c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d4c, value : 32'h81370ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d4d, value : 32'h27003031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d4e, value : 32'h10201680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d4f, value : 32'h75100080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d50, value : 32'hd0bf299},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d51, value : 32'h70f61271},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d52, value : 32'h248af295},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d53, value : 32'h70ec7001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d54, value : 32'h706d700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d55, value : 32'h70cc702d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d56, value : 32'h20a8706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d57, value : 32'h40c30d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d58, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d59, value : 32'h261f791b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d5a, value : 32'h211f2002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d5b, value : 32'hb8223041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d5c, value : 32'h615978ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d5d, value : 32'h40a1611a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d5e, value : 32'h184209a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d5f, value : 32'h20156058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d60, value : 32'h213401c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d61, value : 32'h60d0200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d62, value : 32'h3250829},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d63, value : 32'heb174050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d64, value : 32'h2c7222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d65, value : 32'h207212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d66, value : 32'h222f4953},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d67, value : 32'h212f0187},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d68, value : 32'h79420247},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d69, value : 32'h23ca7170},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d6a, value : 32'h20ca1189},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d6b, value : 32'hf0071249},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d6c, value : 32'h26ca7074},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d6d, value : 32'h210a01c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d6e, value : 32'h203d11c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d6f, value : 32'h71e40303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d70, value : 32'h2c7212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d71, value : 32'h207202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d72, value : 32'h212f4832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d73, value : 32'h202f0187},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d74, value : 32'h78220247},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d75, value : 32'h23ca7050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d76, value : 32'h20ca118a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d77, value : 32'h222f124a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d78, value : 32'h232f22c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d79, value : 32'h23002207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d7a, value : 32'h242f2480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d7b, value : 32'h16002002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d7c, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d7d, value : 32'he82600ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d7e, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d7f, value : 32'h158000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d80, value : 32'h9f0841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d81, value : 32'h5c008ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d82, value : 32'h40a1e80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d83, value : 32'h184209a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d84, value : 32'h20157002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d85, value : 32'h21340500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d86, value : 32'h60d02001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d87, value : 32'hf0047822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d88, value : 32'h24802302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d89, value : 32'h3086120b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d8a, value : 32'h6252f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d8b, value : 32'h180253f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d8c, value : 32'h23741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d8d, value : 32'h42c20005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d8e, value : 32'hfae43e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d8f, value : 32'h44a1fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d90, value : 32'h209a40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d91, value : 32'h20000184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d92, value : 32'h26562010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d93, value : 32'h70021800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d94, value : 32'h5e0087e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d95, value : 32'h5021800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d96, value : 32'h2015e80d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d97, value : 32'h60d12500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d98, value : 32'h20002134},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d99, value : 32'h791d6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d9a, value : 32'h2f802000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d9b, value : 32'h1b488000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d9c, value : 32'h71a5b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d9d, value : 32'h6bee58a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d9e, value : 32'h71e5ffc5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51d9f, value : 32'hc6daf14c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da0, value : 32'h7034c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da1, value : 32'h3012a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da2, value : 32'h79654608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da3, value : 32'h47cbc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da4, value : 32'h409004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da5, value : 32'h27c07825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da6, value : 32'h28401222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da7, value : 32'he688008b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da8, value : 32'h404846c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51da9, value : 32'h26126ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51daa, value : 32'h45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dab, value : 32'h702dffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dac, value : 32'h706c708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dad, value : 32'h1a50b37},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dae, value : 32'he137890},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51daf, value : 32'h20001275},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db0, value : 32'h10201680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db1, value : 32'hb1f0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db2, value : 32'h21050000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db3, value : 32'h78e512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db4, value : 32'hfeef0902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db5, value : 32'h79b09000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db6, value : 32'h4d2009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db7, value : 32'h20087990},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db8, value : 32'h2180004c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51db9, value : 32'h71641010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dba, value : 32'h79b0f1e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dbb, value : 32'h781d6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dbc, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dbd, value : 32'h44cbc0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dbe, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dbf, value : 32'h108814b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc0, value : 32'h14008ce1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc1, value : 32'hf9b1086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc2, value : 32'h8931184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc3, value : 32'h244a11ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc4, value : 32'h265a7280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc5, value : 32'h20a8028b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc6, value : 32'h446900c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc7, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc8, value : 32'h249ac14c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dc9, value : 32'h2432100e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dca, value : 32'h80001f89},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dcb, value : 32'h927c44c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dcc, value : 32'h659e10f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dcd, value : 32'h10b00915},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dce, value : 32'h7135659e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dcf, value : 32'h702d70ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd0, value : 32'h2434f417},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd1, value : 32'hf0131347},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd2, value : 32'h13472434},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd3, value : 32'h11091602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd4, value : 32'h2434f00f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd5, value : 32'h16021347},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd6, value : 32'hdd801109},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd7, value : 32'h21029682},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd8, value : 32'h7d8211c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dd9, value : 32'h3450c0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dda, value : 32'h218a4781},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ddb, value : 32'h21001002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ddc, value : 32'h211411cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ddd, value : 32'h7e9d02cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dde, value : 32'h18c20f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ddf, value : 32'hb58064dc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de0, value : 32'h2cd2214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de1, value : 32'h18c20f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de2, value : 32'hb58074e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de3, value : 32'h2cd2314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de4, value : 32'h18c20f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de5, value : 32'h74217165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de6, value : 32'h71c4b580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de7, value : 32'hc4c6f1b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de8, value : 32'h706cc0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51de9, value : 32'h2240dc3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dea, value : 32'h248a008b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51deb, value : 32'h18007001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dec, value : 32'ha9800003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ded, value : 32'h1c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dee, value : 32'h15081304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51def, value : 32'h10110809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df0, value : 32'hf0037164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df1, value : 32'h2280a860},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df2, value : 32'h248a0f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df3, value : 32'h20a87001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df4, value : 32'h12fc01c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df5, value : 32'heb858503},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df6, value : 32'h89807785},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df7, value : 32'ha980f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df8, value : 32'h7b8f8840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51df9, value : 32'hca0b4b51},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dfa, value : 32'h44207110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dfb, value : 32'hf649700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dfc, value : 32'h21e41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dfd, value : 32'hf120003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dfe, value : 32'hd8c9feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51dff, value : 32'hc0d1760c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e00, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e01, value : 32'h7002248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e02, value : 32'h20a8706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e03, value : 32'h41000480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e04, value : 32'h182235a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e05, value : 32'he219a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e06, value : 32'h41c3623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e07, value : 32'hc14c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e08, value : 32'h61596234},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e09, value : 32'h90d9121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e0a, value : 32'h71640305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e0b, value : 32'hd8807fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e0c, value : 32'h786f7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e0d, value : 32'hf717e1ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e0e, value : 32'h7a22da80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e0f, value : 32'h7080240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e10, value : 32'h44020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e11, value : 32'h215a4200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e12, value : 32'h229a0183},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e13, value : 32'h635b000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e14, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e15, value : 32'h6354c14c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e16, value : 32'h9241627a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e17, value : 32'h3040a09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e18, value : 32'hd9807124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e19, value : 32'h78307fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e1a, value : 32'h1422053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e1b, value : 32'ha941b826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e1c, value : 32'ha9007fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e1d, value : 32'hc1a3c3ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e1e, value : 32'h700c4210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e1f, value : 32'h458b4130},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e20, value : 32'hb504b505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e21, value : 32'h18f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e22, value : 32'hb5030000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e23, value : 32'he7ab502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e24, value : 32'h740cfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e25, value : 32'h4122710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e26, value : 32'h32822440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e27, value : 32'h200eee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e28, value : 32'h31832440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e29, value : 32'h4122700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e2a, value : 32'hee2c282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e2b, value : 32'hc3810020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e2c, value : 32'h3140140a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e2d, value : 32'h2042d980},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e2e, value : 32'h40c38443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e2f, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e30, value : 32'h23ca9582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e31, value : 32'h8840002c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e32, value : 32'he411e4ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e33, value : 32'h24ca95e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e34, value : 32'h1406104d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e35, value : 32'h7e703110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e36, value : 32'h740c7d90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e37, value : 32'h19041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e38, value : 32'h43420007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e39, value : 32'h45c1718c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e3a, value : 32'h400260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e3b, value : 32'he1a47e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e3c, value : 32'hc540feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e3d, value : 32'h13840d1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e3e, value : 32'h23e40817},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e3f, value : 32'h27cc7512},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e40, value : 32'hf7599385},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e41, value : 32'h41224042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e42, value : 32'h43e1704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e43, value : 32'h4042f00d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e44, value : 32'h704c4122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e45, value : 32'h44a143e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e46, value : 32'hfcaf0dd2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e47, value : 32'h404270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e48, value : 32'h704c4122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e49, value : 32'h240a43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e4a, value : 32'hdc20400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e4b, value : 32'h71acfcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e4c, value : 32'he15c7cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e4d, value : 32'hdeb13c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e4e, value : 32'h40429424},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e4f, value : 32'h704c4122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e50, value : 32'hf00f43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e51, value : 32'h14250d13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e52, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e53, value : 32'h191},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e54, value : 32'hfe8f0db6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e55, value : 32'h4042c7cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e56, value : 32'h704c4122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e57, value : 32'h44a143e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e58, value : 32'h78e0f1e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e59, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e5a, value : 32'h24aa0458},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e5b, value : 32'h21aa1144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e5c, value : 32'h82610104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e5d, value : 32'h200e8200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e5e, value : 32'ha2008040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e5f, value : 32'h90c12403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e60, value : 32'ha2217fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e61, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e62, value : 32'hc1b6b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e63, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e64, value : 32'h8ea0122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e65, value : 32'h780f4310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e66, value : 32'h714cc180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e67, value : 32'h1c04706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e68, value : 32'h24403001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e69, value : 32'hbae3019},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e6a, value : 32'h1c000020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e6b, value : 32'h23403001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e6c, value : 32'h23402a18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e6d, value : 32'hd962a9b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e6e, value : 32'h255f0360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e6f, value : 32'h16001251},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e70, value : 32'h272f1092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e71, value : 32'h8e011487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e72, value : 32'h3e40885},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e73, value : 32'h2f412354},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e74, value : 32'h33cd21f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e75, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e76, value : 32'h103e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e77, value : 32'hfeaf0d2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e78, value : 32'h2f4042a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e79, value : 32'hc8091315},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e7a, value : 32'h26c12505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e7b, value : 32'h900447cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e7c, value : 32'h78250000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e7d, value : 32'hb802708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e7e, value : 32'h2440270a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e7f, value : 32'h902078e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e80, value : 32'h1502153},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e81, value : 32'he5207502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e82, value : 32'h2348262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e83, value : 32'h5c7222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e84, value : 32'h7854c082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e85, value : 32'h3e741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e86, value : 32'h43020004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e87, value : 32'hb0a04440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e88, value : 32'hce6740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e89, value : 32'h250afeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e8a, value : 32'h71860580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e8b, value : 32'h507202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e8c, value : 32'h827408dd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e8d, value : 32'h250571e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e8e, value : 32'hc8092601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e8f, value : 32'h21007825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e90, value : 32'hb8022511},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e91, value : 32'h78e57146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e92, value : 32'hf1bdb0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e93, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e94, value : 32'h714cc182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e95, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e96, value : 32'h6200976},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e97, value : 32'hc0b670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e98, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e99, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e9a, value : 32'hd820c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e9b, value : 32'h900745cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e9c, value : 32'h1d00c40c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e9d, value : 32'hc921045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e9e, value : 32'h1d000220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51e9f, value : 32'hd8201005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea0, value : 32'h2200c86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea1, value : 32'h10451d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea2, value : 32'h10051d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea3, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea4, value : 32'h803c2042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea5, value : 32'h42c3f208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea6, value : 32'h12f28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea7, value : 32'h10020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea8, value : 32'h521a14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ea9, value : 32'h620006d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eaa, value : 32'h78e0712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eab, value : 32'h2496c3ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eac, value : 32'h70ed3bef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ead, value : 32'h42e14508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eae, value : 32'h38802455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eaf, value : 32'he42ba8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb0, value : 32'h702cfc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb1, value : 32'h78b8710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb2, value : 32'hdeab802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb3, value : 32'h200f0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb4, value : 32'hdee0350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb5, value : 32'h20400020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb6, value : 32'h208c0791},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb7, value : 32'hdefe8e82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb8, value : 32'hddef705},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eb9, value : 32'h20540000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eba, value : 32'h740c088e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ebb, value : 32'h40441c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ebc, value : 32'h714c0002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ebd, value : 32'hfeaf0c12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ebe, value : 32'h120943a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ebf, value : 32'hc084360d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec0, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec1, value : 32'hde2104a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec2, value : 32'hda78fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec3, value : 32'hfbec084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec4, value : 32'hd97805e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec5, value : 32'h1e00d80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec6, value : 32'h900773c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec7, value : 32'h8cac29c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec8, value : 32'hd90ffdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ec9, value : 32'h212f78cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eca, value : 32'hd960447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ecb, value : 32'h222f0160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ecc, value : 32'h46cb0407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ecd, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ece, value : 32'h25058e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ecf, value : 32'h11f8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed0, value : 32'h8e20002a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed1, value : 32'h640827},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed2, value : 32'hb90e7822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed3, value : 32'h6d527104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed4, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed5, value : 32'h2c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed6, value : 32'h402205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed7, value : 32'h71c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed8, value : 32'hb89c4000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ed9, value : 32'h1800b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eda, value : 32'h70ed0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51edb, value : 32'h87ad80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51edc, value : 32'hd90ffdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51edd, value : 32'hf1e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ede, value : 32'h712cfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51edf, value : 32'h8e208e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee0, value : 32'h64084d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee1, value : 32'h6f417822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee2, value : 32'h240a7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee3, value : 32'h20a87000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee4, value : 32'h29400800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee5, value : 32'h245502c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee6, value : 32'h60783880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee7, value : 32'h30c2940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee8, value : 32'h26f460fb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ee9, value : 32'h80007040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eea, value : 32'h7885048c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eeb, value : 32'hb8027124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eec, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eed, value : 32'h2dc9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eee, value : 32'h20799000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eef, value : 32'hab000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef0, value : 32'h13402405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef1, value : 32'hb89cb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef2, value : 32'hb040b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef3, value : 32'h3400b7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef4, value : 32'hf9d71e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef5, value : 32'h9f84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef6, value : 32'h8ea00800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef7, value : 32'h38912455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef8, value : 32'h2d40700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ef9, value : 32'h210012c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51efa, value : 32'h8e012011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51efb, value : 32'h36408bd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51efc, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51efd, value : 32'h10405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51efe, value : 32'hfeaf0b0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51eff, value : 32'h70ed42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f00, value : 32'h9fdf278c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f01, value : 32'h2d0098},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f02, value : 32'h278bd981},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f03, value : 32'h1c0c9803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f04, value : 32'h1c083400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f05, value : 32'hf4123400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f06, value : 32'h18002756},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f07, value : 32'h11822f41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f08, value : 32'hf802004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f09, value : 32'hffc00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f0a, value : 32'h41c3b826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f0b, value : 32'h20406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f0c, value : 32'had66869},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f0d, value : 32'h740cfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f0e, value : 32'h702cda08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f0f, value : 32'h700cc382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f10, value : 32'h244a633b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f11, value : 32'h736d7100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f12, value : 32'h1440200a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f13, value : 32'h31b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f14, value : 32'h20020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f15, value : 32'h148c1001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f16, value : 32'h12cc2c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f17, value : 32'h78857765},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f18, value : 32'h71247426},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f19, value : 32'hb3f228d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f1a, value : 32'h140dab00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f1b, value : 32'h140b3087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f1c, value : 32'h140c3085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f1d, value : 32'h140a3086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f1e, value : 32'hc2223084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f1f, value : 32'h30831409},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f20, value : 32'h3081140e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f21, value : 32'h3080140f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f22, value : 32'h41c3c140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f23, value : 32'h80407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f24, value : 32'ha76c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f25, value : 32'h740cfeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f26, value : 32'hf1b4e720},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f27, value : 32'ha6a740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f28, value : 32'hb913feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f29, value : 32'hf1a371a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f2a, value : 32'h78e0c7ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f2b, value : 32'h82e43e3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f2c, value : 32'h20780000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f2d, value : 32'h16000001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f2e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f2f, value : 32'h8110008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f30, value : 32'h217800b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f31, value : 32'hb8020000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f32, value : 32'h7b007404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f33, value : 32'h2178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f34, value : 32'h7204781b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f35, value : 32'h78e07b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f36, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f37, value : 32'h88201228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f38, value : 32'h219f8841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f39, value : 32'h229f0582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f3a, value : 32'h10bc02c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f3b, value : 32'h60380000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f3c, value : 32'h8a03621a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f3d, value : 32'h86002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f3e, value : 32'h2002078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f3f, value : 32'h20ca7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f40, value : 32'h78e000a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f41, value : 32'h244ac5e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f42, value : 32'h706c71c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f43, value : 32'h702c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f44, value : 32'h900c44cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f45, value : 32'h20a80240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f46, value : 32'h21050280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f47, value : 32'h7424030d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f48, value : 32'h651d95a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f49, value : 32'h7144ad40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f4a, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f4b, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f4c, value : 32'h244ae90e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f4d, value : 32'h704c71c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f4e, value : 32'h28020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f4f, value : 32'h1381244f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f50, value : 32'h74447945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f51, value : 32'h61199120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f52, value : 32'h7164a967},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f53, value : 32'h78e0c4c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f54, value : 32'h4310c2f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f55, value : 32'h4570710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f56, value : 32'h42304450},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f57, value : 32'hfcaf0d42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f58, value : 32'h4cd2800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f59, value : 32'h10512553},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f5a, value : 32'hd90b700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f5b, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f5c, value : 32'h250a708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f5d, value : 32'hd6e0440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f5e, value : 32'h70ccfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f5f, value : 32'hd9ff700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f60, value : 32'hfd2f0856},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f61, value : 32'h6d12704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f62, value : 32'h200f762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f63, value : 32'hda2204c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f64, value : 32'h700c7e0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f65, value : 32'h20300d1d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f66, value : 32'h244adb40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f67, value : 32'h45c10a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f68, value : 32'hfcef0d42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f69, value : 32'hd88070cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f6a, value : 32'h744cd919},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f6b, value : 32'hf00cdb83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f6c, value : 32'h940244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f6d, value : 32'hd2e45c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f6e, value : 32'h70ccfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f6f, value : 32'hd919d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f70, value : 32'hdb81744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f71, value : 32'h250a708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f72, value : 32'hd1a0440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f73, value : 32'h70ccfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f74, value : 32'hcc2700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f75, value : 32'h712cfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f76, value : 32'h92e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f77, value : 32'hb88b0220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f78, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f79, value : 32'h9ae9c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f7a, value : 32'hd9080220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f7b, value : 32'h20300d0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f7c, value : 32'hd92640c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f7d, value : 32'hd923f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f7e, value : 32'hfe8f0f6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f7f, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f80, value : 32'h8fa0122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f81, value : 32'h82b8f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f82, value : 32'h79af0344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f83, value : 32'hb3e4062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f84, value : 32'h403000a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f85, value : 32'h4002e809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f86, value : 32'hb92742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f87, value : 32'h42620360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f88, value : 32'h23412214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f89, value : 32'h8f01b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f8a, value : 32'h71a57510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f8b, value : 32'hd0df7af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f8c, value : 32'h40c12030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f8d, value : 32'hf003d927},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f8e, value : 32'hf2ed924},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f8f, value : 32'h8fa0fe8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f90, value : 32'hb7d8f61},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f91, value : 32'h7eaf0364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f92, value : 32'hb024062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f93, value : 32'h41c100a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f94, value : 32'h40c1e834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f95, value : 32'hb56742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f96, value : 32'h42620360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f97, value : 32'h22f4b808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f98, value : 32'h22142341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f99, value : 32'h78252342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f9a, value : 32'h1600b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f9b, value : 32'h80007101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f9c, value : 32'h218c0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f9d, value : 32'hf70581c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f9e, value : 32'h451a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51f9f, value : 32'h7810f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa0, value : 32'h95080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa1, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa2, value : 32'hf009ffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa3, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa4, value : 32'h88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa5, value : 32'h2905b911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa6, value : 32'hb2000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa7, value : 32'hd117b10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa8, value : 32'h740c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fa9, value : 32'h35641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51faa, value : 32'hf0050002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fab, value : 32'h35741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fac, value : 32'h8560002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fad, value : 32'h42a1feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fae, value : 32'hf1c471a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51faf, value : 32'hb298fa0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb0, value : 32'h79af0364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb1, value : 32'ha00a86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb2, value : 32'he88b4062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb3, value : 32'h103f0d0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb4, value : 32'h23402214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb5, value : 32'hf0049021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb6, value : 32'h810110fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb7, value : 32'h8f61b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb8, value : 32'hf1ef71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fb9, value : 32'hb438f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fba, value : 32'hc3f0084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fbb, value : 32'h23782030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fbc, value : 32'hd0f2000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fbd, value : 32'h20782030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fbe, value : 32'h48ac0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fbf, value : 32'h489cf002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc0, value : 32'h68614b50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc1, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc2, value : 32'h70c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc3, value : 32'h20a86892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc4, value : 32'h2a400340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc5, value : 32'h22f40380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc6, value : 32'h78852081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc7, value : 32'hb8927144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc8, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fc9, value : 32'hb7ab020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fca, value : 32'h700cfc8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fcb, value : 32'h744cd90c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fcc, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fcd, value : 32'h440250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fce, value : 32'hfcef0baa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fcf, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd0, value : 32'h764cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd1, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd2, value : 32'hb9a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd3, value : 32'h268afcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd4, value : 32'h700c0fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd5, value : 32'h744cd910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd6, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd7, value : 32'h440250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd8, value : 32'hfcef0b82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fd9, value : 32'hd88070cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fda, value : 32'h764cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fdb, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fdc, value : 32'hb7270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fdd, value : 32'h268afcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fde, value : 32'h700c0fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fdf, value : 32'hfcef0b16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe0, value : 32'hc26712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe1, value : 32'hc6d20380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe2, value : 32'hc1a4c3ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe3, value : 32'h45484668},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe4, value : 32'h41104030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe5, value : 32'hf7970ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe6, value : 32'h244a11f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe7, value : 32'h40c37200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe8, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fe9, value : 32'h20300925},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fea, value : 32'h706c8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51feb, value : 32'h34020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fec, value : 32'h209f4020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fed, value : 32'h2000001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fee, value : 32'h2f402002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fef, value : 32'h60581200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff0, value : 32'he8156068},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff1, value : 32'hf022e312},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff2, value : 32'h20a8db7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff3, value : 32'h40200400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff4, value : 32'h1c209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff5, value : 32'h20022000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff6, value : 32'h12002f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff7, value : 32'h60786058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff8, value : 32'h801080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ff9, value : 32'hbb72e808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ffa, value : 32'hc080f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ffb, value : 32'h18541c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ffc, value : 32'hf0060002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ffd, value : 32'h41c3c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51ffe, value : 32'h20186},
                          '{ step_type : REG_WRITE, reg_addr : 32'h51fff, value : 32'hb06078f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52000, value : 32'hf06740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52001, value : 32'h42e1fe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52002, value : 32'hf1c771e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52003, value : 32'h31001400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52004, value : 32'h71c0244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52005, value : 32'hb500c280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52006, value : 32'h20a8b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52007, value : 32'h120203c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52008, value : 32'h95600501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52009, value : 32'hc50909},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5200a, value : 32'h9600b520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5200b, value : 32'h450809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5200c, value : 32'hb6204020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5200d, value : 32'hc7ca78e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5200e, value : 32'he808702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5200f, value : 32'h8002222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52010, value : 32'h6119b8c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52011, value : 32'hf5fc4040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52012, value : 32'h78307fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52013, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52014, value : 32'h2909008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52015, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52016, value : 32'h9b6c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52017, value : 32'ha0afd8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52018, value : 32'h4508fdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52019, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5201a, value : 32'h1c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5201b, value : 32'he80ce906},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5201c, value : 32'hd87ded8b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5201d, value : 32'hf019b807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5201e, value : 32'hed8ce80b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5201f, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52020, value : 32'hf0134650},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52021, value : 32'h40c3ed0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52022, value : 32'h4a380000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52023, value : 32'hed0af00d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52024, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52025, value : 32'hf0095208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52026, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52027, value : 32'hf0052ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52028, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52029, value : 32'hefe36b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5202a, value : 32'h742c01e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5202b, value : 32'hc6c2780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5202c, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5202d, value : 32'h7ed12e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5202e, value : 32'h8000fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5202f, value : 32'h45cbc2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52030, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52031, value : 32'h8d218d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52032, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52033, value : 32'h2c1219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52034, value : 32'h100215bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52035, value : 32'h60386058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52036, value : 32'hb8248801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52037, value : 32'hfcaf09b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52038, value : 32'h58e205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52039, value : 32'h832079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5203a, value : 32'h8d418d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5203b, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5203c, value : 32'h2c1229f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5203d, value : 32'h100115bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5203e, value : 32'h285239f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5203f, value : 32'h60586038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52040, value : 32'h63db8803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52041, value : 32'hd80ab8e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52042, value : 32'h22120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52043, value : 32'h2332631b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52044, value : 32'h80000f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52045, value : 32'hc6c407e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52046, value : 32'h4568c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52047, value : 32'h4050db7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52048, value : 32'h44604220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52049, value : 32'h248ae983},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5204a, value : 32'h8d850fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5204b, value : 32'h11041d06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5204c, value : 32'hea14e80e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5204d, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5204e, value : 32'h1468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5204f, value : 32'h40c3e91e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52050, value : 32'h1408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52051, value : 32'hb5268861},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52052, value : 32'hf0158820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52053, value : 32'h1d08710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52054, value : 32'hb8901001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52055, value : 32'hc6c8a503},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52056, value : 32'h20100831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52057, value : 32'h71011600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52058, value : 32'h1428000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52059, value : 32'h40c3e92e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5205a, value : 32'h1388000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5205b, value : 32'hb5269062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5205c, value : 32'hb5249020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5205d, value : 32'hf031b565},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5205e, value : 32'h11041d0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5205f, value : 32'h10051d08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52060, value : 32'h1d0cec2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52061, value : 32'hf0291085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52062, value : 32'h71011600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52063, value : 32'h1448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52064, value : 32'h40c3e918},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52065, value : 32'h13e8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52066, value : 32'h10fc9060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52067, value : 32'hb5268100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52068, value : 32'hb504b565},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52069, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5206a, value : 32'hb8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5206b, value : 32'h17e082b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5206c, value : 32'h8008238c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5206d, value : 32'h10051d08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5206e, value : 32'h238af78f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5206f, value : 32'hf1dc0fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52070, value : 32'hfc7238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52071, value : 32'h11041d0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52072, value : 32'h10051d08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52073, value : 32'h1d0cec04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52074, value : 32'hf0031205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52075, value : 32'h41c3b506},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52076, value : 32'h30227},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52077, value : 32'hfc2f0c0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52078, value : 32'hc0243d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52079, value : 32'h1104150c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5207a, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5207b, value : 32'h95059544},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5207c, value : 32'h1d0e4851},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5207d, value : 32'h29081104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5207e, value : 32'h78220101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5207f, value : 32'h22841c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52080, value : 32'hb5050004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52081, value : 32'hd027b10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52082, value : 32'h740cfe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52083, value : 32'h78e0c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52084, value : 32'hb5082b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52085, value : 32'hdc32c5e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52086, value : 32'hd2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52087, value : 32'h8c00bc9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52088, value : 32'h14f3b8c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52089, value : 32'h78a7908b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5208a, value : 32'h712ca900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5208b, value : 32'hc2900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5208c, value : 32'h90002311},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5208d, value : 32'h708daa80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5208e, value : 32'hdc4df012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5208f, value : 32'h8d2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52090, value : 32'h8c00bc9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52091, value : 32'h14f3b8c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52092, value : 32'h78a7908b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52093, value : 32'ha900718d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52094, value : 32'h10012c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52095, value : 32'h2311aa20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52096, value : 32'h722c9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52097, value : 32'hf208710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52098, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52099, value : 32'hab201228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5209a, value : 32'h700ca880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5209b, value : 32'h78e0c4c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5209c, value : 32'h700821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5209d, value : 32'h7de07014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5209e, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5209f, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a0, value : 32'hc02078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a1, value : 32'ha1007104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a2, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a3, value : 32'hf015122c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a4, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a5, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a6, value : 32'h50080f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a7, value : 32'hd10811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a8, value : 32'h811900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520a9, value : 32'h1900f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520aa, value : 32'hf0040041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ab, value : 32'h11900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ac, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ad, value : 32'h8820122e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ae, value : 32'h8801aa20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520af, value : 32'hab007fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b0, value : 32'h883c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b1, value : 32'h45080030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b2, value : 32'h71021600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b3, value : 32'h148000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b4, value : 32'hcc41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b5, value : 32'hc320001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b6, value : 32'hd8fffe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b7, value : 32'h8676d09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b8, value : 32'h120d01d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520b9, value : 32'h120c3083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ba, value : 32'h120d3604},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520bb, value : 32'h20253605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520bc, value : 32'hf0080000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520bd, value : 32'hf010f00b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520be, value : 32'hf018f013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520bf, value : 32'hf024f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c0, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c1, value : 32'h300cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c2, value : 32'h700cf022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c3, value : 32'hce41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c4, value : 32'hf01e0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c5, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c6, value : 32'h300cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c7, value : 32'h700cf018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c8, value : 32'hd041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520c9, value : 32'hf0140003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ca, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520cb, value : 32'h300d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520cc, value : 32'h120bf00e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520cd, value : 32'h41c33082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ce, value : 32'h400d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520cf, value : 32'hfc2f0aaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d0, value : 32'hc6c2700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d1, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d2, value : 32'h300d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d3, value : 32'h43804260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d4, value : 32'hfc2f0a96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d5, value : 32'h140240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d6, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d7, value : 32'h43cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d8, value : 32'h242f28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520d9, value : 32'h201f12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520da, value : 32'h7b8a02c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520db, value : 32'h108b2b41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520dc, value : 32'h2c1211f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520dd, value : 32'h184229f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520de, value : 32'h60386078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520df, value : 32'h42c36058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e0, value : 32'h1a468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e1, value : 32'h8012256},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e2, value : 32'h78356029},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e3, value : 32'h61116a2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e4, value : 32'h4a306052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e5, value : 32'h71047230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e6, value : 32'h20ca7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e7, value : 32'h78e00025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e8, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520e9, value : 32'hc1a6b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ea, value : 32'h16004608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520eb, value : 32'h80007100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ec, value : 32'h4528000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ed, value : 32'hc3414358},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ee, value : 32'h781dc043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ef, value : 32'h87812044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f0, value : 32'hc045710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f1, value : 32'hc042d810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f2, value : 32'h90df207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f3, value : 32'h700c00b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f4, value : 32'hf003c045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f5, value : 32'h208ac142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f6, value : 32'hb6010004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f7, value : 32'hae00d820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f8, value : 32'h81fc003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520f9, value : 32'hd8c8007e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520fa, value : 32'h8d409561},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520fb, value : 32'h21b41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520fc, value : 32'h121e0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520fd, value : 32'hb123705},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520fe, value : 32'h121ffe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h520ff, value : 32'h8d003704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52100, value : 32'hc2014363},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52101, value : 32'h95e14210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52102, value : 32'hc8e41e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52103, value : 32'h41f1fdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52104, value : 32'hc0034010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52105, value : 32'h7e081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52106, value : 32'h9561d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52107, value : 32'h41c38d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52108, value : 32'h4021c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52109, value : 32'h400240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5210a, value : 32'hfe6f0ade},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5210b, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5210c, value : 32'h7014c002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5210d, value : 32'h7216f2bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5210e, value : 32'h250174},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5210f, value : 32'hc002746e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52110, value : 32'h70ce8de0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52111, value : 32'hb82295a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52112, value : 32'h1410c044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52113, value : 32'h22003015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52114, value : 32'h240a24c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52115, value : 32'h210a2440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52116, value : 32'h20533400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52117, value : 32'h22020150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52118, value : 32'hd1124c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52119, value : 32'h20531521},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5211a, value : 32'hf1b0151},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5211b, value : 32'h70ee1460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5211c, value : 32'h4022c201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5211d, value : 32'hc224182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5211e, value : 32'h4363fdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5211f, value : 32'h15210d0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52120, value : 32'hf254710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52121, value : 32'hc2011400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52122, value : 32'h41824002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52123, value : 32'hfdaf0c0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52124, value : 32'hf154363},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52125, value : 32'h81f2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52126, value : 32'h47100664},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52127, value : 32'h220a474a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52128, value : 32'hf00b2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52129, value : 32'ha640270c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5212a, value : 32'h148627ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5212b, value : 32'h244622ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5212c, value : 32'h270af743},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5212d, value : 32'h24002640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5212e, value : 32'h240224c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5212f, value : 32'h205324d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52130, value : 32'h21530218},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52131, value : 32'h77522211},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52132, value : 32'h944125cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52133, value : 32'hd21f405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52134, value : 32'h700e1621},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52135, value : 32'hc201f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52136, value : 32'h41224042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52137, value : 32'hfdaf0bba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52138, value : 32'h40104363},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52139, value : 32'h25cc7752},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5213a, value : 32'hf2119601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5213b, value : 32'h4042c201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5213c, value : 32'hba64103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5213d, value : 32'h4363fdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5213e, value : 32'h20050813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5213f, value : 32'h5e40819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52140, value : 32'h2600210a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52141, value : 32'h4010458a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52142, value : 32'h200cf00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52143, value : 32'h25caa5c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52144, value : 32'hf7461506},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52145, value : 32'h2500210a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52146, value : 32'h25c0200a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52147, value : 32'h26610817},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52148, value : 32'h30141410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52149, value : 32'hf547262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5214a, value : 32'h2542f204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5214b, value : 32'hf0032054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5214c, value : 32'hc003708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5214d, value : 32'h7e082d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5214e, value : 32'h2507252f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5214f, value : 32'h41c3d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52150, value : 32'h7021d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52151, value : 32'h434242c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52152, value : 32'h440240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52153, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52154, value : 32'h400260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52155, value : 32'h4c0270a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52156, value : 32'hfe6f09ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52157, value : 32'h35401c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52158, value : 32'h8178e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52159, value : 32'hd170481},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5215a, value : 32'h96012010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5215b, value : 32'h440080f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5215c, value : 32'h2500250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5215d, value : 32'hdfdf012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5215e, value : 32'h1410a011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5215f, value : 32'h202f3015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52160, value : 32'h431084c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52161, value : 32'h716ef404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52162, value : 32'h2500250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52163, value : 32'h12079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52164, value : 32'h2005c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52165, value : 32'hf20c807e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52166, value : 32'hc00271c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52167, value : 32'ha000260c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52168, value : 32'h14441e02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52169, value : 32'hffe506aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5216a, value : 32'h14821e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5216b, value : 32'hc0a64002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5216c, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5216d, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5216e, value : 32'h44cbc0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5216f, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52170, value : 32'h8c204028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52171, value : 32'h7100244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52172, value : 32'h70ad70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52173, value : 32'h20a8708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52174, value : 32'h91b0240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52175, value : 32'h7185030f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52176, value : 32'h75c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52177, value : 32'h702c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52178, value : 32'h900345cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52179, value : 32'h706dc000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5217a, value : 32'h6892f015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5217b, value : 32'h10812800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5217c, value : 32'h79647d85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5217d, value : 32'h1f8c2505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5217e, value : 32'h9038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5217f, value : 32'h25059480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52180, value : 32'h903b1f8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52181, value : 32'h2406c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52182, value : 32'h7c6410cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52183, value : 32'h2c0179e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52184, value : 32'hc43108b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52185, value : 32'hb5200031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52186, value : 32'h708c1600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52187, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52188, value : 32'h1600ec88},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52189, value : 32'h8000708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5218a, value : 32'hec140040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5218b, value : 32'hbe0cde07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5218c, value : 32'h28007e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5218d, value : 32'h6e52108c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5218e, value : 32'h22057c64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5218f, value : 32'h90000f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52190, value : 32'h91200000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52191, value : 32'hf8d2205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52192, value : 32'hc0009003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52193, value : 32'h79857966},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52194, value : 32'h4061b520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52195, value : 32'h78e0c4c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52196, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52197, value : 32'hc1acb6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52198, value : 32'h4508c71c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52199, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5219a, value : 32'h148000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5219b, value : 32'h21c0230a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5219c, value : 32'h40384150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5219d, value : 32'h70ce708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5219e, value : 32'h31801c28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5219f, value : 32'h31401c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a0, value : 32'h31001c24},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a1, value : 32'h13e081b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a2, value : 32'h1600c348},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a3, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a4, value : 32'h80f001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a5, value : 32'h71ce003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a6, value : 32'h540086e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a7, value : 32'h97c44610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a8, value : 32'h8336d0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521a9, value : 32'h17020175},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521aa, value : 32'hdfa1110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ab, value : 32'he815fe4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ac, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ad, value : 32'h8841122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ae, value : 32'ha1f8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521af, value : 32'h790f0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b0, value : 32'h27147104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b1, value : 32'h19241041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b2, value : 32'h790f0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b3, value : 32'h80450af3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b4, value : 32'hddbf003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b5, value : 32'h20789050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b6, value : 32'h731730cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b7, value : 32'h24ca4d19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b8, value : 32'hc0412261},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521b9, value : 32'h23922038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ba, value : 32'hcbec01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521bb, value : 32'hc04b0360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521bc, value : 32'hfcef0832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521bd, value : 32'h83ed8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521be, value : 32'h970efcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521bf, value : 32'h208a70d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c0, value : 32'h208a0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c1, value : 32'h43db2002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c2, value : 32'h1d09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c3, value : 32'h200220ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c4, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c5, value : 32'h211f28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c6, value : 32'h781b2001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c7, value : 32'h2000231f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c8, value : 32'h45cb70b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521c9, value : 32'h3dd09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ca, value : 32'h702f757f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521cb, value : 32'h45d3700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521cc, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521cd, value : 32'hc0436038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ce, value : 32'h209f4082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521cf, value : 32'hc1030184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d0, value : 32'h20006038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d1, value : 32'h80000f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d2, value : 32'h70c31a44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d3, value : 32'h1a468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d4, value : 32'h2050c047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d5, value : 32'hc0453000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d6, value : 32'hc044710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d7, value : 32'hc146720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d8, value : 32'h40c3c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521d9, value : 32'hc2cc9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521da, value : 32'h1030081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521db, value : 32'hfc7218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521dc, value : 32'h736db020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521dd, value : 32'h6441804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521de, value : 32'h819c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521df, value : 32'h976800b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e0, value : 32'hf009bb07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e1, value : 32'h716d706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e2, value : 32'h6441800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e3, value : 32'hf003b022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e4, value : 32'h15b7bb08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e5, value : 32'h15012086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e6, value : 32'h15002089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e7, value : 32'h784f2082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e8, value : 32'h1024095f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521e9, value : 32'he57702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ea, value : 32'h2714002e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521eb, value : 32'h28401001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ec, value : 32'h27050387},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ed, value : 32'h90040f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ee, value : 32'h91323ed4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ef, value : 32'h2105b90a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f0, value : 32'hb42002c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f1, value : 32'h21f4c108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f2, value : 32'he2b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f3, value : 32'h60782030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f4, value : 32'h10300817},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f5, value : 32'h21557910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f6, value : 32'h218a0800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f7, value : 32'h208c0fcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f8, value : 32'hf7c98fcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521f9, value : 32'h218cf008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521fa, value : 32'h702c8002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521fb, value : 32'h2080f784},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521fc, value : 32'h4100003e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521fd, value : 32'h3402705},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521fe, value : 32'h7144b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h521ff, value : 32'habef1d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52200, value : 32'h4002fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52201, value : 32'hf2737056},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52202, value : 32'h208915b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52203, value : 32'h20881501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52204, value : 32'h15008f05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52205, value : 32'he830208b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52206, value : 32'hfc7278a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52207, value : 32'h2c7222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52208, value : 32'h108408c9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52209, value : 32'h108e094d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5220a, value : 32'hf80221f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5220b, value : 32'ha3c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5220c, value : 32'h611bc106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5220d, value : 32'h611cc107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5220e, value : 32'hc1014082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5220f, value : 32'h450835},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52210, value : 32'he988c100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52211, value : 32'h6812200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52212, value : 32'h811120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52213, value : 32'h400819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52214, value : 32'h7001248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52215, value : 32'h41814660},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52216, value : 32'h18020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52217, value : 32'h151904},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52218, value : 32'h1d41e04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52219, value : 32'h1842380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5221a, value : 32'h11842480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5221b, value : 32'hf1e77104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5221c, value : 32'hf1d67165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5221d, value : 32'h128c235f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5221e, value : 32'h222f7482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5221f, value : 32'h86d02c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52220, value : 32'h9631084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52221, value : 32'h468110ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52222, value : 32'hc0014182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52223, value : 32'h50957},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52224, value : 32'he888c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52225, value : 32'h6802200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52226, value : 32'h801020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52227, value : 32'h941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52228, value : 32'h187202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52229, value : 32'h7002248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5222a, value : 32'he209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5222b, value : 32'hf832000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5222c, value : 32'hc14c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5222d, value : 32'h20a8c00b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5222e, value : 32'h1b0601c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5222f, value : 32'h1bfc0014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52230, value : 32'h225f8005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52231, value : 32'h60f80500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52232, value : 32'h20300e0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52233, value : 32'h18347834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52234, value : 32'hf0060fc5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52235, value : 32'h23f4c309},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52236, value : 32'hb07a0083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52237, value : 32'h712471c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52238, value : 32'he40af1d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52239, value : 32'hf1cb7165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5223a, value : 32'hd06704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5223b, value : 32'h1500fc4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5223c, value : 32'h15012091},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5223d, value : 32'h262f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5223e, value : 32'h47d31447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5223f, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52240, value : 32'h3a40871},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52241, value : 32'h1700710d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52242, value : 32'h8652080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52243, value : 32'h2e4003ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52244, value : 32'h230a1397},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52245, value : 32'hc0012500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52246, value : 32'h20050b55},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52247, value : 32'he888c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52248, value : 32'h16802600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52249, value : 32'h801020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5224a, value : 32'h20000b41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5224b, value : 32'h22802b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5224c, value : 32'h20ca7317},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5224d, value : 32'h20050021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5224e, value : 32'h200505c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5224f, value : 32'hc10a06c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52250, value : 32'ha2c7034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52251, value : 32'h9000fda1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52252, value : 32'h1502265f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52253, value : 32'h7034c104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52254, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52255, value : 32'h2214be2c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52256, value : 32'hf20504c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52257, value : 32'hb1006159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52258, value : 32'h6159f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52259, value : 32'h41950},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5225a, value : 32'hf1d77166},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5225b, value : 32'hf1c37126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5225c, value : 32'h7724c102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5225d, value : 32'h7034c142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5225e, value : 32'h5ea702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5225f, value : 32'hc144ffe2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52260, value : 32'h20921500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52261, value : 32'h2487212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52262, value : 32'ha000210c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52263, value : 32'hd012a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52264, value : 32'h20811700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52265, value : 32'h84402111},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52266, value : 32'h225ef28d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52267, value : 32'h468a2296},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52268, value : 32'h7610c001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52269, value : 32'h6010a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5226a, value : 32'he888c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5226b, value : 32'h26802100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5226c, value : 32'h801020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5226d, value : 32'h10000ea1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5226e, value : 32'h2503215f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5226f, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52270, value : 32'h2314be2c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52271, value : 32'h60590382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52272, value : 32'h11506215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52273, value : 32'h8f050113},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52274, value : 32'h9724e82e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52275, value : 32'h9701db3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52276, value : 32'h97074831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52277, value : 32'h12904},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52278, value : 32'h41c37830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52279, value : 32'h2023e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5227a, value : 32'h20bc4200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5227b, value : 32'hbfa0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5227c, value : 32'h4050fbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5227d, value : 32'h2f81211f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5227e, value : 32'ha3c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5227f, value : 32'h6119c003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52280, value : 32'h209a40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52281, value : 32'h60380184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52282, value : 32'h4012015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52283, value : 32'hf802100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52284, value : 32'h1a448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52285, value : 32'hf822100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52286, value : 32'h1a468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52287, value : 32'h23650b33},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52288, value : 32'hfc7218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52289, value : 32'h51a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5228a, value : 32'hf016b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5228b, value : 32'h23640b29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5228c, value : 32'h79d46779},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5228d, value : 32'h82d911a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5228e, value : 32'hf81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5228f, value : 32'h2300ffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52290, value : 32'he0ff2340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52291, value : 32'h700cf70a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52292, value : 32'h51934},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52293, value : 32'hb0a0f00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52294, value : 32'h4c41a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52295, value : 32'hf1a671c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52296, value : 32'h2080781d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52297, value : 32'hb11a003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52298, value : 32'h78109728},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52299, value : 32'h75104d12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5229a, value : 32'h4c0200e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5229b, value : 32'h23832600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5229c, value : 32'h4b2a04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5229d, value : 32'h28047c6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5229e, value : 32'h23ca0040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5229f, value : 32'h7a101025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a0, value : 32'h2c8212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a1, value : 32'h80640ad1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a2, value : 32'h215f4081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a3, value : 32'h209f0181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a4, value : 32'h6119000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a5, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a6, value : 32'h6038c14c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a7, value : 32'hb0219721},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a8, value : 32'h90609721},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522a9, value : 32'hc50907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522aa, value : 32'h7165b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ab, value : 32'h1501f1ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ac, value : 32'h71462080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ad, value : 32'hc0acf168},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ae, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522af, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b0, value : 32'h47cbc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b1, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b2, value : 32'h240a8fc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b3, value : 32'h250a2180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b4, value : 32'h260a2140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b5, value : 32'h47702100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b6, value : 32'h41384058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b7, value : 32'h8f014110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b8, value : 32'h3840899},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522b9, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ba, value : 32'h880012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522bb, value : 32'h3ae0889},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522bc, value : 32'h1105704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522bd, value : 32'h700e2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522be, value : 32'h27f4e883},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522bf, value : 32'h265a2390},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c0, value : 32'h11051293},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c1, value : 32'he81d2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c2, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c3, value : 32'h791b28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c4, value : 32'h3002211f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c5, value : 32'h3041201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c6, value : 32'h78ccb822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c7, value : 32'h611a6159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c8, value : 32'h209a4042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522c9, value : 32'h621a0184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ca, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522cb, value : 32'h60591a44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522cc, value : 32'h91016215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522cd, value : 32'h345081b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ce, value : 32'h700c70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522cf, value : 32'hccaf009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d0, value : 32'h4062ff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d1, value : 32'h40624508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d2, value : 32'hff6f0cee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d3, value : 32'h60b941a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d4, value : 32'h24c22614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d5, value : 32'h7502793d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d6, value : 32'h71467102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d7, value : 32'h2514b220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d8, value : 32'hb1a024c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522d9, value : 32'h4012000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522da, value : 32'h24c02414},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522db, value : 32'ha977166},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522dc, value : 32'hb020a2b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522dd, value : 32'hf1b571c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522de, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522df, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e0, value : 32'h8901122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e1, value : 32'h71108920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e2, value : 32'h7cd20e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e3, value : 32'h29407822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e4, value : 32'h71040382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e5, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e6, value : 32'h30020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e7, value : 32'hf812205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e8, value : 32'h1d09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522e9, value : 32'h72c39100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ea, value : 32'h40000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522eb, value : 32'hb100e020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ec, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ed, value : 32'h343236f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ee, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ef, value : 32'h93000460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f0, value : 32'h208cda08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f1, value : 32'hd8088059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f2, value : 32'h2a520ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f3, value : 32'h9300b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f4, value : 32'h8059208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f5, value : 32'h20cad808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f6, value : 32'hb10102a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f7, value : 32'h208c9300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f8, value : 32'hd8088059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522f9, value : 32'h2a520ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522fa, value : 32'h9300b102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522fb, value : 32'h8059208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522fc, value : 32'h2a522ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522fd, value : 32'hb1437fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522fe, value : 32'hc1a2c3ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h522ff, value : 32'h42104728},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52300, value : 32'hc0d2055},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52301, value : 32'hf464020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52302, value : 32'h702cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52303, value : 32'h40424010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52304, value : 32'hcee702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52305, value : 32'hdacafbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52306, value : 32'h208a71cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52307, value : 32'hb5c20016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52308, value : 32'h20041ac2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52309, value : 32'hc15208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5230a, value : 32'h1600b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5230b, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5230c, value : 32'h20440009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5230d, value : 32'h710c8091},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5230e, value : 32'ha120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5230f, value : 32'h22431ac6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52310, value : 32'h2e00f22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52311, value : 32'h20021ac9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52312, value : 32'h22408d24},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52313, value : 32'hadc82403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52314, value : 32'h200d2178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52315, value : 32'h424240e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52316, value : 32'h71ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52317, value : 32'hfeef0d0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52318, value : 32'h12c546a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52319, value : 32'h22402081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5231a, value : 32'h22402202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5231b, value : 32'h40e12603},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5231c, value : 32'h71ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5231d, value : 32'hfeef0cf2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5231e, value : 32'h47cb46a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5231f, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52320, value : 32'h8f018fc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52321, value : 32'h3840841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52322, value : 32'h238d2214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52323, value : 32'hecec180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52324, value : 32'h9500fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52325, value : 32'hec69504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52326, value : 32'hc181fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52327, value : 32'haf2c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52328, value : 32'h712c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52329, value : 32'hfe2f0b16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5232a, value : 32'hb500c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5232b, value : 32'hae2c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5232c, value : 32'h712c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5232d, value : 32'hfe2f0b06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5232e, value : 32'hb504c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5232f, value : 32'h76108f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52330, value : 32'hf7a471c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52331, value : 32'h5000986},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52332, value : 32'h70148fc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52333, value : 32'h2040740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52334, value : 32'h20ca2413},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52335, value : 32'h204001e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52336, value : 32'h1ac72491},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52337, value : 32'h8f012002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52338, value : 32'h3a4085f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52339, value : 32'h13102e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5233a, value : 32'h265a70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5233b, value : 32'h2d401503},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5233c, value : 32'h22051202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5233d, value : 32'hc8090402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5233e, value : 32'h41c37a05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5233f, value : 32'h9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52340, value : 32'h4402205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52341, value : 32'h4c22205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52342, value : 32'hb8027342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52343, value : 32'h78257bb4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52344, value : 32'h1051000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52345, value : 32'h1b206a12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52346, value : 32'h78250144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52347, value : 32'h1041000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52348, value : 32'h1b70740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52349, value : 32'h41c30104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5234a, value : 32'h401c9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5234b, value : 32'h9da42c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5234c, value : 32'h43a1fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5234d, value : 32'hdb771a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5234e, value : 32'h71c59254},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5234f, value : 32'hc7cef1d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52350, value : 32'h40c3c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52351, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52352, value : 32'hc8098880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52353, value : 32'h7885bc0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52354, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52355, value : 32'hfd80003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52356, value : 32'h5200bd6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52357, value : 32'hc809702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52358, value : 32'h6c127c05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52359, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5235a, value : 32'h364900c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5235b, value : 32'h7fe0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5235c, value : 32'h51800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5235d, value : 32'hd9ffd838},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5235e, value : 32'h1803b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5235f, value : 32'h18fc0052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52360, value : 32'h18018042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52361, value : 32'h18160052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52362, value : 32'h18010052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52363, value : 32'ha8200052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52364, value : 32'h7fe0a823},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52365, value : 32'h78e0a824},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52366, value : 32'hd9ffd83a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52367, value : 32'h1803b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52368, value : 32'h18fc0052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52369, value : 32'h18018042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5236a, value : 32'h18160052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5236b, value : 32'h18010052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5236c, value : 32'ha8200052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5236d, value : 32'h7fe0a823},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5236e, value : 32'h78e0a824},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5236f, value : 32'h200ac2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52370, value : 32'h47682100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52371, value : 32'h45284648},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52372, value : 32'h135080b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52373, value : 32'hba0e4200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52374, value : 32'ha0ff00d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52375, value : 32'h700c03f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52376, value : 32'hba0eda1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52377, value : 32'h41c3f008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52378, value : 32'h10030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52379, value : 32'hfbcf0802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5237a, value : 32'hba92704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5237b, value : 32'h900040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5237c, value : 32'h22053a90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5237d, value : 32'h74040001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5237e, value : 32'h2205b1a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5237f, value : 32'h74040001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52380, value : 32'h2205b1c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52381, value : 32'h74040001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52382, value : 32'hb1e07845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52383, value : 32'h4041800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52384, value : 32'h78e0c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52385, value : 32'h4110c2ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52386, value : 32'h230a4040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52387, value : 32'h220a2140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52388, value : 32'h45682100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52389, value : 32'hfeaf0bca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5238a, value : 32'h46084030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5238b, value : 32'hfeaf0bc2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5238c, value : 32'h470840a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5238d, value : 32'hfeaf0bba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5238e, value : 32'h45084042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5238f, value : 32'hfeaf0bb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52390, value : 32'h9214062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52391, value : 32'h92d2090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52392, value : 32'h9472050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52393, value : 32'h42222031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52394, value : 32'h901c42c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52395, value : 32'h41c3006c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52396, value : 32'hf8a89007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52397, value : 32'hf011b2c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52398, value : 32'h901c42c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52399, value : 32'hb2c000ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5239a, value : 32'h900741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5239b, value : 32'hf009f928},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5239c, value : 32'h901c42c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5239d, value : 32'hb2c000ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5239e, value : 32'h900741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5239f, value : 32'hb2e2f8e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a0, value : 32'hb102b1a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a1, value : 32'h84041ad4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a2, value : 32'h840419d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a3, value : 32'h41c3c6ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a4, value : 32'h1002f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a5, value : 32'hfbaf0f52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a6, value : 32'hc6ce700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a7, value : 32'h45cbc5e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a8, value : 32'h6c901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523a9, value : 32'h10141d04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523aa, value : 32'h900744cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ab, value : 32'h1d3cf8a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ac, value : 32'h1c041054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ad, value : 32'h1c3c1094},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ae, value : 32'h1d0410d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523af, value : 32'hb5201014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b0, value : 32'h10941c04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b1, value : 32'hb51eb460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b2, value : 32'h10441d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b3, value : 32'h1c40b45e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b4, value : 32'hc4c210c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b5, value : 32'h1600c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b6, value : 32'h90307100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b7, value : 32'h45cb0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b8, value : 32'h4fcc8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523b9, value : 32'h1a11dab0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ba, value : 32'h206d3003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523bb, value : 32'h40c30081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523bc, value : 32'h4a88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523bd, value : 32'h40a1a820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523be, value : 32'hfbaf0a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523bf, value : 32'h42c3702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c0, value : 32'hfffc7fff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c1, value : 32'h10802504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c2, value : 32'h2000b822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c3, value : 32'h50f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c4, value : 32'h12688000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c5, value : 32'h20790600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c6, value : 32'h1a680000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c7, value : 32'h1a090058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c8, value : 32'hc6c23002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523c9, value : 32'hb7ac3ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ca, value : 32'hc1a1fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523cb, value : 32'h800040d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523cc, value : 32'h205410dc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523cd, value : 32'h70cd280f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ce, value : 32'h254270ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523cf, value : 32'h8111700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d0, value : 32'h160001d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d1, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d2, value : 32'he8130131},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d3, value : 32'h14032532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d4, value : 32'h1700700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d5, value : 32'h762c1084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d6, value : 32'h254a704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d7, value : 32'hb8603c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d8, value : 32'h70ccfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523d9, value : 32'hd922700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523da, value : 32'hfc6f0e6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523db, value : 32'h71a5704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523dc, value : 32'h98f40dcb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523dd, value : 32'h700c71e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523de, value : 32'hfc6f0b1a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523df, value : 32'hdd25712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e0, value : 32'hbd9f714e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e1, value : 32'h702c722e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e2, value : 32'h8d40720e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e3, value : 32'h7a058d1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e4, value : 32'h20402a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e5, value : 32'h200fb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e6, value : 32'h7f4b004f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e7, value : 32'he4ef21b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e8, value : 32'h40c10060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523e9, value : 32'hafae817},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ea, value : 32'h252ffc0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523eb, value : 32'h700c03c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ec, value : 32'h704c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ed, value : 32'h244adbd0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ee, value : 32'hb2a0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ef, value : 32'h70ccfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f0, value : 32'hd922700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f1, value : 32'hfc6f0e12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f2, value : 32'h700c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f3, value : 32'hfc6f0ac6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f4, value : 32'h208d712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f5, value : 32'h712c277f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f6, value : 32'h25ff218d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f7, value : 32'hd98271cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f8, value : 32'hb99f70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523f9, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523fa, value : 32'h712e1228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523fb, value : 32'h4801101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523fc, value : 32'h140206c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523fd, value : 32'he002045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523fe, value : 32'h8900c060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h523ff, value : 32'h140206c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52400, value : 32'he002045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52401, value : 32'h30021c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52402, value : 32'h206c8901},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52403, value : 32'h20450140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52404, value : 32'h1c020e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52405, value : 32'h89023002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52406, value : 32'h140206c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52407, value : 32'he002045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52408, value : 32'h30021c03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52409, value : 32'h790f700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5240a, value : 32'hb50979},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5240b, value : 32'he906af00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5240c, value : 32'he8888d1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5240d, value : 32'hf034710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5240e, value : 32'h70148d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5240f, value : 32'hf230700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52410, value : 32'h20402900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52411, value : 32'hfeaf0842},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52412, value : 32'ha56780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52413, value : 32'h702cfc0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52414, value : 32'h8d60720e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52415, value : 32'h7b058d1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52416, value : 32'h20402900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52417, value : 32'h200fb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52418, value : 32'h7a6b0042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52419, value : 32'h8f60f20f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5241a, value : 32'h252fc080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5241b, value : 32'h704c0087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5241c, value : 32'h440244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5241d, value : 32'h787470cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5241e, value : 32'h700c602b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5241f, value : 32'hfc6f0a66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52420, value : 32'h208d762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52421, value : 32'h712c2a7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52422, value : 32'hd922700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52423, value : 32'hfc6f0d4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52424, value : 32'h700c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52425, value : 32'hfc6f09fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52426, value : 32'h8f00712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52427, value : 32'hf1c57104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52428, value : 32'hfe6f0fe6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52429, value : 32'hb7c0730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5242a, value : 32'h78e0c7cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5242b, value : 32'hf16c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5242c, value : 32'h208a00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5242d, value : 32'h7910041f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5242e, value : 32'hd1e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5242f, value : 32'h704cfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52430, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52431, value : 32'h4508c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52432, value : 32'hb813d841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52433, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52434, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52435, value : 32'ha0e70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52436, value : 32'h70ccfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52437, value : 32'hfc4f0cb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52438, value : 32'hd90740a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52439, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5243a, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5243b, value : 32'hfc6f09f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5243c, value : 32'hc8670cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5243d, value : 32'h40a1fc4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5243e, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5243f, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52440, value : 32'h9e270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52441, value : 32'h70ccfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52442, value : 32'hd907d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52443, value : 32'h744cb893},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52444, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52445, value : 32'h9ce70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52446, value : 32'h70ccfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52447, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52448, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52449, value : 32'h8a40122d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5244a, value : 32'h42223c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5244b, value : 32'h16007854},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5244c, value : 32'h80007082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5244d, value : 32'h22110121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5244e, value : 32'h21448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5244f, value : 32'h20f90040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52450, value : 32'h7fe00022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52451, value : 32'h2120f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52452, value : 32'h4608c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52453, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52454, value : 32'h8800122d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52455, value : 32'h203c4528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52456, value : 32'hc920040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52457, value : 32'h41c10060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52458, value : 32'h710c7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52459, value : 32'h38120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5245a, value : 32'hffe10fb8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5245b, value : 32'hc6c441a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5245c, value : 32'h923682b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5245d, value : 32'h71140175},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5245e, value : 32'h71011600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5245f, value : 32'h148000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52460, value : 32'h710cb9e3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52461, value : 32'h21047de0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52462, value : 32'hf80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52463, value : 32'hb82e4000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52464, value : 32'h700cf003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52465, value : 32'h7ee0f3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52466, value : 32'h4220c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52467, value : 32'h2144b923},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52468, value : 32'hbac50601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52469, value : 32'h81006119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5246a, value : 32'hfbaf0b22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5246b, value : 32'hb8c08121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5246c, value : 32'h7fe0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5246d, value : 32'h2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5246e, value : 32'h2482c3ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5246f, value : 32'h45083708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52470, value : 32'h9c2c087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52471, value : 32'h41a1ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52472, value : 32'hc18240a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52473, value : 32'hfd6f087e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52474, value : 32'h31c22440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52475, value : 32'hc7cce802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52476, value : 32'h30801407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52477, value : 32'hb00811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52478, value : 32'h80f72cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52479, value : 32'h704e00f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5247a, value : 32'hf00370cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5247b, value : 32'h702e714e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5247c, value : 32'hc080c182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5247d, value : 32'h42a179d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5247e, value : 32'hffaf09aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5247f, value : 32'h80fc387},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52480, value : 32'hc7200444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52481, value : 32'h14024110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52482, value : 32'h76523110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52483, value : 32'hf63277c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52484, value : 32'ha03009c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52485, value : 32'h1d82750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52486, value : 32'h2580141c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52487, value : 32'h700c1084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52488, value : 32'hc7ccade0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52489, value : 32'hc1a2c3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5248a, value : 32'h70ad4708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5248b, value : 32'h800146cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5248c, value : 32'hc5414d84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5248d, value : 32'h71080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5248e, value : 32'hd864c540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5248f, value : 32'hf066b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52490, value : 32'hb606d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52491, value : 32'h80ff062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52492, value : 32'he8890050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52493, value : 32'hb808d87f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52494, value : 32'hd87ff003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52495, value : 32'hc040b810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52496, value : 32'hd9fbf006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52497, value : 32'hb8a700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52498, value : 32'hb910fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52499, value : 32'h10710f0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5249a, value : 32'h26f44e1c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5249b, value : 32'hf0041340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5249c, value : 32'h34020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5249d, value : 32'hb0eb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5249e, value : 32'h7810fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5249f, value : 32'hd907d841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a0, value : 32'hda08b813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a1, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a2, value : 32'h85a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a3, value : 32'h70ccfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a4, value : 32'h742c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a5, value : 32'hfc6f0b42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a6, value : 32'hc080714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a7, value : 32'ha9a41e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a8, value : 32'h724cfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524a9, value : 32'hd914700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524aa, value : 32'hfc6f0b2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ab, value : 32'h706c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ac, value : 32'h4060d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ad, value : 32'hb892744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ae, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524af, value : 32'hfc6f0826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b0, value : 32'h160070cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b1, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b2, value : 32'h811000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b3, value : 32'h700c003e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b4, value : 32'hb06d914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b5, value : 32'h714cfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b6, value : 32'hd907d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b7, value : 32'hda08b893},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b8, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524b9, value : 32'hffe70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ba, value : 32'h70ccfc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524bb, value : 32'hfbcf0f9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524bc, value : 32'h13412614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524bd, value : 32'h10710f0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524be, value : 32'hb1016849},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524bf, value : 32'hb14c71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c0, value : 32'hb107f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c1, value : 32'hb15271a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c2, value : 32'h90b40d3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c3, value : 32'hc7c678b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c4, value : 32'h702cc2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c5, value : 32'h4508da4b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c6, value : 32'hfb6f0de6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c7, value : 32'h90e2055},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c8, value : 32'h704cd95a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524c9, value : 32'h1104b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ca, value : 32'had010480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524cb, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524cc, value : 32'h1104ad02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524cd, value : 32'had030480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ce, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524cf, value : 32'h1104ad0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d0, value : 32'had0b0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d1, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d2, value : 32'h1104ad0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d3, value : 32'had0d0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d4, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d5, value : 32'h1104ad0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d6, value : 32'had0f0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d7, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d8, value : 32'h1104ad10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524d9, value : 32'had110480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524da, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524db, value : 32'h1104ad12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524dc, value : 32'had130480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524dd, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524de, value : 32'h1104ad14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524df, value : 32'had150480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e0, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e1, value : 32'h1104ad16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e2, value : 32'had180480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e3, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e4, value : 32'h1104ad19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e5, value : 32'had1a0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e6, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e7, value : 32'h1104ad1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e8, value : 32'had1c0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524e9, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ea, value : 32'h1104ad1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524eb, value : 32'had1f0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ec, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ed, value : 32'h10021d20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ee, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ef, value : 32'h10021d21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f0, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f1, value : 32'h10021d22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f2, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f3, value : 32'h10021d25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f4, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f5, value : 32'h10021d28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f6, value : 32'h4801108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f7, value : 32'h10021d29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f8, value : 32'h10821d2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524f9, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524fa, value : 32'h10021d3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524fb, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524fc, value : 32'h10021d45},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524fd, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524fe, value : 32'h10021d46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h524ff, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52500, value : 32'h10021d47},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52501, value : 32'h84801179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52502, value : 32'h10021d48},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52503, value : 32'h80118b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52504, value : 32'h10021d49},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52505, value : 32'h80118f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52506, value : 32'h10021d4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52507, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52508, value : 32'h10021d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52509, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5250a, value : 32'h10021d4d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5250b, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5250c, value : 32'h10021d4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5250d, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5250e, value : 32'h10021d55},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5250f, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52510, value : 32'h10021d56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52511, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52512, value : 32'h10021d57},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52513, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52514, value : 32'h10021d58},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52515, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52516, value : 32'h10021d59},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52517, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52518, value : 32'h10021d5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52519, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5251a, value : 32'h10021d5b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5251b, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5251c, value : 32'h10021d5c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5251d, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5251e, value : 32'h10021d5d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5251f, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52520, value : 32'h10021d5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52521, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52522, value : 32'h10021d5f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52523, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52524, value : 32'h10021d60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52525, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52526, value : 32'h10021d61},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52527, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52528, value : 32'h10021d63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52529, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5252a, value : 32'h10021d64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5252b, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5252c, value : 32'h10021d65},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5252d, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5252e, value : 32'h10021d66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5252f, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52530, value : 32'h10021d67},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52531, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52532, value : 32'h10021d69},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52533, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52534, value : 32'h10021d6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52535, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52536, value : 32'h10021d6b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52537, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52538, value : 32'h10021d6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52539, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5253a, value : 32'h10021d6d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5253b, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5253c, value : 32'h10021d70},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5253d, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5253e, value : 32'h10021d73},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5253f, value : 32'h4801108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52540, value : 32'h10021d74},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52541, value : 32'h10821d79},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52542, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52543, value : 32'h10021d85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52544, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52545, value : 32'h1104ae00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52546, value : 32'h1d910480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52547, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52548, value : 32'h1d920480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52549, value : 32'h11791002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5254a, value : 32'h1d938480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5254b, value : 32'h118b1002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5254c, value : 32'hae040080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5254d, value : 32'h80118f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5254e, value : 32'h10021d95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5254f, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52550, value : 32'h10021d97},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52551, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52552, value : 32'h1104ae08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52553, value : 32'h1d990480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52554, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52555, value : 32'hae100480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52556, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52557, value : 32'h10021da1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52558, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52559, value : 32'h10021da2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5255a, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5255b, value : 32'h10021da3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5255c, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5255d, value : 32'h1104ae14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5255e, value : 32'h1da50480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5255f, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52560, value : 32'h1da60480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52561, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52562, value : 32'h1da70480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52563, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52564, value : 32'hae180480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52565, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52566, value : 32'h10021da9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52567, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52568, value : 32'h10021daa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52569, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5256a, value : 32'h10021dab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5256b, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5256c, value : 32'h1104ae1c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5256d, value : 32'h1dae0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5256e, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5256f, value : 32'h1daf0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52570, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52571, value : 32'h1e200480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52572, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52573, value : 32'h1db10480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52574, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52575, value : 32'h1db20480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52576, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52577, value : 32'h1e240480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52578, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52579, value : 32'h1db50480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5257a, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5257b, value : 32'h1db60480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5257c, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5257d, value : 32'h1db70480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5257e, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5257f, value : 32'h1e280480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52580, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52581, value : 32'h1dbb0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52582, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52583, value : 32'h1dbe0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52584, value : 32'h11081002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52585, value : 32'h1dbf0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52586, value : 32'h1e341002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52587, value : 32'h11041082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52588, value : 32'h1e400480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52589, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5258a, value : 32'h1ddb0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5258b, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5258c, value : 32'h1e4c0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5258d, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5258e, value : 32'h1ddd0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5258f, value : 32'h11791002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52590, value : 32'h1dde8480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52591, value : 32'h118b1002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52592, value : 32'h1ddf0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52593, value : 32'h118f1002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52594, value : 32'h1e500080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52595, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52596, value : 32'h1de20480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52597, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52598, value : 32'h1de30480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52599, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5259a, value : 32'h1e540480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5259b, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5259c, value : 32'h1deb0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5259d, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5259e, value : 32'h1e5c0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5259f, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a0, value : 32'h1ded0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a1, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a2, value : 32'h1dee0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a3, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a4, value : 32'h1def0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a5, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a6, value : 32'h1e600480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a7, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a8, value : 32'h1df10480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525a9, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525aa, value : 32'h1df20480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ab, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ac, value : 32'h1df30480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ad, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ae, value : 32'h1e640480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525af, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b0, value : 32'h1df50480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b1, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b2, value : 32'h1df60480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b3, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b4, value : 32'h1df70480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b5, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b6, value : 32'h1df90480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b7, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b8, value : 32'h1dfa0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525b9, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ba, value : 32'h1dfb0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525bb, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525bc, value : 32'h1e6c0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525bd, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525be, value : 32'h1dfd0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525bf, value : 32'h11041002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c0, value : 32'h1dff0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c1, value : 32'h25561002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c2, value : 32'h11041800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c3, value : 32'ha8600483},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c4, value : 32'h238043a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c5, value : 32'h11040044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c6, value : 32'hab000480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c7, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c8, value : 32'h1104ab01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525c9, value : 32'hab020480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ca, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525cb, value : 32'h1104ab05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525cc, value : 32'hab080480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525cd, value : 32'h4801108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ce, value : 32'hab4eab09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525cf, value : 32'h4801104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d0, value : 32'h1104ab1a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d1, value : 32'h1b250480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d2, value : 32'h11040002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d3, value : 32'h1b260480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d4, value : 32'h25560002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d5, value : 32'h11041940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d6, value : 32'ha8400482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d7, value : 32'h1b288900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d8, value : 32'h89040002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525d9, value : 32'h21b29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525da, value : 32'h1b2a8908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525db, value : 32'hc6c40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525dc, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525dd, value : 32'h256fb6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525de, value : 32'h8d001243},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525df, value : 32'h17e084f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e0, value : 32'h42c3c1ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e1, value : 32'h349018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e2, value : 32'h5001204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e3, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e4, value : 32'h1902018c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e5, value : 32'h12040014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e6, value : 32'h19020500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e7, value : 32'h12040014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e8, value : 32'h19020500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525e9, value : 32'h12e00014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ea, value : 32'hb1008500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525eb, value : 32'h6872c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ec, value : 32'h802305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ed, value : 32'hb1039000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ee, value : 32'h3002242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ef, value : 32'h90007865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f0, value : 32'h6a0cb101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f1, value : 32'h90007865},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f2, value : 32'hc08bb102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f3, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f4, value : 32'h916063d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f5, value : 32'h764cfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f6, value : 32'haf2c08b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f7, value : 32'h762c0520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f8, value : 32'hd9258d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525f9, value : 32'hb99fb8c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525fa, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525fb, value : 32'h22c9008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525fc, value : 32'h42c38900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525fd, value : 32'h1c8901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525fe, value : 32'h891bb200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h525ff, value : 32'h11f4b202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52600, value : 32'he8968080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52601, value : 32'h300095e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52602, value : 32'h2042c805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52603, value : 32'hf210803c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52604, value : 32'h20a8700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52605, value : 32'h20050380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52606, value : 32'h90040f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52607, value : 32'h9220028c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52608, value : 32'h70c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52609, value : 32'h21444000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5260a, value : 32'hb2200301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5260b, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5260c, value : 32'h68000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5260d, value : 32'hf85082b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5260e, value : 32'hc810000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5260f, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52610, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52611, value : 32'h20049024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52612, value : 32'h8179800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52613, value : 32'h41c30013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52614, value : 32'hff810000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52615, value : 32'h902c40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52616, value : 32'hb0200c98},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52617, value : 32'h41c3b022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52618, value : 32'hc98902c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52619, value : 32'h91229100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5261a, value : 32'hb8e07825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5261b, value : 32'hfc810fc4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5261c, value : 32'hb7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5261d, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5261e, value : 32'h11d8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5261f, value : 32'h3647014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52620, value : 32'h16000002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52621, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52622, value : 32'h701400f3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52623, value : 32'h10336},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52624, value : 32'h702e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52625, value : 32'h1e00b88c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52626, value : 32'h90077444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52627, value : 32'h47cbc3e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52628, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52629, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5262a, value : 32'hc3649007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5262b, value : 32'h6892c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5262c, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5262d, value : 32'h270001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5262e, value : 32'h1f832405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5262f, value : 32'h83c9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52630, value : 32'h24059320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52631, value : 32'h90071f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52632, value : 32'h2104c83c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52633, value : 32'hf81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52634, value : 32'h2185ff78},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52635, value : 32'hb2200182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52636, value : 32'h1f812405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52637, value : 32'hc09c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52638, value : 32'hb802c04a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52639, value : 32'hc14478e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5263a, value : 32'h9020c047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5263b, value : 32'hb9a0c004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5263c, value : 32'h1600b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5263d, value : 32'h90047100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5263e, value : 32'hb8a00ab0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5263f, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52640, value : 32'hcab09007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52641, value : 32'h20459300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52642, value : 32'hb2a0014d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52643, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52644, value : 32'h88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52645, value : 32'h1002079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52646, value : 32'h2040b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52647, value : 32'h2b40030b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52648, value : 32'hde61240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52649, value : 32'h20960120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5264a, value : 32'hc8090208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5264b, value : 32'h46cbbda0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5264c, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5264d, value : 32'h22056852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5264e, value : 32'h90070f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5264f, value : 32'hb1a0c83c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52650, value : 32'hae208e22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52651, value : 32'h16048e23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52652, value : 32'h218c1092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52653, value : 32'h22ca8fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52654, value : 32'hae212022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52655, value : 32'h21012250},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52656, value : 32'h34401c0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52657, value : 32'h1c08b90e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52658, value : 32'h79453440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52659, value : 32'h34401c04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5265a, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5265b, value : 32'h8249004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5265c, value : 32'h793b9120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5265d, value : 32'hf872184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5265e, value : 32'h231f7124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5265f, value : 32'h21551041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52660, value : 32'hc1450dc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52661, value : 32'hf812205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52662, value : 32'h1909038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52663, value : 32'hc1499120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52664, value : 32'hb962c181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52665, value : 32'h202fc148},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52666, value : 32'h42c32487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52667, value : 32'ha809004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52668, value : 32'h23132840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52669, value : 32'h4c02005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5266a, value : 32'h21056832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5266b, value : 32'h90000080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5266c, value : 32'hb3024383},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5266d, value : 32'h21056a04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5266e, value : 32'h74040002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5266f, value : 32'hb3439240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52670, value : 32'h22105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52671, value : 32'h74049240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52672, value : 32'h2105b344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52673, value : 32'h92400002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52674, value : 32'hb3457404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52675, value : 32'h208a7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52676, value : 32'h91200fcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52677, value : 32'h2840b307},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52678, value : 32'hb3262380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52679, value : 32'hf8d2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5267a, value : 32'hab09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5267b, value : 32'h9520c046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5267c, value : 32'h214f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5267d, value : 32'hb9a0b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5267e, value : 32'hc006b520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5267f, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52680, value : 32'h3549004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52681, value : 32'hc0099020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52682, value : 32'h25f0807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52683, value : 32'h140c793d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52684, value : 32'h252f3107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52685, value : 32'h140a2048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52686, value : 32'h740c3106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52687, value : 32'h31031404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52688, value : 32'h5a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52689, value : 32'h14080007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5268a, value : 32'h42023105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5268b, value : 32'h311b1406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5268c, value : 32'h6c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5268d, value : 32'hfdaf0cd2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5268e, value : 32'h35401c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5268f, value : 32'h26c0255f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52690, value : 32'h30161420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52691, value : 32'h70ee708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52692, value : 32'h9012885},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52693, value : 32'h20192502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52694, value : 32'h5582000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52695, value : 32'h21011602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52696, value : 32'h71021600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52697, value : 32'h68000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52698, value : 32'ha11783b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52699, value : 32'hf85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5269a, value : 32'hd2d0c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5269b, value : 32'hf0202005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5269c, value : 32'h5440825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5269d, value : 32'h20300f19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5269e, value : 32'h30402302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5269f, value : 32'h21001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a0, value : 32'h8154910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a1, value : 32'h8113002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a2, value : 32'hf0120642},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a3, value : 32'h30020809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a4, value : 32'h64308e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a5, value : 32'h2779d95d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a6, value : 32'hb4e2100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a7, value : 32'hb910fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a8, value : 32'h72c671e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526a9, value : 32'ha1740fb1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526aa, value : 32'h758e7186},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ab, value : 32'h2305c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ac, value : 32'h12f86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ad, value : 32'h2005020f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ae, value : 32'h200504c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526af, value : 32'hb9020180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b0, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b1, value : 32'hab49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b2, value : 32'h5041900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b3, value : 32'h1e00d99c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b4, value : 32'h90077044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b5, value : 32'hc10ac364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b6, value : 32'h4c12105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b7, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b8, value : 32'h130003cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526b9, value : 32'h214f1109},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ba, value : 32'h1b001001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526bb, value : 32'h68321044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526bc, value : 32'h110079e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526bd, value : 32'h206c0108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526be, value : 32'hb8801040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526bf, value : 32'hc0ab100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c0, value : 32'hc0050120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c1, value : 32'h10002150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c2, value : 32'h10022050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c3, value : 32'h10041b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c4, value : 32'h2005c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c5, value : 32'hb9020181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c6, value : 32'hb14079e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c7, value : 32'h224f9540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c8, value : 32'hb5200001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526c9, value : 32'h4c12005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ca, value : 32'hbaa0b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526cb, value : 32'h2105b540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526cc, value : 32'h90040f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526cd, value : 32'hc1060abc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ce, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526cf, value : 32'h3589004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d0, value : 32'hb2209120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d1, value : 32'h80d8e23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d2, value : 32'h218c2065},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d3, value : 32'hf4108fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d4, value : 32'h20610813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d5, value : 32'h8e258e44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d6, value : 32'h72304250},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d7, value : 32'h206d21ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d8, value : 32'h815f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526d9, value : 32'h8e252084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526da, value : 32'h2045080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526db, value : 32'h70367146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526dc, value : 32'hf006f313},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526dd, value : 32'hf1fd712e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526de, value : 32'hf19a708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526df, value : 32'hb802c107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e0, value : 32'hc10491a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e1, value : 32'h1002254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e2, value : 32'h2005b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e3, value : 32'h90070f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e4, value : 32'h2005c83c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e5, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e6, value : 32'h90c0083c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e7, value : 32'h1040266c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e8, value : 32'hb100b880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526e9, value : 32'h1200b62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ea, value : 32'hc004c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526eb, value : 32'hbea0bda0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ec, value : 32'hc809b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ed, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ee, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ef, value : 32'hb0c0c83c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f0, value : 32'h1600f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f1, value : 32'h80007101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f2, value : 32'h1600018a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f3, value : 32'h80007100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f4, value : 32'h8110006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f5, value : 32'he820044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f6, value : 32'h7014fc8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f7, value : 32'hffc104b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f8, value : 32'h2c00c7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526f9, value : 32'h1404c0ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526fa, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526fb, value : 32'hc809c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526fc, value : 32'h21056832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526fd, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526fe, value : 32'h2105c83c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h526ff, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52700, value : 32'h9120083c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52701, value : 32'hf812104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52702, value : 32'hff780000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52703, value : 32'h1812145},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52704, value : 32'h1600b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52705, value : 32'h80007087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52706, value : 32'hb1e0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52707, value : 32'h710c0320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52708, value : 32'h47cb712d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52709, value : 32'h84900c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5270a, value : 32'hf9574cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5270b, value : 32'h1f000030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5270c, value : 32'h700c1244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5270d, value : 32'h1200b5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5270e, value : 32'h702c742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5270f, value : 32'h901840c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52710, value : 32'hb7200008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52711, value : 32'h2441800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52712, value : 32'h824418fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52713, value : 32'h70441e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52714, value : 32'hc40902c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52715, value : 32'h804418f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52716, value : 32'h9840c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52717, value : 32'hb369680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52718, value : 32'h46280120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52719, value : 32'h47cbd833},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5271a, value : 32'h8009008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5271b, value : 32'h45cbb700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5271c, value : 32'h2889008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5271d, value : 32'ha92d820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5271e, value : 32'hb5c00120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5271f, value : 32'h900743cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52720, value : 32'h1d58c11c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52721, value : 32'h208a9244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52722, value : 32'h1b000010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52723, value : 32'h1b001145},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52724, value : 32'h234f1184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52725, value : 32'h1b0014cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52726, value : 32'h1b001145},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52727, value : 32'h1d001184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52728, value : 32'ha661085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52729, value : 32'h1d580120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5272a, value : 32'h700c9384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5272b, value : 32'hb5c0d920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5272c, value : 32'h1200ae2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5272d, value : 32'h1b0cb7c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5272e, value : 32'hf0659244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5272f, value : 32'h1200a4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52730, value : 32'h46cb740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52731, value : 32'h189018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52732, value : 32'h950016f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52733, value : 32'h2004702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52734, value : 32'hf80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52735, value : 32'h1e00fdff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52736, value : 32'h901b7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52737, value : 32'h40c3c018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52738, value : 32'h4240000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52739, value : 32'hb7204528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5273a, value : 32'h4708b620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5273b, value : 32'h70441e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5273c, value : 32'hc40902c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5273d, value : 32'h90441efc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5273e, value : 32'h90441ef8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5273f, value : 32'h1200a96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52740, value : 32'h10c51e04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52741, value : 32'h78fd720d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52742, value : 32'ha8a702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52743, value : 32'h1e040120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52744, value : 32'h702c1204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52745, value : 32'h9840c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52746, value : 32'ha7a9680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52747, value : 32'hb6a20120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52748, value : 32'h900843cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52749, value : 32'h47c301e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5274a, value : 32'hc11c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5274b, value : 32'h12441b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5274c, value : 32'h1f00d833},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5274d, value : 32'h47cb0145},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5274e, value : 32'h8009008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5274f, value : 32'h1841f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52750, value : 32'h4c7274f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52751, value : 32'h1a8e2355},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52752, value : 32'h1451f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52753, value : 32'h1841f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52754, value : 32'h760cb700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52755, value : 32'h12009b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52756, value : 32'h700cb6a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52757, value : 32'h41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52758, value : 32'h1b002710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52759, value : 32'ha2e1204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5275a, value : 32'h1e000120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5275b, value : 32'h700c1204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5275c, value : 32'h1b00d920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5275d, value : 32'hb6a01344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5275e, value : 32'h1200a1a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5275f, value : 32'h1f0cb7a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52760, value : 32'h9de8244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52761, value : 32'h710c01e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52762, value : 32'h120097e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52763, value : 32'h46cbd878},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52764, value : 32'hc11c900f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52765, value : 32'h14cf2650},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52766, value : 32'h1e00710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52767, value : 32'h1e001185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52768, value : 32'h1f001105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52769, value : 32'h8261185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5276a, value : 32'h1f0000e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5276b, value : 32'hf2a1105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5276c, value : 32'h208afdcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5276d, value : 32'h45cb0d07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5276e, value : 32'h3e09008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5276f, value : 32'h9d6d920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52770, value : 32'h1d000120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52771, value : 32'h700c1045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52772, value : 32'h1eb2b88c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52773, value : 32'hd820101c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52774, value : 32'h101d1f84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52775, value : 32'h1200932},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52776, value : 32'h10051d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52777, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52778, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52779, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5277a, value : 32'h16007a1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5277b, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5277c, value : 32'h7859001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5277d, value : 32'h7fe07839},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5277e, value : 32'h78e0b8c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5277f, value : 32'h2079c2f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52780, value : 32'h43500050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52781, value : 32'h45cb4728},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52782, value : 32'h11e28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52783, value : 32'h3200b8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52784, value : 32'h204e2014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52785, value : 32'h66a8704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52786, value : 32'h20250a2b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52787, value : 32'h20166f14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52788, value : 32'h70420400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52789, value : 32'h60a9e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5278a, value : 32'hcfad880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5278b, value : 32'h41300320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5278c, value : 32'h23912940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5278d, value : 32'h21057146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5278e, value : 32'h90042f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5278f, value : 32'hb1000230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52790, value : 32'h40c3f1eb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52791, value : 32'h4e200000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52792, value : 32'h120094a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52793, value : 32'h66a8702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52794, value : 32'h21d3234f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52795, value : 32'h702ee82b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52796, value : 32'h20166f14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52797, value : 32'h70220400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52798, value : 32'h60a9e024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52799, value : 32'hcbe4062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5279a, value : 32'h42300320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5279b, value : 32'h23942a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5279c, value : 32'h2f812405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5279d, value : 32'h2309004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5279e, value : 32'h8f2b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5279f, value : 32'h740c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a0, value : 32'h2fc7228a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a1, value : 32'h2f802405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a2, value : 32'h2249004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a3, value : 32'h4841800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a4, value : 32'h12008da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a5, value : 32'h2405740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a6, value : 32'h90042f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a7, value : 32'h1800022c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a8, value : 32'h71260484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527a9, value : 32'h9b566a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527aa, value : 32'hd90ca004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ab, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ac, value : 32'h8e21388},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ad, value : 32'h44100120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ae, value : 32'he81a66a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527af, value : 32'h2213234f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b0, value : 32'h6f14704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b1, value : 32'h4002016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b2, value : 32'he0247042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b3, value : 32'h406260a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b4, value : 32'h3200c52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b5, value : 32'h29404130},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b6, value : 32'h71462391},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b7, value : 32'h2f812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b8, value : 32'h2309004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527b9, value : 32'h66a8b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ba, value : 32'ha0040adb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527bb, value : 32'h8a64082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527bc, value : 32'hd90c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527bd, value : 32'he82666a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527be, value : 32'h6f14702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527bf, value : 32'h4002016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c0, value : 32'he0247022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c1, value : 32'h208a60a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c2, value : 32'hc1a0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c3, value : 32'h42300320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c4, value : 32'h23932a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c5, value : 32'h2f812305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c6, value : 32'h2249004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c7, value : 32'h84eb100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c8, value : 32'h740c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527c9, value : 32'h6208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ca, value : 32'h3200bfa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527cb, value : 32'h23054142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527cc, value : 32'h90042f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527cd, value : 32'hb100022c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ce, value : 32'h66a87126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527cf, value : 32'ha00409bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d0, value : 32'h340c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d1, value : 32'h84ed090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d2, value : 32'h702c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d3, value : 32'h3000a86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d4, value : 32'h78e0c6d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d5, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d6, value : 32'h2496b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d7, value : 32'h702c3def},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d8, value : 32'hfcef0bea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527d9, value : 32'h1207c045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527da, value : 32'hc0443091},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527db, value : 32'hc051700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527dc, value : 32'hc04fc050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527dd, value : 32'hc04dc04e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527de, value : 32'hff2f093a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527df, value : 32'h47cbc04c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e0, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e1, value : 32'h40108f61},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e2, value : 32'hb338f20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e3, value : 32'h750c0064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e4, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e5, value : 32'hc8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e6, value : 32'h700cb8e3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e7, value : 32'h2100f208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e8, value : 32'h10200680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527e9, value : 32'h20780080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ea, value : 32'hb8080000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527eb, value : 32'h70422614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ec, value : 32'h48c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ed, value : 32'hb2007124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ee, value : 32'hc205f1e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ef, value : 32'h3ee46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f0, value : 32'hf460001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f1, value : 32'h41c1fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f2, value : 32'hfe2f0822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f3, value : 32'h45cbc005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f4, value : 32'h1268000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f5, value : 32'h264f8d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f6, value : 32'hf2e1401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f7, value : 32'h740cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f8, value : 32'h214a7036},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527f9, value : 32'h8d003480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527fa, value : 32'h33e121ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527fb, value : 32'hf490b8e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527fc, value : 32'h712ec005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527fd, value : 32'h41c3c204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527fe, value : 32'h103f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h527ff, value : 32'h20002900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52800, value : 32'hf0668d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52801, value : 32'h740cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52802, value : 32'h712cc004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52803, value : 32'hfcaf0916},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52804, value : 32'heea704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52805, value : 32'ha8afe0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52806, value : 32'h976fb8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52807, value : 32'h94e0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52808, value : 32'h700c0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52809, value : 32'hfbef0a6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5280a, value : 32'h1600712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5280b, value : 32'h80007082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5280c, value : 32'h22780008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5280d, value : 32'h68210080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5280e, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5280f, value : 32'h510901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52810, value : 32'h2044c047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52811, value : 32'h20002040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52812, value : 32'h1e002003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52813, value : 32'h901c7044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52814, value : 32'ha0f0510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52815, value : 32'h218a00b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52816, value : 32'h218a0048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52817, value : 32'hc0050090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52818, value : 32'h1010260f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52819, value : 32'h2340c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5281a, value : 32'hb802078e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5281b, value : 32'hf822005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5281c, value : 32'h4f8901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5281d, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5281e, value : 32'h4f4901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5281f, value : 32'h714cb220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52820, value : 32'h712cb020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52821, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52822, value : 32'h508901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52823, value : 32'hb887c048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52824, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52825, value : 32'h508901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52826, value : 32'hfcaf088a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52827, value : 32'h83ec004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52828, value : 32'h4210fb8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52829, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5282a, value : 32'hd76ffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5282b, value : 32'h410002e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5282c, value : 32'h208a7056},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5282d, value : 32'hd9ff0fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5282e, value : 32'hb6a711c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5282f, value : 32'h710c02e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52830, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52831, value : 32'hc8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52832, value : 32'hdf080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52833, value : 32'h74441e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52834, value : 32'hc2d49007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52835, value : 32'h1e00d80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52836, value : 32'h901f7085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52837, value : 32'h1e00c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52838, value : 32'h90077085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52839, value : 32'hb02f880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5283a, value : 32'hd90ffcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5283b, value : 32'h2000e5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5283c, value : 32'h9e678cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5283d, value : 32'h212f0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5283e, value : 32'h8d000407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5283f, value : 32'hff081f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52840, value : 32'h141070ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52841, value : 32'h2340301b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52842, value : 32'hf0e83a9b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52843, value : 32'hd80ad93f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52844, value : 32'hfd6f0df6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52845, value : 32'h3f7b914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52846, value : 32'hc0920000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52847, value : 32'h702c42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52848, value : 32'hfaef0fde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52849, value : 32'hc305ba8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5284a, value : 32'h714c740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5284b, value : 32'h3f541c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5284c, value : 32'h1c2c0002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5284d, value : 32'hdd23fc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5284e, value : 32'h1c28fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5284f, value : 32'h8fc03fc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52850, value : 32'h301b1410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52851, value : 32'h3a9b2340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52852, value : 32'h9fdf258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52853, value : 32'h2d008c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52854, value : 32'h12c02e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52855, value : 32'h8f81c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52856, value : 32'h6c02005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52857, value : 32'hc236872},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52858, value : 32'h2e4013a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52859, value : 32'h78651380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5285a, value : 32'hb89cb892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5285b, value : 32'hed86b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5285c, value : 32'h9020c28a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5285d, value : 32'hb2207ad4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5285e, value : 32'h71c5b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5285f, value : 32'hdcef1f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52860, value : 32'hd80f0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52861, value : 32'hfcaf0a62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52862, value : 32'h700cd90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52863, value : 32'hfbef0906},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52864, value : 32'h8f01712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52865, value : 32'h8418fc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52866, value : 32'h78c203a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52867, value : 32'h710443c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52868, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52869, value : 32'h60020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5286a, value : 32'h2c12b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5286b, value : 32'h6038c092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5286c, value : 32'h26f460b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5286d, value : 32'h800070c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5286e, value : 32'h6852048c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5286f, value : 32'h3802b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52870, value : 32'h71647845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52871, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52872, value : 32'h2dc9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52873, value : 32'h20799000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52874, value : 32'ha9000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52875, value : 32'hf1ba71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52876, value : 32'h651dc592},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52877, value : 32'h8f01702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52878, value : 32'h3a408c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52879, value : 32'h41c342c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5287a, value : 32'h103f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5287b, value : 32'hfd6f0d1a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5287c, value : 32'h700e740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5287d, value : 32'h2f8508a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5287e, value : 32'h8000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5287f, value : 32'ha803208b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52880, value : 32'h34401c0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52881, value : 32'h34401c08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52882, value : 32'h2056f411},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52883, value : 32'h28412800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52884, value : 32'h20042182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52885, value : 32'hf80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52886, value : 32'hb826ffc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52887, value : 32'h3f741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52888, value : 32'h68690002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52889, value : 32'hfd6f0ce2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5288a, value : 32'hda08740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5288b, value : 32'h702c40a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5288c, value : 32'h700cc382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5288d, value : 32'h244a633b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5288e, value : 32'h736d7100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5288f, value : 32'h1200210a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52890, value : 32'h31b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52891, value : 32'h20020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52892, value : 32'h148c1101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52893, value : 32'h12cc2c00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52894, value : 32'h78857765},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52895, value : 32'h71247405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52896, value : 32'hb3f228d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52897, value : 32'h140dab00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52898, value : 32'h140b3087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52899, value : 32'h140c3085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5289a, value : 32'h140a3086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5289b, value : 32'hc2223084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5289c, value : 32'h30831409},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5289d, value : 32'h3081140e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5289e, value : 32'h3080140f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5289f, value : 32'h41c3c140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a0, value : 32'h803f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a1, value : 32'hc82c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a2, value : 32'h740cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a3, value : 32'h2040e520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a4, value : 32'hf1b22810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a5, value : 32'h3f941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a6, value : 32'hc6e0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a7, value : 32'h740cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a8, value : 32'hf19f71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528a9, value : 32'h8318f20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528aa, value : 32'h78220064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ab, value : 32'hc8096861},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ac, value : 32'h6c02005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ad, value : 32'h70c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ae, value : 32'h20a86852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528af, value : 32'hc08a0380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b0, value : 32'h4320f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b1, value : 32'h3802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b2, value : 32'h71247845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b3, value : 32'hb89cb892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b4, value : 32'hb060b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b5, value : 32'h2000c76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b6, value : 32'h3fa41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b7, value : 32'hc2a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b8, value : 32'h740cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528b9, value : 32'h42d3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ba, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528bb, value : 32'h202fc046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528bc, value : 32'hc0498648},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528bd, value : 32'h1600f2f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528be, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528bf, value : 32'h817000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c0, value : 32'h700c00fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c1, value : 32'hfbaf0f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c2, value : 32'hd80f712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c3, value : 32'hfcaf08da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c4, value : 32'h700cd90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c5, value : 32'hfbaf0f7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c6, value : 32'h8fc0712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c7, value : 32'h76108f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c8, value : 32'h2d01a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528c9, value : 32'h2440d80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ca, value : 32'h27143c17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528cb, value : 32'h17002397},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528cc, value : 32'h70142100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528cd, value : 32'h2614f4c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ce, value : 32'h80007395},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528cf, value : 32'h2e40048c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d0, value : 32'h24401301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d1, value : 32'h15003e11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d2, value : 32'h21052100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d3, value : 32'h10f98},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d4, value : 32'h200500b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d5, value : 32'h21050600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d6, value : 32'hb80206c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d7, value : 32'h23912114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d8, value : 32'h4802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528d9, value : 32'h2490224f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528da, value : 32'hc8099040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528db, value : 32'h78254350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528dc, value : 32'h20841900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528dd, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528de, value : 32'hc0902010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528df, value : 32'h21141000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e0, value : 32'h3962014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e1, value : 32'h21001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e2, value : 32'hb3fe80e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e3, value : 32'h740c2031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e4, value : 32'h3fb41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e5, value : 32'h42c10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e6, value : 32'hb6e4382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e7, value : 32'h1f00fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e8, value : 32'hf0922045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528e9, value : 32'h20110b23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ea, value : 32'h7014ca07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528eb, value : 32'h20cad812},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ec, value : 32'hc10903e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ed, value : 32'h610813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ee, value : 32'h740cd9ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ef, value : 32'hfd6f0b4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f0, value : 32'h710cb912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f1, value : 32'h2453c046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f2, value : 32'h24ad214d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f3, value : 32'h740c2982},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f4, value : 32'h3fd41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f5, value : 32'h42c10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f6, value : 32'h44a14382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f7, value : 32'hfd6f0b2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f8, value : 32'h4c0250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528f9, value : 32'h20812440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528fa, value : 32'h20056916},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528fb, value : 32'hca070353},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528fc, value : 32'hd8227014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528fd, value : 32'h72120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528fe, value : 32'h4508c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h528ff, value : 32'h8b1c006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52900, value : 32'h16000010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52901, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52902, value : 32'h29090008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52903, value : 32'hf2508014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52904, value : 32'h3fe41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52905, value : 32'haf20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52906, value : 32'h740cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52907, value : 32'hd90fd80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52908, value : 32'hfc6f0fc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52909, value : 32'h23441800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5290a, value : 32'h2000b22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5290b, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5290c, value : 32'h303ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5290d, value : 32'h706c42c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5290e, value : 32'hfd6f0ace},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5290f, value : 32'h160044a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52910, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52911, value : 32'h817000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52912, value : 32'h700c00fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52913, value : 32'hfbaf0e46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52914, value : 32'hd80f712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52915, value : 32'hfc6f0f92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52916, value : 32'h700cd90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52917, value : 32'hfbaf0e36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52918, value : 32'h1500712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52919, value : 32'h20052100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5291a, value : 32'hb8020600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5291b, value : 32'h4802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5291c, value : 32'h19009000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5291d, value : 32'he8122004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5291e, value : 32'h2c40732c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5291f, value : 32'hb99a2184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52920, value : 32'h3442405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52921, value : 32'h42c1740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52922, value : 32'ha7e4382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52923, value : 32'h1800fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52924, value : 32'h1f002104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52925, value : 32'hf0182045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52926, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52927, value : 32'h30401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52928, value : 32'h706c42c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52929, value : 32'hfd6f0a62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5292a, value : 32'h43b144a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5292b, value : 32'h40241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5292c, value : 32'h9360000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5292d, value : 32'h700cfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5292e, value : 32'h24c41800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5292f, value : 32'h21001100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52930, value : 32'h20041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52931, value : 32'hf12c71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52932, value : 32'hfc6f0f1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52933, value : 32'ha7ed90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52934, value : 32'h77270220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52935, value : 32'hc007f10d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52936, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52937, value : 32'h510901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52938, value : 32'h1e00c008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52939, value : 32'h901c7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5293a, value : 32'h9aa0508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5293b, value : 32'hc004fe4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5293c, value : 32'hc32702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5293d, value : 32'h704cfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5293e, value : 32'h40341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5293f, value : 32'ha0a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52940, value : 32'h750cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52941, value : 32'hfdef0ae6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52942, value : 32'h2496c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52943, value : 32'h14043250},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52944, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52945, value : 32'hc1a4c3e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52946, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52947, value : 32'h8ea11228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52948, value : 32'h40d371ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52949, value : 32'h4e7c8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5294a, value : 32'h40027014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5294b, value : 32'h7fb8d912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5294c, value : 32'hd92f209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5294d, value : 32'h40020280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5294e, value : 32'hcced912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5294f, value : 32'hda800060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52950, value : 32'hf0ef003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52951, value : 32'hbf20200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52952, value : 32'hc08002e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52953, value : 32'hc46c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52954, value : 32'hd912fdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52955, value : 32'h259f8e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52956, value : 32'h209f12c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52957, value : 32'h704c0582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52958, value : 32'h708cc380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52959, value : 32'h6f12651d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5295a, value : 32'h250078e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5295b, value : 32'hf6a1401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5295c, value : 32'h780f0460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5295d, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5295e, value : 32'ha1a4e20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5295f, value : 32'h702c00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52960, value : 32'h78e0c7c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52961, value : 32'h2482c3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52962, value : 32'h44103104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52963, value : 32'h702cc081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52964, value : 32'hfaef0b6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52965, value : 32'h4228a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52966, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52967, value : 32'h8d401228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52968, value : 32'h20502479},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52969, value : 32'h22102040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5296a, value : 32'ha0432442},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5296b, value : 32'h41c3750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5296c, value : 32'h30151},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5296d, value : 32'hfd6f0952},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5296e, value : 32'h400240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5296f, value : 32'h24408da0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52970, value : 32'hc8093081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52971, value : 32'h7d05bd0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52972, value : 32'hfcaf0d06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52973, value : 32'h46084082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52974, value : 32'h1f802505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52975, value : 32'hd90003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52976, value : 32'hb56d940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52977, value : 32'h43100460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52978, value : 32'h2200916},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52979, value : 32'h1402be68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5297a, value : 32'h7fd03102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5297b, value : 32'h41e14082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5297c, value : 32'h80a41f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5297d, value : 32'h4250fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5297e, value : 32'h41c3e807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5297f, value : 32'h155},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52980, value : 32'hfaef0fe6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52981, value : 32'h2840700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52982, value : 32'h70cd2200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52983, value : 32'h47cb7d05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52984, value : 32'h4848000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52985, value : 32'h1f952505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52986, value : 32'hd80003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52987, value : 32'h258c7dd0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52988, value : 32'hf7139fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52989, value : 32'hb0a40a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5298a, value : 32'h41a10460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5298b, value : 32'h20008ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5298c, value : 32'h41224082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5298d, value : 32'hfb2f0fc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5298e, value : 32'hc1814242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5298f, value : 32'ha90061b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52990, value : 32'h661e8f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52991, value : 32'h40a2f1ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52992, value : 32'h4600ae6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52993, value : 32'h2b40702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52994, value : 32'h70ad2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52995, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52996, value : 32'h220089e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52997, value : 32'hd92bb0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52998, value : 32'h8a6740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52999, value : 32'hb913fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5299a, value : 32'h21c22042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5299b, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5299c, value : 32'h20159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5299d, value : 32'hfd6f0892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5299e, value : 32'h8f804302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5299f, value : 32'h7200244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a0, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a1, value : 32'h30020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a2, value : 32'h659ec081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a3, value : 32'h224e60a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a4, value : 32'h714401c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a5, value : 32'h290045c9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a6, value : 32'h7b050000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a7, value : 32'h41c37a6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a8, value : 32'h1015a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529a9, value : 32'hfd6f0862},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529aa, value : 32'h268c740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ab, value : 32'h45c99004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ac, value : 32'h41c3f6a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ad, value : 32'h15b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ae, value : 32'hfd6f084e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529af, value : 32'h8f40740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b0, value : 32'h208c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b1, value : 32'hf7088fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b2, value : 32'h6109c181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b3, value : 32'h20c07034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b4, value : 32'hf3f90081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b5, value : 32'h3f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b6, value : 32'h268c7e0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b7, value : 32'hf6889004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b8, value : 32'h700cd957},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529b9, value : 32'hfaef0f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ba, value : 32'hf009b912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529bb, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529bc, value : 32'h1015d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529bd, value : 32'hfd6f0812},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529be, value : 32'h40c342c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529bf, value : 32'h1258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c0, value : 32'h6d2988a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c1, value : 32'h114090b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c2, value : 32'h180074ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c3, value : 32'h47cb0103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c4, value : 32'h1015e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c5, value : 32'h41e1740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c6, value : 32'hfd2f0fee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c7, value : 32'hbd0542a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c8, value : 32'h1401274f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529c9, value : 32'hfe2740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ca, value : 32'h42a1fd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529cb, value : 32'h780e4eb0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529cc, value : 32'h78e0c7d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529cd, value : 32'hc1a4c3e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ce, value : 32'h800145cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529cf, value : 32'h40a14e7c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d0, value : 32'h2a00b82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d1, value : 32'h40a1d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d2, value : 32'habed910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d3, value : 32'hda410060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d4, value : 32'hd91040a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d5, value : 32'hfbef0bc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d6, value : 32'h40a1daf3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d7, value : 32'h2a00b66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d8, value : 32'h40a1d929},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529d9, value : 32'hbb6d929},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529da, value : 32'hda1ffbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529db, value : 32'h2e009ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529dc, value : 32'hc080c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529dd, value : 32'hfdef0a1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529de, value : 32'hc080d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529df, value : 32'hfdef0a16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e0, value : 32'h40a1d929},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e1, value : 32'hc280702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e2, value : 32'ha52dbff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e3, value : 32'h708c04a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e4, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e5, value : 32'hffe4e20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e6, value : 32'h702c00a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e7, value : 32'hcb240a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e8, value : 32'hd9290220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529e9, value : 32'h78e0c7c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ea, value : 32'hc1a2c3ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529eb, value : 32'h800145cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ec, value : 32'h41304d6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ed, value : 32'hd8644010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ee, value : 32'h254070cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ef, value : 32'hb5001312},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f0, value : 32'hc640c641},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f1, value : 32'h731478cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f2, value : 32'hd00f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f3, value : 32'h20100919},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f4, value : 32'hd00829},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f5, value : 32'h50081f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f6, value : 32'h900829},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f7, value : 32'hd87fe896},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f8, value : 32'hf01eb808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529f9, value : 32'hd0082d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529fa, value : 32'h500831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529fb, value : 32'h90080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529fc, value : 32'hd87fe898},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529fd, value : 32'hf014b810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529fe, value : 32'h7f0040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h529ff, value : 32'hf0107f7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a00, value : 32'h7f7f40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a01, value : 32'hf00c007f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a02, value : 32'h700cd987},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a03, value : 32'hf00eb911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a04, value : 32'h7f40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a05, value : 32'hf0047f7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a06, value : 32'hb818d87f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a07, value : 32'hf008c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a08, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a09, value : 32'h115},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a0a, value : 32'hfacf0dbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a0b, value : 32'h15001502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a0c, value : 32'hd52b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a0d, value : 32'h7810fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a0e, value : 32'hd907d841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a0f, value : 32'hda08b813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a10, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a11, value : 32'ha9e70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a12, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a13, value : 32'h742c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a14, value : 32'hfbaf0d86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a15, value : 32'hc080714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a16, value : 32'hcde4102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a17, value : 32'h724cfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a18, value : 32'hd914700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a19, value : 32'hfbaf0d72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a1a, value : 32'h706c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a1b, value : 32'h4060d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a1c, value : 32'hb892744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a1d, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a1e, value : 32'hfbaf0a6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a1f, value : 32'h160070cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a20, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a21, value : 32'h811000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a22, value : 32'h700c003e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a23, value : 32'hd4ad914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a24, value : 32'h714cfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a25, value : 32'hd907d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a26, value : 32'hda08b893},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a27, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a28, value : 32'ha4270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a29, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a2a, value : 32'hfb4f09de},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a2b, value : 32'h7704b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a2c, value : 32'h20141a02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a2d, value : 32'hf18871c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a2e, value : 32'h78e0c7cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a2f, value : 32'h4608c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a30, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a31, value : 32'hc8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a32, value : 32'h47284050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a33, value : 32'h8e00204b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a34, value : 32'h40c3f2b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a35, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a36, value : 32'h20812078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a37, value : 32'h219f8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a38, value : 32'h209f02c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a39, value : 32'h61190582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a3a, value : 32'hf8f2132},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a3b, value : 32'h4e8e8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a3c, value : 32'hfb4f09ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a3d, value : 32'hd907706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a3e, value : 32'h744c4568},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a3f, value : 32'h708cbd9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a40, value : 32'h70ac40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a41, value : 32'hfbaf09de},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a42, value : 32'h43e170cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a43, value : 32'h238540a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a44, value : 32'h762c0201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a45, value : 32'h244a744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a46, value : 32'h250a0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a47, value : 32'h9c60400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a48, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a49, value : 32'hd90740a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a4a, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a4b, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a4c, value : 32'hfbaf09b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a4d, value : 32'hfc1268a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a4e, value : 32'hfb8f0c56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a4f, value : 32'h13c0254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a50, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a51, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a52, value : 32'h99a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a53, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a54, value : 32'hd90740a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a55, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a56, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a57, value : 32'hfbaf0986},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a58, value : 32'h3c0264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a59, value : 32'hd9077ebd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a5a, value : 32'h744c40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a5b, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a5c, value : 32'h97270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a5d, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a5e, value : 32'hd90740a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a5f, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a60, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a61, value : 32'hfbaf095e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a62, value : 32'hfc3268a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a63, value : 32'hd90740c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a64, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a65, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a66, value : 32'hfbaf094a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a67, value : 32'h40a170cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a68, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a69, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a6a, value : 32'h93a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a6b, value : 32'h268afbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a6c, value : 32'h40c10fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a6d, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a6e, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a6f, value : 32'h92670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a70, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a71, value : 32'hd90740a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a72, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a73, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a74, value : 32'hfbaf0912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a75, value : 32'hfc3268a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a76, value : 32'h1480254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a77, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a78, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a79, value : 32'h8fe70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a7a, value : 32'h71ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a7b, value : 32'hfb8f0b8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a7c, value : 32'hd90740a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a7d, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a7e, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a7f, value : 32'hfbaf08e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a80, value : 32'h40a173cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a81, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a82, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a83, value : 32'h8d670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a84, value : 32'h268afbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a85, value : 32'h40a10fc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a86, value : 32'h744c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a87, value : 32'h244a43e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a88, value : 32'h250a0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a89, value : 32'h8be0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a8a, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a8b, value : 32'hd90740a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a8c, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a8d, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a8e, value : 32'hfc0264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a8f, value : 32'h862f03f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a90, value : 32'h700cfb4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a91, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a92, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a93, value : 32'h89670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a94, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a95, value : 32'hfb8f0b3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a96, value : 32'hd907706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a97, value : 32'h724c4568},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a98, value : 32'h708cbd99},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a99, value : 32'h70ac40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a9a, value : 32'hfbaf087a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a9b, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a9c, value : 32'h42c1d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a9d, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a9e, value : 32'h86a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52a9f, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa0, value : 32'hbd2d740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa1, value : 32'h712cb892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa2, value : 32'h43a142e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa3, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa4, value : 32'hfbaf0852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa5, value : 32'h6d1370cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa6, value : 32'hda0cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa7, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa8, value : 32'h84270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aa9, value : 32'h71ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aaa, value : 32'hfb8f0ace},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aab, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aac, value : 32'h706cda10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aad, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aae, value : 32'h82a70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aaf, value : 32'hd880fb8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab0, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab1, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab2, value : 32'h81a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab3, value : 32'h70ccfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab4, value : 32'h78e0c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab5, value : 32'h4510c2f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab6, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab7, value : 32'h508901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab8, value : 32'h20534330},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ab9, value : 32'hf4098196},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aba, value : 32'h3e241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52abb, value : 32'hc1a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52abc, value : 32'h740cfd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52abd, value : 32'h265f71ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52abe, value : 32'h2e4020cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52abf, value : 32'h710c2094},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac0, value : 32'h200e241f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac1, value : 32'h93a50ffd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac2, value : 32'hf967104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac3, value : 32'h740cfb0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac4, value : 32'h3e341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac5, value : 32'hbf20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac6, value : 32'h42c2fd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac7, value : 32'hfb8f0a72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac8, value : 32'h2280265f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ac9, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aca, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52acb, value : 32'h770470ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52acc, value : 32'h2007212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52acd, value : 32'hfae700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ace, value : 32'h260afb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52acf, value : 32'h6f010440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad0, value : 32'h7b0f702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad1, value : 32'h986d807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad2, value : 32'h704c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad3, value : 32'h45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad4, value : 32'h232f12c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad5, value : 32'hd81d0580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad6, value : 32'h426241a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad7, value : 32'h20096e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad8, value : 32'hd81e4270},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ad9, value : 32'h426241a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ada, value : 32'h200962},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52adb, value : 32'hd81f4342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52adc, value : 32'h426241a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52add, value : 32'h200956},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ade, value : 32'hd8204342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52adf, value : 32'h704c41a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae0, value : 32'h20094a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae1, value : 32'h78f24342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae2, value : 32'h661e702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae3, value : 32'h7bcfd807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae4, value : 32'h93a704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae5, value : 32'h40700020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae6, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae7, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae8, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ae9, value : 32'hfb6f0f3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aea, value : 32'h440260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aeb, value : 32'h20402242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aec, value : 32'h262fd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aed, value : 32'h700c0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aee, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aef, value : 32'hf26708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af0, value : 32'h70acfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af1, value : 32'h710cdd08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af2, value : 32'hb7a41c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af3, value : 32'h4262fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af4, value : 32'h41c2700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af5, value : 32'hfbaf0b6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af6, value : 32'h258c4262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af7, value : 32'h700c1dff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af8, value : 32'hda5cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52af9, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52afa, value : 32'h70cc70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52afb, value : 32'hfb6f0ef6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52afc, value : 32'h708c71ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52afd, value : 32'h458874cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52afe, value : 32'hbd8cbe92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52aff, value : 32'hd92e40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b00, value : 32'h43a142a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b01, value : 32'hede70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b02, value : 32'h70ccfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b03, value : 32'hd92f40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b04, value : 32'h43a142a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b05, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b06, value : 32'hfb6f0eca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b07, value : 32'h6d1370cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b08, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b09, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b0a, value : 32'heba70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b0b, value : 32'h71ccfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b0c, value : 32'h540202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b0d, value : 32'hc8d2054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b0e, value : 32'h2580241f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b0f, value : 32'h8fd46ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b10, value : 32'h71c68364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b11, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b12, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b13, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b14, value : 32'hfb6f0e92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b15, value : 32'h440260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b16, value : 32'h1500261e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b17, value : 32'h704c702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b18, value : 32'h671f78a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b19, value : 32'h7b0f6f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b1a, value : 32'h200862},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b1b, value : 32'hdd25d807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b1c, value : 32'hbd07d81d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b1d, value : 32'h41a14262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b1e, value : 32'h200852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b1f, value : 32'hd81e4342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b20, value : 32'h426241a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b21, value : 32'h200846},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b22, value : 32'hd81f4342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b23, value : 32'h426241a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b24, value : 32'h20083a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b25, value : 32'hd8204342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b26, value : 32'h704c41a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b27, value : 32'h20082e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b28, value : 32'hd8074342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b29, value : 32'h704c702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b2a, value : 32'h200822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b2b, value : 32'h700c4302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b2c, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b2d, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b2e, value : 32'he2a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b2f, value : 32'h260afb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b30, value : 32'h8b60440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b31, value : 32'hc6d4fb8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b32, value : 32'h4648c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b33, value : 32'h40104728},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b34, value : 32'h6b09eb0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b35, value : 32'h68a1780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b36, value : 32'h4102700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b37, value : 32'h43e1704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b38, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b39, value : 32'hfb6f0dfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b3a, value : 32'h258c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b3b, value : 32'hc6c81e3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b3c, value : 32'h4050c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b3d, value : 32'h47cb4528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b3e, value : 32'h4988000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b3f, value : 32'h8703e81b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b40, value : 32'he8877104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b41, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b42, value : 32'h25c9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b43, value : 32'h720ca703},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b44, value : 32'h900746cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b45, value : 32'ha56c25c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b46, value : 32'h1e0000a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b47, value : 32'h16001005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b48, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b49, value : 32'h2053000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b4a, value : 32'hf223817e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b4b, value : 32'h90051ecc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b4c, value : 32'hc809f021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b4d, value : 32'h46cb70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b4e, value : 32'hc3ec9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b4f, value : 32'h21056832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b50, value : 32'h903b0f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b51, value : 32'hb0a0c02c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b52, value : 32'h268079c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b53, value : 32'hd8141939},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b54, value : 32'h9b6b1a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b55, value : 32'hb6a000a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b56, value : 32'h90451e2c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b57, value : 32'h93441ed8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b58, value : 32'h93441ed4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b59, value : 32'hb6068703},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b5a, value : 32'h93441ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b5b, value : 32'h1eccc6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b5c, value : 32'h740c9344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b5d, value : 32'h900746cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b5e, value : 32'h9f2c224},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b5f, value : 32'hb6a000a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b60, value : 32'h10051e08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b61, value : 32'h20300819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b62, value : 32'h90051e58},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b63, value : 32'h20710823},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b64, value : 32'h1e00700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b65, value : 32'h90077285},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b66, value : 32'hf010c254},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b67, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b68, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b69, value : 32'hc3ec9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b6a, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b6b, value : 32'h41c3f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b6c, value : 32'h34a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b6d, value : 32'hfacf0832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b6e, value : 32'h74041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b6f, value : 32'hc2509007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b70, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b71, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b72, value : 32'hc02c903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b73, value : 32'h851800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b74, value : 32'h78e0c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b75, value : 32'hc1a2c3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b76, value : 32'hb99fd925},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b77, value : 32'h1c068900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b78, value : 32'h891b3002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b79, value : 32'h30021c07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b7a, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b7b, value : 32'h8820122c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b7c, value : 32'h8822c161},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b7d, value : 32'h30421c05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b7e, value : 32'h88038821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b7f, value : 32'h30421c02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b80, value : 32'hfeaf0a4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b81, value : 32'h30021c03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b82, value : 32'h70ed4110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b83, value : 32'h218121ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b84, value : 32'hfa9714e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b85, value : 32'h2a001465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b86, value : 32'h70cd23d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b87, value : 32'he99c806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b88, value : 32'h24401005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b89, value : 32'h60c83180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b8a, value : 32'ha000250b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b8b, value : 32'h2714f242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b8c, value : 32'h700e1380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b8d, value : 32'h20142a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b8e, value : 32'h30802440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b8f, value : 32'h3932032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b90, value : 32'h60cdc081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b91, value : 32'hb6d78af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b92, value : 32'h78cf2024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b93, value : 32'hff6f0f9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b94, value : 32'h6e3479ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b95, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b96, value : 32'he81311e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b97, value : 32'h20402040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b98, value : 32'h3c32116},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b99, value : 32'h6d817910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b9a, value : 32'h61596179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b9b, value : 32'h3021920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b9c, value : 32'h408212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b9d, value : 32'h61596179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b9e, value : 32'h3421920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52b9f, value : 32'h232ff016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba0, value : 32'h79f60408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba1, value : 32'h16006179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba2, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba3, value : 32'h240b0121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba4, value : 32'h6d01a000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba5, value : 32'hf2066159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba6, value : 32'h21920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba7, value : 32'hf005a9a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba8, value : 32'h1920a900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ba9, value : 32'h40020342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52baa, value : 32'h204072a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bab, value : 32'hf1cc0050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bac, value : 32'hf1b671c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bad, value : 32'hf1af71e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bae, value : 32'h78e0c7d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52baf, value : 32'hdb24c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb0, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb1, value : 32'hbb9f122c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb2, value : 32'h31a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb3, value : 32'he0078b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb4, value : 32'hc12841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb5, value : 32'h69898b1c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb6, value : 32'he80faa81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb7, value : 32'h791dc805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb8, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bb9, value : 32'h3f8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bba, value : 32'hb9c6e007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bbb, value : 32'haa22b823},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bbc, value : 32'h68c96038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bbd, value : 32'h4689f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bbe, value : 32'h12b5aa22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bbf, value : 32'h788f008d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc0, value : 32'haac37104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc1, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc2, value : 32'h20a8770c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc3, value : 32'h71040180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc4, value : 32'h100d250f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc5, value : 32'h42c378cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc6, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc7, value : 32'h64081b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc8, value : 32'h7822aaa0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bc9, value : 32'h240a7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bca, value : 32'h20a87000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bcb, value : 32'h250f0180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bcc, value : 32'h7124104d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bcd, value : 32'h70adaaa0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bce, value : 32'h800044cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bcf, value : 32'hd4311e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd0, value : 32'h408910b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd1, value : 32'h706d70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd2, value : 32'hb3179af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd3, value : 32'h70751095},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd4, value : 32'h20ca4060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd5, value : 32'h80000f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd6, value : 32'h88e0003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd7, value : 32'hff6f0e8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd8, value : 32'he80578cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bd9, value : 32'hb8236f07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bda, value : 32'h4f1ff003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bdb, value : 32'h1802b824},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bdc, value : 32'h71c51012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bdd, value : 32'hf1eb7165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bde, value : 32'h71a57185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bdf, value : 32'hc6c6f1e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be0, value : 32'h8bac0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be1, value : 32'hc0d10100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be2, value : 32'h700c7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be3, value : 32'he9058840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be4, value : 32'h1f0a0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be5, value : 32'hbae07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be6, value : 32'h88217de0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be7, value : 32'hf78ae1c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be8, value : 32'h20e07354},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52be9, value : 32'h218007cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bea, value : 32'ha821003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52beb, value : 32'hf0086a21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bec, value : 32'h7ce07054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bed, value : 32'h8012154},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bee, value : 32'h6a29a821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bef, value : 32'ha8207fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf0, value : 32'h443216f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf1, value : 32'h11fe8940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf2, value : 32'h229f8101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf3, value : 32'h790c041f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf4, value : 32'h802905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf5, value : 32'h71047fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf6, value : 32'h2482c3f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf7, value : 32'h16003302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf8, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bf9, value : 32'hb8c30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bfa, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bfb, value : 32'h205f1228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bfc, value : 32'h752c0b16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bfd, value : 32'h702eb916},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bfe, value : 32'h15802700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52bff, value : 32'h11808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c00, value : 32'hfcef0f06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c01, value : 32'hf32d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c02, value : 32'h42d3ff8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c03, value : 32'h11408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c04, value : 32'h448202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c05, value : 32'h31812440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c06, value : 32'h31422440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c07, value : 32'hfeaf09f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c08, value : 32'h31c32440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c09, value : 32'hf4e37014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c0a, value : 32'h30801407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c0b, value : 32'hfdaf085a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c0c, value : 32'h20431a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c0d, value : 32'h30801405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c0e, value : 32'ha4e712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c0f, value : 32'h4310fdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c10, value : 32'h406270ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c11, value : 32'h704c712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c12, value : 32'hffaf0f62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c13, value : 32'h23421a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c14, value : 32'h30801406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c15, value : 32'h724cc182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c16, value : 32'h708c716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c17, value : 32'hfaaf0eb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c18, value : 32'hc0834010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c19, value : 32'h89a702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c1a, value : 32'hda80faaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c1b, value : 32'h2002258a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c1c, value : 32'h70cd708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c1d, value : 32'h222f8f20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c1e, value : 32'h40620507},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c1f, value : 32'hff6f0d82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c20, value : 32'h4002c540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c21, value : 32'h724cc180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c22, value : 32'he86716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c23, value : 32'h708cfaaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c24, value : 32'h30801401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c25, value : 32'h81be2053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c26, value : 32'hc083f205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c27, value : 32'h180060d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c28, value : 32'h71860043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c29, value : 32'h2a3f258d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c2a, value : 32'h8f6071c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c2b, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c2c, value : 32'h20142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c2d, value : 32'hfcef0e52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c2e, value : 32'h70ad4202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c2f, value : 32'hc083de80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c30, value : 32'h14341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c31, value : 32'h60aa0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c32, value : 32'hfcef0e3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c33, value : 32'h268d740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c34, value : 32'h71a51e7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c35, value : 32'h740cd951},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c36, value : 32'hfcef0e2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c37, value : 32'h248ab912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c38, value : 32'h77ad7002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c39, value : 32'h776d700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c3a, value : 32'h20a8776c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c3b, value : 32'hc1830740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c3c, value : 32'h610977b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c3d, value : 32'he0fff207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c3e, value : 32'he914f202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c3f, value : 32'h6829e906},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c40, value : 32'he98ff005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c41, value : 32'hf00e4508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c42, value : 32'h2302d97f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c43, value : 32'h49b210cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c44, value : 32'h25ca7291},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c45, value : 32'h21ca10cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c46, value : 32'h43a102cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c47, value : 32'h77ad4328},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c48, value : 32'h77747104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c49, value : 32'h77b5f404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c4a, value : 32'hf404de7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c4b, value : 32'h46694568},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c4c, value : 32'h41a18f60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c4d, value : 32'h21b94eb0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c4e, value : 32'h207f0fff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c4f, value : 32'h78240100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c50, value : 32'h14641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c51, value : 32'hca20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c52, value : 32'h4202faaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c53, value : 32'h41c366b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c54, value : 32'h30147},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c55, value : 32'h942844},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c56, value : 32'h42a1740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c57, value : 32'hdaa43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c58, value : 32'h240afcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c59, value : 32'h8f200500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c5a, value : 32'h843e2105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c5b, value : 32'h26144620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c5c, value : 32'h70022040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c5d, value : 32'h180860f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c5e, value : 32'hf20b0502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c5f, value : 32'h2011081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c60, value : 32'h510e19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c61, value : 32'h75021e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c62, value : 32'h4e8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c63, value : 32'h1e00f013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c64, value : 32'h80007502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c65, value : 32'hf00f0033},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c66, value : 32'h20510813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c67, value : 32'h110e0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c68, value : 32'h75021e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c69, value : 32'h348000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c6a, value : 32'h1e00f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c6b, value : 32'h80007502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c6c, value : 32'h242f004f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c6d, value : 32'h250a0507},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c6e, value : 32'h245f0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c6f, value : 32'h20540140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c70, value : 32'h78300c81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c71, value : 32'h2822845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c72, value : 32'h209e4040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c73, value : 32'h60380dbf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c74, value : 32'h14841c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c75, value : 32'h7b100005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c76, value : 32'hfcef0d2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c77, value : 32'h4062750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c78, value : 32'hb36702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c79, value : 32'h1a00fdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c7a, value : 32'h71262043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c7b, value : 32'h448202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c7c, value : 32'h6207414},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c7d, value : 32'h40c3ffc5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c7e, value : 32'h12e08000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c7f, value : 32'h431800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c80, value : 32'h78e0c7d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c81, value : 32'h88606038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c82, value : 32'ha8607b45},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c83, value : 32'h83104b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c84, value : 32'h184b7b45},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c85, value : 32'h109600c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c86, value : 32'h7b450083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c87, value : 32'hc21896},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c88, value : 32'h8310e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c89, value : 32'h7fe07a65},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c8a, value : 32'h8218e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c8b, value : 32'h2482c3ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c8c, value : 32'h266f3206},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c8d, value : 32'hc0801243},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c8e, value : 32'hff2f08da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c8f, value : 32'h10901600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c90, value : 32'h800140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c91, value : 32'h88404e7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c92, value : 32'h7a058813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c93, value : 32'h30811403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c94, value : 32'h30801416},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c95, value : 32'h78477825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c96, value : 32'h1be080b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c97, value : 32'h99e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c98, value : 32'h256f03c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c99, value : 32'h150016c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c9a, value : 32'h81110c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c9b, value : 32'hc0800032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c9c, value : 32'h8aad913},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c9d, value : 32'hdaf3fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c9e, value : 32'h3bc02456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52c9f, value : 32'hfd6f0dfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca0, value : 32'h20d02053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca1, value : 32'h3bc02456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca2, value : 32'h2600eba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca3, value : 32'hc080d90b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca4, value : 32'hda45d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca5, value : 32'hffef0f72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca6, value : 32'h30112440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca7, value : 32'h3bc02456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca8, value : 32'h2600ea2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ca9, value : 32'h2456d946},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52caa, value : 32'he9a3bc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cab, value : 32'hd9470260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cac, value : 32'h3bc02456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cad, value : 32'h2600e8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cae, value : 32'h2456d948},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52caf, value : 32'he863bc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb0, value : 32'hd9490260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb1, value : 32'h3bc02456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb2, value : 32'h2600e7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb3, value : 32'hca0ed94a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb4, value : 32'h47cb704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb5, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb6, value : 32'h50a31},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb7, value : 32'h2b01205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb8, value : 32'hf832232},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cb9, value : 32'h4788000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cba, value : 32'h79557322},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cbb, value : 32'h673f7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cbc, value : 32'hab208f28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cbd, value : 32'h1b968f2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cbe, value : 32'h8f290042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cbf, value : 32'h421b4b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc0, value : 32'h1be18f2b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc1, value : 32'hf1e70042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc2, value : 32'h3bc22456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc3, value : 32'h712cc080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc4, value : 32'hecadbff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc5, value : 32'h708c0420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc6, value : 32'hd910c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc7, value : 32'hfb6f0ffe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc8, value : 32'h8d00dabc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cc9, value : 32'h5e0815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cca, value : 32'h8118e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ccb, value : 32'hc080017f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ccc, value : 32'hed6d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ccd, value : 32'hda40ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cce, value : 32'h2600dfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ccf, value : 32'h3bc02456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd0, value : 32'h3bc02456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd1, value : 32'hfd6f0e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd2, value : 32'hc027d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd3, value : 32'h17f0819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd4, value : 32'hd91cc080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd5, value : 32'hffef0eb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd6, value : 32'h2456724c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd7, value : 32'he363bc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd8, value : 32'hd91cfd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cd9, value : 32'h3bc22456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cda, value : 32'h702cc080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cdb, value : 32'he6edbff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cdc, value : 32'h708c0420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cdd, value : 32'h80f8d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cde, value : 32'h8e00005e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cdf, value : 32'hba8b8e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce0, value : 32'hb76fec1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce1, value : 32'hf1afccf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce2, value : 32'h8d00facf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce3, value : 32'hf29eb8e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce4, value : 32'hb8e58e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce5, value : 32'hb66f49a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce6, value : 32'hdf6fd8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce7, value : 32'hd8100240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce8, value : 32'hb16d940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ce9, value : 32'hda0ffb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cea, value : 32'h762c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ceb, value : 32'hfb6f0a2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cec, value : 32'h8f20714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ced, value : 32'h582219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cee, value : 32'h100017bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cef, value : 32'h88216038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf0, value : 32'hdf090d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf1, value : 32'h20538814},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf2, value : 32'hf23580fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf3, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf4, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf5, value : 32'hd2a012c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf6, value : 32'hda4bfa6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf7, value : 32'h3a002456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf8, value : 32'h2600d8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cf9, value : 32'h831800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cfa, value : 32'heaa700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cfb, value : 32'h712cfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cfc, value : 32'hfacf0eae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cfd, value : 32'h2400d9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cfe, value : 32'h752c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52cff, value : 32'hfb6f09da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d00, value : 32'h40c3714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d01, value : 32'h3a980000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d02, value : 32'h600b8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d03, value : 32'hae2742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d04, value : 32'h710c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d05, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d06, value : 32'h12c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d07, value : 32'h2400ec2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d08, value : 32'h340c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d09, value : 32'hb6e0d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d0a, value : 32'hd9080060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d0b, value : 32'h1200b32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d0c, value : 32'hd810710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d0d, value : 32'ha82702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d0e, value : 32'hda0ffb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d0f, value : 32'h762c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d10, value : 32'hfb6f0996},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d11, value : 32'h700c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d12, value : 32'h704cd932},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d13, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d14, value : 32'he9273ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d15, value : 32'h70ccfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d16, value : 32'hd933700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d17, value : 32'h706cda20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d18, value : 32'h73ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d19, value : 32'hfb2f0e7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d1a, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d1b, value : 32'h96a762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d1c, value : 32'h714cfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d1d, value : 32'hd938d811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d1e, value : 32'hfb6f0a3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d1f, value : 32'h700cda0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d20, value : 32'h956d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d21, value : 32'h714cfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d22, value : 32'hd930700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d23, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d24, value : 32'h73ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d25, value : 32'hfb2f0e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d26, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d27, value : 32'h704cd931},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d28, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d29, value : 32'he3e73ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d2a, value : 32'h70ccfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d2b, value : 32'h762c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d2c, value : 32'hfb6f0926},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d2d, value : 32'hcb6714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d2e, value : 32'h700c0240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d2f, value : 32'hfb2f0dd6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d30, value : 32'h9d2712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d31, value : 32'hf027fdcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d32, value : 32'hda20d825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d33, value : 32'h706cb89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d34, value : 32'h70cc708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d35, value : 32'h881b8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d36, value : 32'hd90b7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d37, value : 32'h452053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d38, value : 32'hfb2f0e02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d39, value : 32'h700c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d3a, value : 32'h724cd928},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d3b, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d3c, value : 32'hdf273ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d3d, value : 32'h70ccfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d3e, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d3f, value : 32'h706cda1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d40, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d41, value : 32'hfb2f0dde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d42, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d43, value : 32'hfb2f0d86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d44, value : 32'h702c712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d45, value : 32'h70441e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d46, value : 32'hc200901f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d47, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d48, value : 32'h968000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d49, value : 32'h11e0815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d4a, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d4b, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d4c, value : 32'hc0049007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d4d, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d4e, value : 32'h900840c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d4f, value : 32'hb02001b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d50, value : 32'h1cc3266f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d51, value : 32'h8e00b036},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d52, value : 32'hf01ae89e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d53, value : 32'h1600e908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d54, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d55, value : 32'he88b0040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d56, value : 32'hf011710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d57, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d58, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d59, value : 32'h700c7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d5a, value : 32'h710cf209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d5b, value : 32'hb1a7838},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d5c, value : 32'h780ffd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d5d, value : 32'hfb8f0c7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d5e, value : 32'h68218f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d5f, value : 32'h792faf20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d60, value : 32'h809409cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d61, value : 32'hfd6f0b02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d62, value : 32'h70ad730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d63, value : 32'h8e20b7a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d64, value : 32'h9f6e984},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d65, value : 32'h8e200240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d66, value : 32'h900740c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d67, value : 32'hb0a0c2cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d68, value : 32'he989b0a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d69, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d6a, value : 32'h108000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d6b, value : 32'hf647114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d6c, value : 32'h8320202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d6d, value : 32'had6ff4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d6e, value : 32'hc7cafd8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d6f, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d70, value : 32'h7fe0700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d71, value : 32'hc420ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d72, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d73, value : 32'hc1a2b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d74, value : 32'hc8094608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d75, value : 32'h6d41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d76, value : 32'hb8020002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d77, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d78, value : 32'h200c900c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d79, value : 32'h78bd90a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d7a, value : 32'h70901600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d7b, value : 32'h48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d7c, value : 32'h4f2044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d7d, value : 32'h10432544},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d7e, value : 32'h42e1d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d7f, value : 32'hfcef090a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d80, value : 32'h20534078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d81, value : 32'hc04020c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d82, value : 32'hc200ef8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d83, value : 32'h6e41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d84, value : 32'h8f60001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d85, value : 32'hd80afcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d86, value : 32'h3e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d87, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d88, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d89, value : 32'h140c9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d8a, value : 32'h30310821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d8b, value : 32'h1131000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d8c, value : 32'h10c02d41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d8d, value : 32'h1ac125ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d8e, value : 32'hf832084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d8f, value : 32'h60b8742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d90, value : 32'h380205a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d91, value : 32'hf004e038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d92, value : 32'h732cd870},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d93, value : 32'h6038710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d94, value : 32'h1e007017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d95, value : 32'h90037404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d96, value : 32'h1e00d878},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d97, value : 32'h90077404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d98, value : 32'h2f4f87c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d99, value : 32'hc0410022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d9a, value : 32'h2ec70d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d9b, value : 32'h710c0021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d9c, value : 32'h100087e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d9d, value : 32'h45cbc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d9e, value : 32'hc400900f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52d9f, value : 32'h14ce2550},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da0, value : 32'hb802726d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da1, value : 32'h3412005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da2, value : 32'h190078c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da3, value : 32'h180002c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da4, value : 32'h8da02c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da5, value : 32'hd81e0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da6, value : 32'h36091209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da7, value : 32'h702e700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da8, value : 32'h70cc71ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52da9, value : 32'h100f11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52daa, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dab, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dac, value : 32'hf053e888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dad, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dae, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52daf, value : 32'h1008a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db0, value : 32'h52752},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db1, value : 32'h3000264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db2, value : 32'h33002e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db3, value : 32'h70c0704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db4, value : 32'h200572ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db5, value : 32'he090244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db6, value : 32'heab830d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db7, value : 32'h31310e17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db8, value : 32'h8080270b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52db9, value : 32'h1600f207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dba, value : 32'h80007081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dbb, value : 32'h95d0025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dbc, value : 32'he1b0050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dbd, value : 32'h220b3131},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dbe, value : 32'hf2098140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dbf, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc0, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc1, value : 32'h51090f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc2, value : 32'h2678f020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc3, value : 32'h794b3141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc4, value : 32'h215af41c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc5, value : 32'h41c32503},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc6, value : 32'h12e88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc7, value : 32'h71266a94},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc8, value : 32'h43c36179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dc9, value : 32'hff10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dca, value : 32'h43c3b166},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dcb, value : 32'h52c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dcc, value : 32'h1908639a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dcd, value : 32'h82e30003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dce, value : 32'h22058241},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dcf, value : 32'ha1e40102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd0, value : 32'h6462a141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd1, value : 32'ha1407a05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd2, value : 32'h31ff278d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd3, value : 32'h2640714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd4, value : 32'he79305e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd5, value : 32'h46c3b194},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd6, value : 32'h70000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd7, value : 32'h193e238d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd8, value : 32'h40c370ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dd9, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dda, value : 32'h841000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ddb, value : 32'h43c371cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ddc, value : 32'h54c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ddd, value : 32'h22e0c6b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dde, value : 32'h72ac700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ddf, value : 32'h72e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de0, value : 32'h2002014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de1, value : 32'h244ab80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de2, value : 32'h20057180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de3, value : 32'h4308025f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de4, value : 32'h3000264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de5, value : 32'h88020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de6, value : 32'h310c2e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de7, value : 32'h89086399},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de8, value : 32'h8000270b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52de9, value : 32'h215af218},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dea, value : 32'h40c32502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52deb, value : 32'h12e88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dec, value : 32'h60587126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ded, value : 32'h42c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dee, value : 32'hb0460ff1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52def, value : 32'h81218143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df0, value : 32'h7c12105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df1, value : 32'h1821808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df2, value : 32'h6461a021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df3, value : 32'h2c12105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df4, value : 32'ha020a044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df5, value : 32'h305e2640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df6, value : 32'h4bf258d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df7, value : 32'h7105710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df8, value : 32'h91140895},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52df9, value : 32'h41c34022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dfa, value : 32'h10068},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dfb, value : 32'h24120bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dfc, value : 32'hfa6f0df6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dfd, value : 32'h21424222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dfe, value : 32'h42d3a03c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52dff, value : 32'h12ec8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e00, value : 32'h2344f20b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e01, value : 32'h22402042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e02, value : 32'hd9f12140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e03, value : 32'h14020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e04, value : 32'h1814a822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e05, value : 32'h706d0092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e06, value : 32'h79eddff1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e07, value : 32'hfe2f0a76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e08, value : 32'h71654022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e09, value : 32'h14310b11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e0a, value : 32'h702c4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e0b, value : 32'h1a0082a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e0c, value : 32'h706dda10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e0d, value : 32'h7f0d6f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e0e, value : 32'h94120fe3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e0f, value : 32'h702c4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e10, value : 32'h1a00816},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e11, value : 32'h21424261},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e12, value : 32'hf20da03c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e13, value : 32'h2006710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e14, value : 32'h224004c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e15, value : 32'h20a82140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e16, value : 32'h180201c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e17, value : 32'h181403c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e18, value : 32'h706d0052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e19, value : 32'h4022df0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e1a, value : 32'hfe2f0a2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e1b, value : 32'h716541e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e1c, value : 32'h14310b11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e1d, value : 32'h712c4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e1e, value : 32'h1600fde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e1f, value : 32'h706dda10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e20, value : 32'h7f0d6f09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e21, value : 32'h9c3f278c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e22, value : 32'h4022f62f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e23, value : 32'hfca712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e24, value : 32'h42610160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e25, value : 32'h2030098f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e26, value : 32'h230a708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e27, value : 32'h702f3440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e28, value : 32'h350f215a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e29, value : 32'h23d32200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e2a, value : 32'h20d51308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e2b, value : 32'h23f10d1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e2c, value : 32'h20d61309},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e2d, value : 32'h14822730},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e2e, value : 32'hdb0f740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e2f, value : 32'h6341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e30, value : 32'he460003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e31, value : 32'h240afcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e32, value : 32'h268c0580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e33, value : 32'hf40dac7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e34, value : 32'h14822730},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e35, value : 32'h43a2740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e36, value : 32'h6441c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e37, value : 32'he2a0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e38, value : 32'h248afcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e39, value : 32'h26000c7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e3a, value : 32'h27302540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e3b, value : 32'h28441482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e3c, value : 32'h13040097},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e3d, value : 32'h252f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e3e, value : 32'he80705c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e3f, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e40, value : 32'h40065},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e41, value : 32'h740cf005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e42, value : 32'h6641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e43, value : 32'h43a20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e44, value : 32'hfcaf0df6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e45, value : 32'h580240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e46, value : 32'h238d7127},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e47, value : 32'h1b06313f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e48, value : 32'h402225c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e49, value : 32'h42009ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e4a, value : 32'hc809702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e4b, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e4c, value : 32'h78c50341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e4d, value : 32'h5041900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e4e, value : 32'h5041800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e4f, value : 32'he00e22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e50, value : 32'hc809710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e51, value : 32'h7d05b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e52, value : 32'h1d007e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e53, value : 32'h1e001045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e54, value : 32'hf0061045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e55, value : 32'h74041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e56, value : 32'hc02c9003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e57, value : 32'h2200db2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e58, value : 32'h4008710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e59, value : 32'h200e06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e5a, value : 32'h45cbd80d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e5b, value : 32'he008900f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e5c, value : 32'h255070cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e5d, value : 32'hb5c014cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e5e, value : 32'h13841b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e5f, value : 32'h200d8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e60, value : 32'h1d00c001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e61, value : 32'h8231404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e62, value : 32'h1b003031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e63, value : 32'hc8091404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e64, value : 32'h40c36832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e65, value : 32'hc400900f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e66, value : 32'h22105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e67, value : 32'h7825b8b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e68, value : 32'hb0c0b2c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e69, value : 32'h40c3f00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e6a, value : 32'hc02c9003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e6b, value : 32'hb8afb0c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e6c, value : 32'h70451e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e6d, value : 32'h802c9001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e6e, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e6f, value : 32'h1e0070cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e70, value : 32'h90037384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e71, value : 32'h1e00d878},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e72, value : 32'h90077384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e73, value : 32'hd42f87c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e74, value : 32'h40010220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e75, value : 32'h45cbd820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e76, value : 32'h3e09008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e77, value : 32'h200d2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e78, value : 32'h10451d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e79, value : 32'hd22d820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e7a, value : 32'hb5c00020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e7b, value : 32'hd80ac200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e7c, value : 32'h6f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e7d, value : 32'hd120002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e7e, value : 32'h4303fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e7f, value : 32'h1404c0a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e80, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e81, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e82, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e83, value : 32'h46303902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e84, value : 32'hb911d955},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e85, value : 32'h30001c84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e86, value : 32'h4078740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e87, value : 32'hfcaf0cea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e88, value : 32'hd9204450},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e89, value : 32'h89a0b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e8a, value : 32'h11002553},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e8b, value : 32'h8961a900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e8c, value : 32'h1002353},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e8d, value : 32'ha9017ba5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e8e, value : 32'h813e2353},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e8f, value : 32'h808c11f7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e90, value : 32'h11002453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e91, value : 32'h800219f7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e92, value : 32'h808211f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e93, value : 32'h1002253},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e94, value : 32'h800219f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e95, value : 32'h1901f405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e96, value : 32'h19000043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e97, value : 32'h7a850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e98, value : 32'h813e2253},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e99, value : 32'h19f8f405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e9a, value : 32'h19f78043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e9b, value : 32'h81b8043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e9c, value : 32'h740c3030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e9d, value : 32'h30710821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e9e, value : 32'hc8ed9ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52e9f, value : 32'hb910fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea0, value : 32'h706e70ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea1, value : 32'hd92bf00e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea2, value : 32'hfcaf0c7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea3, value : 32'h706eb912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea4, value : 32'hf00871ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea5, value : 32'hc72d9ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea6, value : 32'hb910fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea7, value : 32'h70ee716e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea8, value : 32'hbe9fdeee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ea9, value : 32'h16328ea0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eaa, value : 32'h70b51095},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eab, value : 32'h3a00c3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eac, value : 32'h202225ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ead, value : 32'h30001c9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eae, value : 32'hd957e812},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eaf, value : 32'hc4a740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb0, value : 32'hb911fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb1, value : 32'hb89fd825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb2, value : 32'h9b1000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb3, value : 32'h30412344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb4, value : 32'h885ba820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb5, value : 32'h412244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb6, value : 32'ha83b4158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb7, value : 32'h740cd9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb8, value : 32'hfcaf0c26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eb9, value : 32'h120cb910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eba, value : 32'h41c23085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ebb, value : 32'h30001484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ebc, value : 32'h43034282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ebd, value : 32'hfc2f0892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ebe, value : 32'h540240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ebf, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec0, value : 32'hb8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec1, value : 32'h3e0819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec2, value : 32'h740cd90b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec3, value : 32'hfcaf0bfa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec4, value : 32'h4062b914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec5, value : 32'he964182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec6, value : 32'h42e2fdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec7, value : 32'h24c02705},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec8, value : 32'h710853},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ec9, value : 32'h30001c88},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eca, value : 32'he8a58e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ecb, value : 32'h740cd9b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ecc, value : 32'hfcaf0bd6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ecd, value : 32'h2679b910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ece, value : 32'h40622003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ecf, value : 32'h4282702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed0, value : 32'h1200caa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed1, value : 32'h47084070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed2, value : 32'h4062e888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed3, value : 32'h4282712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed4, value : 32'h1200c9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed5, value : 32'h47084302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed6, value : 32'h740cd959},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed7, value : 32'hfcaf0baa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed8, value : 32'h4062b911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ed9, value : 32'he464182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eda, value : 32'h42e2fdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52edb, value : 32'hfe2f0f56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52edc, value : 32'h70d640e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52edd, value : 32'hfb220cb8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ede, value : 32'hb174082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52edf, value : 32'h740c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee0, value : 32'hb86d9b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee1, value : 32'hb910fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee2, value : 32'h48008fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee3, value : 32'hd92df057},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee4, value : 32'hfcaf0b76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee5, value : 32'h120cb912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee6, value : 32'h26793081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee7, value : 32'h25782003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee8, value : 32'h40e21004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ee9, value : 32'h4600e2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eea, value : 32'hca0c4282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eeb, value : 32'h5ca212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eec, value : 32'h2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eed, value : 32'h84d7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eee, value : 32'hd840003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eef, value : 32'hb89f70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef0, value : 32'h8820720e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef1, value : 32'h808d10e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef2, value : 32'hd237d25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef3, value : 32'h40e113ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef4, value : 32'h70911600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef5, value : 32'h48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef6, value : 32'hfbef0f72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef7, value : 32'h4200712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef8, value : 32'h4122700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ef9, value : 32'hfcef0c62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52efa, value : 32'h208d43e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52efb, value : 32'h71ed2c7f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52efc, value : 32'h740cd9b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52efd, value : 32'hfcaf0b12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52efe, value : 32'hcf6b910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52eff, value : 32'h4082fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f00, value : 32'h343206f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f01, value : 32'h10c29020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f02, value : 32'h9330700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f03, value : 32'he2f0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f04, value : 32'h16002011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f05, value : 32'h80007100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f06, value : 32'h9230188},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f07, value : 32'h8860005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f08, value : 32'h2005fccf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f09, value : 32'h81705c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f0a, value : 32'hd95b0071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f0b, value : 32'hada740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f0c, value : 32'hb911fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f0d, value : 32'hfb2f0dd6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f0e, value : 32'h8e004082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f0f, value : 32'hf47a7114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f10, value : 32'h7014ca06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f11, value : 32'h700cf276},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f12, value : 32'h20300e15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f13, value : 32'h30001c8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f14, value : 32'hfccf0852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f15, value : 32'h710ce804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f16, value : 32'h30001c8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f17, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f18, value : 32'h1700122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f19, value : 32'h262f1090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f1a, value : 32'h8f011407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f1b, value : 32'h38408c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f1c, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f1d, value : 32'h880012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f1e, value : 32'h3ae08b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f1f, value : 32'hea64082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f20, value : 32'h41c10220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f21, value : 32'h1ca0702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f22, value : 32'h14a03000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f23, value : 32'h8973000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f24, value : 32'h720c046e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f25, value : 32'h1c90704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f26, value : 32'hd8253000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f27, value : 32'h8820b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f28, value : 32'h7905881b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f29, value : 32'h2800710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f2a, value : 32'hb8020480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f2b, value : 32'h480200f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f2c, value : 32'hf231782b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f2d, value : 32'h300d148c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f2e, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f2f, value : 32'h791b28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f30, value : 32'h2002221f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f31, value : 32'hb82279aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f32, value : 32'h434278ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f33, value : 32'h704c6159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f34, value : 32'h40226119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f35, value : 32'h184209a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f36, value : 32'h41626038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f37, value : 32'h800070c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f38, value : 32'h1c941a44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f39, value : 32'h26793000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f3a, value : 32'h1c982000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f3b, value : 32'h14943000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f3c, value : 32'h98a3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f3d, value : 32'h14980460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f3e, value : 32'h14943004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f3f, value : 32'h41623000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f40, value : 32'h30041498},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f41, value : 32'h976714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f42, value : 32'h43420460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f43, value : 32'h71ad70b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f44, value : 32'h1490f3d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f45, value : 32'h714e3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f46, value : 32'h8837704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f47, value : 32'h1c908031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f48, value : 32'h71263000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f49, value : 32'ha2940967},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f4a, value : 32'hf19f7106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f4b, value : 32'hc00f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f4c, value : 32'h3000149c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f4d, value : 32'hf2e37014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f4e, value : 32'h3800996},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f4f, value : 32'h200f2679},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f50, value : 32'h30021c05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f51, value : 32'h416240a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f52, value : 32'hbd242e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f53, value : 32'hc380fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f54, value : 32'h740cd9b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f55, value : 32'hfcaf09b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f56, value : 32'h1488b910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f57, value : 32'he81a3000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f58, value : 32'h1243256f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f59, value : 32'h8dc0700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f5a, value : 32'hfbef0de2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f5b, value : 32'h4200712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f5c, value : 32'h41c1700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f5d, value : 32'hfcef0ad2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f5e, value : 32'h8da0706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f5f, value : 32'hdce710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f60, value : 32'h712cfbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f61, value : 32'h700c4200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f62, value : 32'habe41a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f63, value : 32'h716cfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f64, value : 32'h2144de40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f65, value : 32'hbe9f3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f66, value : 32'h2344ae00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f67, value : 32'hbed3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f68, value : 32'h1ee52030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f69, value : 32'hae29002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f6a, value : 32'h710cfd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f6b, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f6c, value : 32'h8d221b44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f6d, value : 32'h478b714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f6e, value : 32'h790a9706},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f6f, value : 32'h60389500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f70, value : 32'hb62790f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f71, value : 32'h710cfaaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f72, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f73, value : 32'h88422580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f74, value : 32'h794a9726},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f75, value : 32'h724c9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f76, value : 32'h790f6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f77, value : 32'hfaaf0b46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f78, value : 32'haa6710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f79, value : 32'h720cfd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f7a, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f7b, value : 32'h88422fbc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f7c, value : 32'h794a9726},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f7d, value : 32'h714c9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f7e, value : 32'h790f6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f7f, value : 32'hfaaf0b26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f80, value : 32'h40c3710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f81, value : 32'h39f88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f82, value : 32'h97268842},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f83, value : 32'h9000794a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f84, value : 32'h6038724c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f85, value : 32'hb0e790f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f86, value : 32'h710cfaaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f87, value : 32'hfd2f0a6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f88, value : 32'h120c730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f89, value : 32'h41c23085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f8a, value : 32'h30001484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f8b, value : 32'h43034282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f8c, value : 32'hfbef0d56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f8d, value : 32'hd917708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f8e, value : 32'h8ce740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f8f, value : 32'hb913fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f90, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f91, value : 32'h10b7122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f92, value : 32'h88810088},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f93, value : 32'hc6d8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f94, value : 32'h8351044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f95, value : 32'h244a106e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f96, value : 32'h700c7280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f97, value : 32'h50020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f98, value : 32'h209a68e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f99, value : 32'h211a0184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f9a, value : 32'hf82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f9b, value : 32'h60580a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f9c, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f9d, value : 32'h621a4434},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f9e, value : 32'h60b860b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52f9f, value : 32'h8802b260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa0, value : 32'h40e1aa02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa1, value : 32'hf1e57124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa2, value : 32'h3085120c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa3, value : 32'h148441c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa4, value : 32'h42823000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa5, value : 32'hcf24303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa6, value : 32'h708cfbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa7, value : 32'h740cd9b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa8, value : 32'hfcaf0866},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fa9, value : 32'h120cb910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52faa, value : 32'h40e23081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fab, value : 32'h43e14282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fac, value : 32'h4600b1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fad, value : 32'hf004708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fae, value : 32'h4400dca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52faf, value : 32'h30001488},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb0, value : 32'h256fe819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb1, value : 32'h700c1243},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb2, value : 32'hc828de0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb3, value : 32'h712cfbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb4, value : 32'h700c4200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb5, value : 32'h97241e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb6, value : 32'h706cfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb7, value : 32'h710c8da0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb8, value : 32'hfbef0c6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fb9, value : 32'h4200712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fba, value : 32'h41a1700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fbb, value : 32'hfcef095a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fbc, value : 32'h1e00716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fbd, value : 32'h1ee51642},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fbe, value : 32'h248096c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fbf, value : 32'h14043902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc0, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc1, value : 32'h68614200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc2, value : 32'h7054ca08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc3, value : 32'h20aa7b19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc4, value : 32'h81700c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc5, value : 32'h23ca003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc6, value : 32'h720c0021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc7, value : 32'hc420ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc8, value : 32'h20ab710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fc9, value : 32'hb1100c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fca, value : 32'h16000415},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fcb, value : 32'h901c7100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fcc, value : 32'hf01b0490},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fcd, value : 32'h10420aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fce, value : 32'ha1b7a12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fcf, value : 32'h24aa00e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd0, value : 32'h21aa1144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd1, value : 32'h8ff0104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd2, value : 32'h4b508044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd3, value : 32'h114424aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd4, value : 32'h6078f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd5, value : 32'h10421aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd6, value : 32'h20e17110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd7, value : 32'h22aa07c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd8, value : 32'hcf50144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fd9, value : 32'h7ee09080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fda, value : 32'h443226f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fdb, value : 32'h8a004300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fdc, value : 32'ha0f239a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fdd, value : 32'h802079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fde, value : 32'h12fe6822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fdf, value : 32'h78398100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe0, value : 32'h70002e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe1, value : 32'h4240000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe2, value : 32'hffef077d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe3, value : 32'h2b05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe4, value : 32'h826c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe5, value : 32'hf720000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe6, value : 32'hc0d1ffcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe7, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe8, value : 32'h4328c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fe9, value : 32'h200812},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fea, value : 32'h7071702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52feb, value : 32'h7fe0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fec, value : 32'h2c520ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fed, value : 32'h343226f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fee, value : 32'h370d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fef, value : 32'h92600d41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff0, value : 32'hf8628c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff1, value : 32'h86a00001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff2, value : 32'hc620da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff3, value : 32'h52628c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff4, value : 32'hc520da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff5, value : 32'hf8528c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff6, value : 32'h8480001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff7, value : 32'h69818a62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff8, value : 32'h71046078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ff9, value : 32'hc02805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ffa, value : 32'h800043c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ffb, value : 32'h8b601140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ffc, value : 32'h12fbeb0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ffd, value : 32'ha178082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52ffe, value : 32'h43c300df},
                          '{ step_type : REG_WRITE, reg_addr : 32'h52fff, value : 32'h12268000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53000, value : 32'hea058b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53001, value : 32'h8b817a2c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53002, value : 32'h74107c4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53003, value : 32'h20ca7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53004, value : 32'h78e0030d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53005, value : 32'h83ac2ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53006, value : 32'h2053fe0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53007, value : 32'h206d00c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53008, value : 32'h50160900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53009, value : 32'h43d3782a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5300a, value : 32'h3f8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5300b, value : 32'h13005015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5300c, value : 32'h13012080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5300d, value : 32'he9102081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5300e, value : 32'h2079d953},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5300f, value : 32'hdaa0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53010, value : 32'hb913fa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53011, value : 32'h1300ca14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53012, value : 32'hb8022081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53013, value : 32'h80206c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53014, value : 32'hf0136119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53015, value : 32'h29941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53016, value : 32'hd8e0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53017, value : 32'h2078fa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53018, value : 32'h16000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53019, value : 32'h80007081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5301a, value : 32'hc8060024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5301b, value : 32'h91080b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5301c, value : 32'h781dc805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5301d, value : 32'h7a2f5015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5301e, value : 32'h807e2153},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5301f, value : 32'h832a41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53020, value : 32'h23c0ba23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53021, value : 32'h21530062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53022, value : 32'h1a028080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53023, value : 32'h22c03002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53024, value : 32'hd80a0062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53025, value : 32'h29a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53026, value : 32'h1a010002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53027, value : 32'he6a30c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53028, value : 32'h1a00fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53029, value : 32'h276f3082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5302a, value : 32'h41c310c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5302b, value : 32'h6029c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5302c, value : 32'hb8e28f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5302d, value : 32'h20cad87f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5302e, value : 32'h1a0301e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5302f, value : 32'hd80a3002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53030, value : 32'h14861705},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53031, value : 32'h11071700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53032, value : 32'h1085170c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53033, value : 32'h1104170a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53034, value : 32'h20831301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53035, value : 32'hfc6f0e32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53036, value : 32'h8f1f8f5f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53037, value : 32'hf28db8e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53038, value : 32'hd80ade66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53039, value : 32'h41c3be9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5303a, value : 32'h502a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5303b, value : 32'h948616fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5303c, value : 32'h948516fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5303d, value : 32'h10841600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5303e, value : 32'h908316fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5303f, value : 32'h908216a6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53040, value : 32'hfc6f0e06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53041, value : 32'h2640bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53042, value : 32'h8e6c1610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53043, value : 32'h20861000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53044, value : 32'h2a645cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53045, value : 32'h10fc0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53046, value : 32'hd80aa085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53047, value : 32'ha08410f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53048, value : 32'h16a641a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53049, value : 32'hde29082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5304a, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5304b, value : 32'h24122040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5304c, value : 32'h20831004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5304d, value : 32'h20861200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5304e, value : 32'h1401254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5304f, value : 32'ha08512fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53050, value : 32'h12f8d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53051, value : 32'h16a6a084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53052, value : 32'hdbe9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53053, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53054, value : 32'h24112240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53055, value : 32'h20831204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53056, value : 32'h24861110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53057, value : 32'h11ecd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53058, value : 32'h41c3a085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53059, value : 32'h502a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5305a, value : 32'ha08411e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5305b, value : 32'h16a64030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5305c, value : 32'hd969082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5305d, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5305e, value : 32'ha48611fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5305f, value : 32'h2401204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53060, value : 32'h20851100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53061, value : 32'h11fcd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53062, value : 32'h11f8a084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53063, value : 32'h16a6a083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53064, value : 32'hd769082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53065, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53066, value : 32'h250d2140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53067, value : 32'h20831108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53068, value : 32'h10861500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53069, value : 32'h2441204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5306a, value : 32'h908515fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5306b, value : 32'h15f8d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5306c, value : 32'h40309084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5306d, value : 32'h908216a6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5306e, value : 32'hfc6f0d4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5306f, value : 32'h1510bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53070, value : 32'h204f1086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53071, value : 32'h150c2401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53072, value : 32'hd80a1085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53073, value : 32'h10841508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53074, value : 32'h16a68d64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53075, value : 32'hd329082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53076, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53077, value : 32'h10841518},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53078, value : 32'h8d74d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53079, value : 32'h2ac41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5307a, value : 32'h16a60003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5307b, value : 32'hd1a9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5307c, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5307d, value : 32'hb8e18f1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5307e, value : 32'hde67f287},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5307f, value : 32'hbe9fd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53080, value : 32'h2af41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53081, value : 32'h16fc0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53082, value : 32'h16fc9486},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53083, value : 32'h16009485},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53084, value : 32'h16fc1084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53085, value : 32'h16a59083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53086, value : 32'hcee9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53087, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53088, value : 32'h160d2640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53089, value : 32'h15108e6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5308a, value : 32'hd80a1486},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5308b, value : 32'h908515ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5308c, value : 32'h2b041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5308d, value : 32'h15e80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5308e, value : 32'h40309084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5308f, value : 32'h908216a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53090, value : 32'hfc6f0cc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53091, value : 32'h15fcbac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53092, value : 32'h204f9486},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53093, value : 32'h15142401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53094, value : 32'hd80a1485},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53095, value : 32'h908415e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53096, value : 32'h908315e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53097, value : 32'h908216a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53098, value : 32'hfc6f0ca6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53099, value : 32'h15fcbac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5309a, value : 32'h204f9486},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5309b, value : 32'h15002441},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5309c, value : 32'hd80a1085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5309d, value : 32'h908415fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5309e, value : 32'h15f84230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5309f, value : 32'h16a59083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a0, value : 32'hc869082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a1, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a2, value : 32'h15112540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a3, value : 32'h11008d68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a4, value : 32'h224f2086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a5, value : 32'h11fc2401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a6, value : 32'hd80aa085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a7, value : 32'ha08411f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a8, value : 32'h908216a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530a9, value : 32'hfc6f0c62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530aa, value : 32'h2140bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ab, value : 32'h1104240d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ac, value : 32'h15002083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ad, value : 32'h204f1086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ae, value : 32'h15fc2481},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530af, value : 32'hd80a9085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b0, value : 32'h908415f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b1, value : 32'h16a54030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b2, value : 32'hc3e9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b3, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b4, value : 32'h10861510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b5, value : 32'h2401204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b6, value : 32'h1085150c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b7, value : 32'h1508d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b8, value : 32'h8d641084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530b9, value : 32'h908216a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ba, value : 32'hfc6f0c1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530bb, value : 32'h1518bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530bc, value : 32'hd80a1084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530bd, value : 32'h41c38d74},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530be, value : 32'h302b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530bf, value : 32'h908216a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c0, value : 32'hfc6f0c06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c1, value : 32'h1301bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c2, value : 32'hb8e02080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c3, value : 32'hde68f28c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c4, value : 32'hbe9fd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c5, value : 32'h2b941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c6, value : 32'h16fc0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c7, value : 32'h16fc9486},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c8, value : 32'h16189485},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530c9, value : 32'h16e41484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ca, value : 32'h168c9083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530cb, value : 32'hbda9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530cc, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530cd, value : 32'h948616fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ce, value : 32'h2ba45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530cf, value : 32'h16000005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d0, value : 32'hd80a1085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d1, value : 32'h908416fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d2, value : 32'h16f841a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d3, value : 32'h16909083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d4, value : 32'hbb69082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d5, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d6, value : 32'h15102640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d7, value : 32'h10008e68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d8, value : 32'h254f2086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530d9, value : 32'h10fc1401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530da, value : 32'hd80aa085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530db, value : 32'ha08410f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530dc, value : 32'h90821690},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530dd, value : 32'hfc6f0b92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530de, value : 32'h2040bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530df, value : 32'h1004240d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e0, value : 32'h15002083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e1, value : 32'hd80a1086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e2, value : 32'h908515fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e3, value : 32'h2bc41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e4, value : 32'h15f80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e5, value : 32'h40309084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e6, value : 32'h90821690},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e7, value : 32'hfc6f0b6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e8, value : 32'h2540bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530e9, value : 32'h8d641411},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ea, value : 32'h20861100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530eb, value : 32'h2401204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ec, value : 32'ha08511fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ed, value : 32'h11f8d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ee, value : 32'h1690a084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ef, value : 32'hb4a9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f0, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f1, value : 32'h240d2140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f2, value : 32'h20831104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f3, value : 32'h10861500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f4, value : 32'h2441204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f5, value : 32'h908515fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f6, value : 32'h15f8d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f7, value : 32'h40309084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f8, value : 32'h90821690},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530f9, value : 32'hfc6f0b22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530fa, value : 32'h1510bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530fb, value : 32'h204f1086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530fc, value : 32'h150c2401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530fd, value : 32'hd80a1085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530fe, value : 32'h10841508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h530ff, value : 32'h16908d64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53100, value : 32'hb069082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53101, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53102, value : 32'h10841518},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53103, value : 32'h8d74d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53104, value : 32'h2c041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53105, value : 32'h16900003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53106, value : 32'haee9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53107, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53108, value : 32'h20801301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53109, value : 32'hf28eb8e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5310a, value : 32'hd80ade69},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5310b, value : 32'h41c3be9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5310c, value : 32'h502c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5310d, value : 32'h948616fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5310e, value : 32'h948516fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5310f, value : 32'h10841600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53110, value : 32'h908316fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53111, value : 32'h908216a3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53112, value : 32'hfc6f0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53113, value : 32'h2640bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53114, value : 32'h8e6c1610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53115, value : 32'h20861000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53116, value : 32'h2c445cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53117, value : 32'h10fc0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53118, value : 32'hd80aa085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53119, value : 32'ha08410f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5311a, value : 32'h16a341a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5311b, value : 32'ha9a9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5311c, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5311d, value : 32'h24112040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5311e, value : 32'h20831004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5311f, value : 32'h20861100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53120, value : 32'h1401254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53121, value : 32'ha08511fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53122, value : 32'h11f8d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53123, value : 32'h16a3a084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53124, value : 32'ha769082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53125, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53126, value : 32'h24122140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53127, value : 32'h20831104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53128, value : 32'h20861200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53129, value : 32'h12fcbd91},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5312a, value : 32'hd80aa085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5312b, value : 32'ha08412f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5312c, value : 32'h16a341a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5312d, value : 32'ha529082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5312e, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5312f, value : 32'h24102240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53130, value : 32'h20831204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53131, value : 32'h20861000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53132, value : 32'h1401254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53133, value : 32'ha08510fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53134, value : 32'h10f8d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53135, value : 32'h16a3a084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53136, value : 32'ha2e9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53137, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53138, value : 32'h240d2040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53139, value : 32'h20831004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5313a, value : 32'h14861510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5313b, value : 32'h15ecd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5313c, value : 32'h41c39085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5313d, value : 32'h502c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5313e, value : 32'h908415e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5313f, value : 32'h16a34030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53140, value : 32'ha069082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53141, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53142, value : 32'h948615fc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53143, value : 32'h2401204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53144, value : 32'h10851500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53145, value : 32'h15fcd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53146, value : 32'h15f89084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53147, value : 32'h16a39083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53148, value : 32'h9e69082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53149, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5314a, value : 32'h1084150c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5314b, value : 32'h8d68d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5314c, value : 32'h2ca41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5314d, value : 32'h16a30003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5314e, value : 32'h9ce9082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5314f, value : 32'hbac3fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53150, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53151, value : 32'h2009030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53152, value : 32'hb822710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53153, value : 32'h20002006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53154, value : 32'h30021a08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53155, value : 32'h82f9700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53156, value : 32'hf85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53157, value : 32'hc8090a6b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53158, value : 32'h7200244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53159, value : 32'h700c6852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5315a, value : 32'h34020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5315b, value : 32'h12205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5315c, value : 32'h70c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5315d, value : 32'h21054000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5315e, value : 32'h90380f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5315f, value : 32'h1900004c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53160, value : 32'he360404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53161, value : 32'h46cbfe0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53162, value : 32'hc1dc901f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53163, value : 32'h1443256f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53164, value : 32'h74041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53165, value : 32'h4a0901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53166, value : 32'h74041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53167, value : 32'hc294900b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53168, value : 32'h10051e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53169, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5316a, value : 32'h102cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5316b, value : 32'hfc6f095a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5316c, value : 32'h8ea8d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5316d, value : 32'h8d00faef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5316e, value : 32'h750cd92d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5316f, value : 32'hfc6f094a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53170, value : 32'h1e24b914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53171, value : 32'h97051404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53172, value : 32'h500813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53173, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53174, value : 32'h48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53175, value : 32'h98cb8e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53176, value : 32'h16000101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53177, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53178, value : 32'h70140114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53179, value : 32'h1820c7c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5317a, value : 32'h78e0c6ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5317b, value : 32'hcb2c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5317c, value : 32'h40c3fa4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5317d, value : 32'hbb80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5317e, value : 32'hffef09aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5317f, value : 32'h252f702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53180, value : 32'hf20d9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53181, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53182, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53183, value : 32'h73ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53184, value : 32'hfaaf0cd2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53185, value : 32'h258c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53186, value : 32'hd8801e3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53187, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53188, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53189, value : 32'hcbe73ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5318a, value : 32'h70ccfaaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5318b, value : 32'hc66700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5318c, value : 32'h712cfaaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5318d, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5318e, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5318f, value : 32'h4610b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53190, value : 32'h70c01600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53191, value : 32'h1f8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53192, value : 32'h320819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53193, value : 32'h34ad2496},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53194, value : 32'h200e66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53195, value : 32'h249640c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53196, value : 32'h14043b92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53197, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53198, value : 32'h740cde51},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53199, value : 32'h8a2be13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5319a, value : 32'h41c1fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5319b, value : 32'h800041d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5319c, value : 32'h1101122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5319d, value : 32'h24002090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5319e, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5319f, value : 32'h702c014c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a0, value : 32'ha7eda24},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a1, value : 32'h1100f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a2, value : 32'h1600208d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a3, value : 32'h80007093},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a4, value : 32'h2344001f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a5, value : 32'h264f2140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a6, value : 32'hf4e1401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a7, value : 32'h2079f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a8, value : 32'h23440140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531a9, value : 32'h23442040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531aa, value : 32'hc0442092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ab, value : 32'h21002344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ac, value : 32'h242fc043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ad, value : 32'hc3030482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ae, value : 32'hc204740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531af, value : 32'h28a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b0, value : 32'h8460003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b1, value : 32'hbb22fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b2, value : 32'h6832c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b3, value : 32'hf802105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b4, value : 32'h89038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b5, value : 32'h275390e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b6, value : 32'hf4129080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b7, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b8, value : 32'h1f8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531b9, value : 32'h720cb8e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ba, value : 32'h6120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531bb, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531bc, value : 32'hc008903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531bd, value : 32'h27537f05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531be, value : 32'hb1e01080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531bf, value : 32'h50080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c0, value : 32'h80b10857},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c1, value : 32'hf003720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c2, value : 32'hc045710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c3, value : 32'hc04178bb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c4, value : 32'h2014710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c5, value : 32'h236d0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c6, value : 32'h41c32902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c7, value : 32'h1028b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c8, value : 32'h740cc049},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531c9, value : 32'hfc2f0fe2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ca, value : 32'had24550},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531cb, value : 32'h40c201a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531cc, value : 32'h212f70ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531cd, value : 32'hbee05c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ce, value : 32'h40c201e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531cf, value : 32'h230e2f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d0, value : 32'h70ad4018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d1, value : 32'h336e08c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d2, value : 32'h12102d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d3, value : 32'h2500275a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d4, value : 32'h23902005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d5, value : 32'h728e706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d6, value : 32'h70c378b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d7, value : 32'h4db48001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d8, value : 32'h4051800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531d9, value : 32'h24554162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531da, value : 32'h219f3bc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531db, value : 32'h23000201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531dc, value : 32'h2340240b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531dd, value : 32'h275a1482},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531de, value : 32'h43c32488},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531df, value : 32'h9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e0, value : 32'h603c44a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e1, value : 32'h7a05c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e2, value : 32'hba027401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e3, value : 32'h7a657cb4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e4, value : 32'h1061200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e5, value : 32'h6159c28b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e6, value : 32'h14022340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e7, value : 32'h1c007845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e8, value : 32'hb8021184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531e9, value : 32'h78657101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ea, value : 32'h100079b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531eb, value : 32'h740c0105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ec, value : 32'h1441900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ed, value : 32'h28c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ee, value : 32'h42620005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ef, value : 32'hfc2f0f4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f0, value : 32'hd4543e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f1, value : 32'h40c32051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f2, value : 32'ha3c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f3, value : 32'h2001271a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f4, value : 32'h231fb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f5, value : 32'h60382000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f6, value : 32'h219a41a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f7, value : 32'h61190184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f8, value : 32'h2005c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531f9, value : 32'h21000400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531fa, value : 32'h80000f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531fb, value : 32'hb8021b48},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531fc, value : 32'h800071c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531fd, value : 32'h20056d28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531fe, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h531ff, value : 32'h90000320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53200, value : 32'hb100b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53201, value : 32'h2c3e248d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53202, value : 32'h71a5716e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53203, value : 32'h92540d39},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53204, value : 32'hf2371e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53205, value : 32'h244aa114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53206, value : 32'hd8987140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53207, value : 32'h24020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53208, value : 32'hf812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53209, value : 32'hc000903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5320a, value : 32'h19007404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5320b, value : 32'hd1300c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5320c, value : 32'h257820b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5320d, value : 32'h46cb2041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5320e, value : 32'h835c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5320f, value : 32'h46cbf004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53210, value : 32'h24b00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53211, value : 32'h20c02a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53212, value : 32'h46cbe904},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53213, value : 32'h2f540001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53214, value : 32'h1002052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53215, value : 32'h8b6c047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53216, value : 32'h700cfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53217, value : 32'h41db710f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53218, value : 32'h50290},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53219, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5321a, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5321b, value : 32'hc008903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5321c, value : 32'h3051080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5321d, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5321e, value : 32'hf005d8a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5321f, value : 32'h1451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53220, value : 32'h141cd8a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53221, value : 32'h706f3010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53222, value : 32'hc809c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53223, value : 32'h7140244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53224, value : 32'h20a8c202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53225, value : 32'h220504c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53226, value : 32'he2100001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53227, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53228, value : 32'h903b0f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53229, value : 32'h2105c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5322a, value : 32'h903b0f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5322b, value : 32'h1b00c004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5322c, value : 32'h19000404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5322d, value : 32'h16000404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5322e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5322f, value : 32'h8110001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53230, value : 32'hdd6400bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53231, value : 32'h708d1600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53232, value : 32'h1208000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53233, value : 32'he88ac003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53234, value : 32'h742cd80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53235, value : 32'h716c42c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53236, value : 32'haae44a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53237, value : 32'h70acfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53238, value : 32'he88ac004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53239, value : 32'h742cd80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5323a, value : 32'h706c42c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5323b, value : 32'ha9a44a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5323c, value : 32'h70acfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5323d, value : 32'h70ae720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5323e, value : 32'hc048c046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5323f, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53240, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53241, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53242, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53243, value : 32'h710c7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53244, value : 32'h5402800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53245, value : 32'h200fb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53246, value : 32'h782b0540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53247, value : 32'h740cf293},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53248, value : 32'h28d41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53249, value : 32'h42030003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5324a, value : 32'hdde4302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5324b, value : 32'h240afc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5324c, value : 32'h11000540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5324d, value : 32'h11012092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5324e, value : 32'h220c2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5324f, value : 32'h106a000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53250, value : 32'h40c3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53251, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53252, value : 32'h8f78800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53253, value : 32'h212f04ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53254, value : 32'h9d20487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53255, value : 32'h40c201e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53256, value : 32'h242f70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53257, value : 32'hc04a2488},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53258, value : 32'h8d9c00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53259, value : 32'h232f036e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5325a, value : 32'hc0042348},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5325b, value : 32'hc003e8ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5325c, value : 32'h40a2e8b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5325d, value : 32'h42624182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5325e, value : 32'h706c7e60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5325f, value : 32'h740c4710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53260, value : 32'h42424123},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53261, value : 32'h44a143a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53262, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53263, value : 32'hfc2f0d7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53264, value : 32'h5c0260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53265, value : 32'h418240a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53266, value : 32'h7e604262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53267, value : 32'h4310716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53268, value : 32'h3401214f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53269, value : 32'h4242740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5326a, value : 32'h44a143a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5326b, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5326c, value : 32'hfc2f0d56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5326d, value : 32'h4c0260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5326e, value : 32'ha5c0230c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5326f, value : 32'h24c527ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53270, value : 32'h40a2f01f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53271, value : 32'h42624182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53272, value : 32'h706c7e60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53273, value : 32'h740c4710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53274, value : 32'h28e41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53275, value : 32'hf00c0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53276, value : 32'h418240a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53277, value : 32'h7e604262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53278, value : 32'h4710716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53279, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5327a, value : 32'h5028f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5327b, value : 32'h43a24242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5327c, value : 32'h250a44a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5327d, value : 32'hd120400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5327e, value : 32'h260afc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5327f, value : 32'h410205c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53280, value : 32'h219a42a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53281, value : 32'h24560804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53282, value : 32'h229f3b80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53283, value : 32'h43a20402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53284, value : 32'h250a44a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53285, value : 32'h260a0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53286, value : 32'h603805c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53287, value : 32'h225a6059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53288, value : 32'h42422900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53289, value : 32'h41c36038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5328a, value : 32'h50292},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5328b, value : 32'h180078b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5328c, value : 32'hcd605c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5328d, value : 32'h740cfc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5328e, value : 32'hd2971a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5328f, value : 32'h71469254},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53290, value : 32'hc008f17b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53291, value : 32'h770471ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53292, value : 32'hc0487014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53293, value : 32'h7106f558},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53294, value : 32'ha800204c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53295, value : 32'hffc50636},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53296, value : 32'h70811600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53297, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53298, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53299, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5329a, value : 32'h710c7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5329b, value : 32'h6c02800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5329c, value : 32'h200fb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5329d, value : 32'h782b06c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5329e, value : 32'h1100f27b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5329f, value : 32'h11012092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a0, value : 32'h8e12080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a1, value : 32'h406304a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a2, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a3, value : 32'h880012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a4, value : 32'h4ae08cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a5, value : 32'h7240244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a6, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a7, value : 32'h14c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a8, value : 32'h10020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532a9, value : 32'h111804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532aa, value : 32'h487212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ab, value : 32'h1e00876},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ac, value : 32'h141c40c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ad, value : 32'h43103010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ae, value : 32'hb6d70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532af, value : 32'h4102236e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b0, value : 32'h219a4263},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b1, value : 32'h24560804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b2, value : 32'h229f3b80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b3, value : 32'h60380402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b4, value : 32'h225a6059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b5, value : 32'h60382900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b6, value : 32'h3f812400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b7, value : 32'h14c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b8, value : 32'h34720f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532b9, value : 32'h2500225a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ba, value : 32'h814079b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532bb, value : 32'h70c378b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532bc, value : 32'h4db48001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532bd, value : 32'h1c50a13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532be, value : 32'h4041800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532bf, value : 32'h400242e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c0, value : 32'h1c01900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c1, value : 32'h9000f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c2, value : 32'h262fc240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c3, value : 32'h740c0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c4, value : 32'h29341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c5, value : 32'h42630007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c6, value : 32'h44a14342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c7, value : 32'hfc2f0bea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c8, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532c9, value : 32'hd9771a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ca, value : 32'h71069254},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532cb, value : 32'ha814088d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532cc, value : 32'h240070ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532cd, value : 32'h3f90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ce, value : 32'hb1d014c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532cf, value : 32'h4006234e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d0, value : 32'h700ce88a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d1, value : 32'h29441c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d2, value : 32'h42630003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d3, value : 32'ha9a4342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d4, value : 32'h44a1f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d5, value : 32'hde771a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d6, value : 32'h74069274},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d7, value : 32'hf1917146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d8, value : 32'h42c3c102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532d9, value : 32'hb5bc0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532da, value : 32'h3e00d2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532db, value : 32'hc00643c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532dc, value : 32'h7704716f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532dd, value : 32'hc0467014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532de, value : 32'hc005f570},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532df, value : 32'hb000200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e0, value : 32'hffe504e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e1, value : 32'h70ad7107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e2, value : 32'hf9a79af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e3, value : 32'h40c201a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e4, value : 32'h13112d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e5, value : 32'h706e4608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e6, value : 32'h14ee0e79},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e7, value : 32'h22102b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e8, value : 32'h2005704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532e9, value : 32'h724e2450},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ea, value : 32'h255a4448},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532eb, value : 32'h249f1488},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ec, value : 32'h24551201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ed, value : 32'h22003bc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ee, value : 32'h43c3040b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ef, value : 32'h9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f0, value : 32'h14812340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f1, value : 32'h4c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f2, value : 32'h20006098},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f3, value : 32'hc8090209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f4, value : 32'h21f47905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f5, value : 32'hb90214c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f6, value : 32'h19007965},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f7, value : 32'h23400184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f8, value : 32'h78251401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532f9, value : 32'h7b05b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532fa, value : 32'h6098c08b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532fb, value : 32'h20f47001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532fc, value : 32'hb32004c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532fd, value : 32'h29541c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532fe, value : 32'h20f40005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h532ff, value : 32'h740c04c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53300, value : 32'h14c621f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53301, value : 32'hfc2f0b02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53302, value : 32'h228d43a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53303, value : 32'h714c243f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53304, value : 32'hb897166},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53305, value : 32'h71a5a254},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53306, value : 32'h91140d71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53307, value : 32'h81240c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53308, value : 32'h712c03a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53309, value : 32'h790fc009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5330a, value : 32'h780fc001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5330b, value : 32'h40927},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5330c, value : 32'h6852c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5330d, value : 32'hb8c4c001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5330e, value : 32'h7845b80e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5330f, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53310, value : 32'h89038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53311, value : 32'hc001b0e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53312, value : 32'hc0417104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53313, value : 32'h9e9780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53314, value : 32'h16008005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53315, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53316, value : 32'hb8e60164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53317, value : 32'h1600f42a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53318, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53319, value : 32'h83b001f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5331a, value : 32'h740c00ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5331b, value : 32'h29641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5331c, value : 32'ha960000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5331d, value : 32'h256ffc0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5331e, value : 32'hd80f1a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5331f, value : 32'h42c2742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53320, value : 32'hd86716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53321, value : 32'h1d00ff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53322, value : 32'hd80f1205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53323, value : 32'h42c2742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53324, value : 32'hff6f0d76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53325, value : 32'hd808706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53326, value : 32'hb500b88f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53327, value : 32'h41c3f00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53328, value : 32'h297},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53329, value : 32'hfc2f0a62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5332a, value : 32'hc06740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5332b, value : 32'h40c2fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5332c, value : 32'hffcf01a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5332d, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5332e, value : 32'hc1bfb6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5332f, value : 32'hc8094410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53330, value : 32'h24056892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53331, value : 32'h90381f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53332, value : 32'h90e00008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53333, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53334, value : 32'h1648000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53335, value : 32'h90832753},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53336, value : 32'h40c3c045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53337, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53338, value : 32'h88218840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53339, value : 32'h1600f411},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5333a, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5333b, value : 32'hb8e6001f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5333c, value : 32'h20ca720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5333d, value : 32'h24050061},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5333e, value : 32'h903b1f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5333f, value : 32'h7f05c008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53340, value : 32'h2753b3e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53341, value : 32'hb111083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53342, value : 32'h710c0070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53343, value : 32'h3227274},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53344, value : 32'h720c0022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53345, value : 32'h71adc043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53346, value : 32'h7d34c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53347, value : 32'h7e5b780d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53348, value : 32'h2044c049},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53349, value : 32'hc0478800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5334a, value : 32'h244af40d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5334b, value : 32'hd8987140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5334c, value : 32'h24020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5334d, value : 32'hf812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5334e, value : 32'hc000903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5334f, value : 32'h19007404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53350, value : 32'hcba00c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53351, value : 32'h40820160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53352, value : 32'h716fd825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53353, value : 32'h8820b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53354, value : 32'h7825881b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53355, value : 32'hc02078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53356, value : 32'hc0487104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53357, value : 32'hc04178af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53358, value : 32'hc04678cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53359, value : 32'h36c7212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5335a, value : 32'h7033c003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5335b, value : 32'h250236},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5335c, value : 32'hc8094082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5335d, value : 32'hb802752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5335e, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5335f, value : 32'hc008903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53360, value : 32'h30710915},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53361, value : 32'h712cc144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53362, value : 32'h2802218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53363, value : 32'h730cb020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53364, value : 32'hf00ac040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53365, value : 32'h1451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53366, value : 32'h218a740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53367, value : 32'hc0402902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53368, value : 32'hc044760c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53369, value : 32'hc00870ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5336a, value : 32'h1f47510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5336b, value : 32'hc0070006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5336c, value : 32'h10182578},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5336d, value : 32'h2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5336e, value : 32'h30182004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5336f, value : 32'h30402178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53370, value : 32'h30182004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53371, value : 32'h3071081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53372, value : 32'h7140244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53373, value : 32'h20a8d898},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53374, value : 32'h20050280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53375, value : 32'h903b0f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53376, value : 32'h7404c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53377, value : 32'h51900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53378, value : 32'hfcaf0b2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53379, value : 32'h1400710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5337a, value : 32'h272f3004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5337b, value : 32'hd8c82347},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5337c, value : 32'h4218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5337d, value : 32'h42c34382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5337e, value : 32'hb5bc0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5337f, value : 32'h5c0250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53380, value : 32'hee270cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53381, value : 32'h43500260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53382, value : 32'h40d3c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53383, value : 32'h4db48001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53384, value : 32'hff0841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53385, value : 32'h3b152440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53386, value : 32'h220a74ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53387, value : 32'h40a22400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53388, value : 32'hac64142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53389, value : 32'hda14f9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5338a, value : 32'h25152540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5338b, value : 32'h2e7f268d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5338c, value : 32'h25122240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5338d, value : 32'h30041410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5338e, value : 32'h218ad8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5338f, value : 32'h42620004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53390, value : 32'h250a4382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53391, value : 32'he9e05c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53392, value : 32'h70cc0260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53393, value : 32'hf005c28b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53394, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53395, value : 32'h746cbf6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53396, value : 32'h7280244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53397, value : 32'h28020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53398, value : 32'h21011000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53399, value : 32'h5001202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5339a, value : 32'h781d6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5339b, value : 32'h20141802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5339c, value : 32'hd3f238c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5339d, value : 32'hfcaf0a96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5339e, value : 32'h4082700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5339f, value : 32'h3600db2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a0, value : 32'h7017702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a1, value : 32'h70ce706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a2, value : 32'h244af284},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a3, value : 32'hd9987140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a4, value : 32'h24020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a5, value : 32'hf802105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a6, value : 32'hc000903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a7, value : 32'h18007424},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a8, value : 32'h73ce04c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533a9, value : 32'hc809f076},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533aa, value : 32'h7140244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ab, value : 32'h3422005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ac, value : 32'h20a84122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ad, value : 32'h220503c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ae, value : 32'he1100040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533af, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b0, value : 32'h903b0f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b1, value : 32'h700cc000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b2, value : 32'h1b00c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b3, value : 32'h14000005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b4, value : 32'h40223004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b5, value : 32'h30061424},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b6, value : 32'h26bfd910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b7, value : 32'h42c30fff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b8, value : 32'h27980000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533b9, value : 32'hdfe4382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ba, value : 32'h250a0260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533bb, value : 32'h203c05c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533bc, value : 32'h14182580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533bd, value : 32'hc04a3010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533be, value : 32'h897c001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533bf, value : 32'hc0020404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c0, value : 32'h402212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c1, value : 32'h2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c2, value : 32'h2840b9c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c3, value : 32'h40820095},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c4, value : 32'h1a00c12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c5, value : 32'h2840704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c6, value : 32'h5021230c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c7, value : 32'h13422405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c8, value : 32'h22054322},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533c9, value : 32'h20440048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ca, value : 32'h21402041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533cb, value : 32'ha57010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533cc, value : 32'h84b22c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533cd, value : 32'h2005056e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ce, value : 32'h42c310c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533cf, value : 32'h9038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d0, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d1, value : 32'h11000089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d2, value : 32'hc10a1106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d3, value : 32'hb040200b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d4, value : 32'h2240f215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d5, value : 32'h79852981},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d6, value : 32'h7a25b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d7, value : 32'hc12653},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d8, value : 32'h3f1091b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533d9, value : 32'h1071200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533da, value : 32'hf00f13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533db, value : 32'h412740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533dc, value : 32'h11841900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533dd, value : 32'h1900b220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533de, value : 32'he3101005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533df, value : 32'h71a67146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e0, value : 32'hc002f1d7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e1, value : 32'h20527106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e2, value : 32'hc0420000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e3, value : 32'h7166f1b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e4, value : 32'h24c7202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e5, value : 32'ha4050e13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e6, value : 32'hf10771a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e7, value : 32'hffef05c9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e8, value : 32'hc8e7167},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533e9, value : 32'h712c0360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ea, value : 32'hc001c106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533eb, value : 32'h440825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ec, value : 32'h6832c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ed, value : 32'h11002653},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ee, value : 32'hb80e71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ef, value : 32'h78257acf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f0, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f1, value : 32'h89038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f2, value : 32'hc001b0e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f3, value : 32'h808508e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f4, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f5, value : 32'h1648000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f6, value : 32'h19f0857},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f7, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f8, value : 32'h1f8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533f9, value : 32'hff0839},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533fa, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533fb, value : 32'h286},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533fc, value : 32'hfbcf0f16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533fd, value : 32'h1a43256f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533fe, value : 32'h742cd80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h533ff, value : 32'h716c4282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53400, value : 32'hff6f0a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53401, value : 32'h12051d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53402, value : 32'h742cd80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53403, value : 32'h9fa4282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53404, value : 32'h706cff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53405, value : 32'hb88fd808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53406, value : 32'hf00bb500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53407, value : 32'h28741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53408, value : 32'hee60000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53409, value : 32'h740cfbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5340a, value : 32'hfb2f0886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5340b, value : 32'hc0bf4082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5340c, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5340d, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5340e, value : 32'h200ac2f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5340f, value : 32'h80f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53410, value : 32'h20292000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53411, value : 32'h206f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53412, value : 32'h100020c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53413, value : 32'h701420c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53414, value : 32'hb0698},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53415, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53416, value : 32'h8f00019a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53417, value : 32'h1600e886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53418, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53419, value : 32'he812019b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5341a, value : 32'hc420aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5341b, value : 32'h3f0811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5341c, value : 32'h20ab720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5341d, value : 32'h710c00c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5341e, value : 32'hc420ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5341f, value : 32'h10420aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53420, value : 32'h20aa5032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53421, value : 32'h50330144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53422, value : 32'h19c3266f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53423, value : 32'h70451e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53424, value : 32'h80900c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53425, value : 32'h903045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53426, value : 32'h16ef03b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53427, value : 32'hc529481},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53428, value : 32'h950002e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53429, value : 32'h41d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5342a, value : 32'h9122408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5342b, value : 32'h1e00fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5342c, value : 32'hdfe1444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5342d, value : 32'h41c30080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5342e, value : 32'h323},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5342f, value : 32'hfbef0e4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53430, value : 32'ha16d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53431, value : 32'h40c3fa4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53432, value : 32'hf4f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53433, value : 32'h902446cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53434, value : 32'hb60020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53435, value : 32'hb602d8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53436, value : 32'h41c3d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53437, value : 32'h10325},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53438, value : 32'hfbef0e26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53439, value : 32'h95424222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5343a, value : 32'h9560d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5343b, value : 32'h32641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5343c, value : 32'h15fc0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5343d, value : 32'h16009104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5343e, value : 32'h90087105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5343f, value : 32'he0a03b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53440, value : 32'h15f8fbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53441, value : 32'hdd29106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53442, value : 32'hcc20fdcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53443, value : 32'h8139620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53444, value : 32'h700c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53445, value : 32'h32741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53446, value : 32'hcce0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53447, value : 32'hcc21f98f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53448, value : 32'h8119622},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53449, value : 32'hd9650060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5344a, value : 32'hcbe700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5344b, value : 32'hb913f9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5344c, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5344d, value : 32'h1858000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5344e, value : 32'hbecb8e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5344f, value : 32'h256f00c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53450, value : 32'h42d31243},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53451, value : 32'h11408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53452, value : 32'hb8c38d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53453, value : 32'hb8149566},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53454, value : 32'h20431a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53455, value : 32'h1600aaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53456, value : 32'hc1e5031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53457, value : 32'hc3efdcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53458, value : 32'hc809fdcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53459, value : 32'h4170bbe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5345a, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5345b, value : 32'h900c0f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5345c, value : 32'h1000003c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5345d, value : 32'hf28e0113},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5345e, value : 32'h70451e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5345f, value : 32'h2889008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53460, value : 32'h200d6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53461, value : 32'h1600710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53462, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53463, value : 32'he8940019},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53464, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53465, value : 32'hd8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53466, value : 32'h5e080b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53467, value : 32'h8198d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53468, value : 32'h8f00011e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53469, value : 32'h1600e888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5346a, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5346b, value : 32'h7014019b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5346c, value : 32'hfa810b50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5346d, value : 32'hff4f0e62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5346e, value : 32'hfecf0d06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5346f, value : 32'h32d41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53470, value : 32'hd460000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53471, value : 32'h740cfbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53472, value : 32'hfe0f0daa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53473, value : 32'hfa0f08d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53474, value : 32'h742c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53475, value : 32'hfa6f0c02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53476, value : 32'h700c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53477, value : 32'hfa6f08b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53478, value : 32'hd7e712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53479, value : 32'h700c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5347a, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5347b, value : 32'hd8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5347c, value : 32'h5e080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5347d, value : 32'hb8e48d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5347e, value : 32'h1410e64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5347f, value : 32'h1a43266f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53480, value : 32'hfbef0e36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53481, value : 32'h10451e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53482, value : 32'hfb0f0fc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53483, value : 32'hfecf0bca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53484, value : 32'h1000dde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53485, value : 32'h233e0937},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53486, value : 32'h70edd933},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53487, value : 32'hd80ab914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53488, value : 32'hfbef0ce6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53489, value : 32'h1600bf8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5348a, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5348b, value : 32'h70140184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5348c, value : 32'h32120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5348d, value : 32'h30021a0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5348e, value : 32'hf9af0e7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5348f, value : 32'hd809b6e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53490, value : 32'hb600b80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53491, value : 32'h200d62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53492, value : 32'hbfed80d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53493, value : 32'h8520340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53494, value : 32'h40c3fa0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53495, value : 32'h3a980000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53496, value : 32'hff6f0d4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53497, value : 32'h780f702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53498, value : 32'h2048d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53499, value : 32'h700c0202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5349a, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5349b, value : 32'h87670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5349c, value : 32'h70ccfa6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5349d, value : 32'h81e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5349e, value : 32'h712cfa6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5349f, value : 32'hfa8f0a82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a0, value : 32'h1a00710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a1, value : 32'hb88f2003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a2, value : 32'hd1eb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a3, value : 32'h700c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a4, value : 32'hfc6f0de6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a5, value : 32'h92d710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a6, value : 32'hd80a207e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a7, value : 32'h2f241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a8, value : 32'hc660000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534a9, value : 32'h266ffbcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534aa, value : 32'h710c1a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ab, value : 32'h1a0094a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ac, value : 32'h10851e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ad, value : 32'hb88f720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ae, value : 32'hceeb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534af, value : 32'h710c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b0, value : 32'h20be094d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b1, value : 32'h1a43266f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b2, value : 32'hfaef0f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b3, value : 32'h11051e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b4, value : 32'h41c3e80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b5, value : 32'h2ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b6, value : 32'hfbef0c2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b7, value : 32'h91ad80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b8, value : 32'hd80901a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534b9, value : 32'hb88f740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ba, value : 32'h750cb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534bb, value : 32'h41c3f00e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534bc, value : 32'h2ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534bd, value : 32'hfbef0c12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534be, value : 32'h8fed80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534bf, value : 32'h700c01a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c0, value : 32'hb88f740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c1, value : 32'h720cb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c2, value : 32'hc9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c3, value : 32'hbf8e70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c4, value : 32'ha3d52104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c5, value : 32'hd92ff212},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c6, value : 32'hbeed80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c7, value : 32'hb914fbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c8, value : 32'h1a43266f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534c9, value : 32'h8d2d80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ca, value : 32'hb6e001a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534cb, value : 32'hb80e730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534cc, value : 32'hc76b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534cd, value : 32'hd8140020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ce, value : 32'ha2142144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534cf, value : 32'h832f204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d0, value : 32'h710c02e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d1, value : 32'h21be0939},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d2, value : 32'hd80ad95f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d3, value : 32'hbbab913},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d4, value : 32'h228afbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d5, value : 32'ha462001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d6, value : 32'h266ffdcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d7, value : 32'hd80b1a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d8, value : 32'h14841e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534d9, value : 32'h1a00892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534da, value : 32'h30431a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534db, value : 32'hb88fd840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534dc, value : 32'hc36b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534dd, value : 32'h760c0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534de, value : 32'h30031a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534df, value : 32'hf445262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e0, value : 32'h3003e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e1, value : 32'hfacf0ed2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e2, value : 32'h41c3e808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e3, value : 32'h2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e4, value : 32'hfbef0b76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e5, value : 32'hf015d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e6, value : 32'h2f941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e7, value : 32'hb6a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e8, value : 32'hd80afbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534e9, value : 32'h266fd880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ea, value : 32'hb6001a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534eb, value : 32'h1a0084a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ec, value : 32'hd880d80d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ed, value : 32'hb600b88f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ee, value : 32'h200bee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ef, value : 32'hd69d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f0, value : 32'h16002010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f1, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f2, value : 32'h8510164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f3, value : 32'hd80a013f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f4, value : 32'h2f141c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f5, value : 32'hb320000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f6, value : 32'h266ffbcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f7, value : 32'hcfe1a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f8, value : 32'hb6e0f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534f9, value : 32'h218a7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534fa, value : 32'hd8ff0fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534fb, value : 32'hffaf0a4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534fc, value : 32'h730c703c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534fd, value : 32'hb600b80e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534fe, value : 32'h200bae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h534ff, value : 32'h8d20d814},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53500, value : 32'h704c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53501, value : 32'hfc2f0c42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53502, value : 32'h8d20706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53503, value : 32'h714c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53504, value : 32'hfc2f0c36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53505, value : 32'hf008716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53506, value : 32'h33141c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53507, value : 32'haea0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53508, value : 32'hd80afbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53509, value : 32'h22be096b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5350a, value : 32'h41c3d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5350b, value : 32'h2fb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5350c, value : 32'hfbef0ad6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5350d, value : 32'h1010278a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5350e, value : 32'hf9cf0ca2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5350f, value : 32'h16004210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53510, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53511, value : 32'hb620163},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53512, value : 32'h712cfaaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53513, value : 32'h1a43266f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53514, value : 32'he724142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53515, value : 32'hb6e00260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53516, value : 32'hb80ad821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53517, value : 32'hca0ab600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53518, value : 32'hd825e894},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53519, value : 32'hb89f70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5351a, value : 32'h8820724e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5351b, value : 32'h7e2588db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5351c, value : 32'h13ee0e13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5351d, value : 32'hed640e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5351e, value : 32'h712cfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5351f, value : 32'hfc2f09c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53520, value : 32'h228d41e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53521, value : 32'h71ed2e3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53522, value : 32'h200b1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53523, value : 32'h92fd80e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53524, value : 32'h16002051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53525, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53526, value : 32'he8980019},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53527, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53528, value : 32'h11d8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53529, value : 32'h41c3e892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5352a, value : 32'h332},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5352b, value : 32'hfbef0a5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5352c, value : 32'hf46d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5352d, value : 32'hd8080160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5352e, value : 32'h90bf008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5352f, value : 32'h710c213f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53530, value : 32'h700cf002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53531, value : 32'h1400ec2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53532, value : 32'h213e096f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53533, value : 32'h1000704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53534, value : 32'h12242080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53535, value : 32'hb8e2370e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53536, value : 32'hf9ef0c02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53537, value : 32'h23e122ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53538, value : 32'h1fc7278a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53539, value : 32'hdfffe882},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5353a, value : 32'h117e0e4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5353b, value : 32'h41c3d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5353c, value : 32'h2fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5353d, value : 32'hfbcf0a12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5353e, value : 32'h404208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5353f, value : 32'h1a43266f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53540, value : 32'h720cb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53541, value : 32'haee4142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53542, value : 32'h42e10020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53543, value : 32'hfacf0d5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53544, value : 32'h41c3e80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53545, value : 32'h2ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53546, value : 32'hfbef09ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53547, value : 32'h730c740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53548, value : 32'had24142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53549, value : 32'h42e10020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5354a, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5354b, value : 32'hb6008110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5354c, value : 32'h200a76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5354d, value : 32'hcafd816},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5354e, value : 32'h704e2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5354f, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53550, value : 32'h90200188},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53551, value : 32'h8700103f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53552, value : 32'h700c7030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53553, value : 32'hf5ef785},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53554, value : 32'h20520000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53555, value : 32'h1a050000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53556, value : 32'h700c3002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53557, value : 32'h2a00e12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53558, value : 32'h34821a0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53559, value : 32'he807ca05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5355a, value : 32'he06700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5355b, value : 32'h1a0c02a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5355c, value : 32'h10003043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5355d, value : 32'h12242080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5355e, value : 32'hb8e2370e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5355f, value : 32'hf9ef0b5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53560, value : 32'h23e122ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53561, value : 32'h1fc7278a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53562, value : 32'hdfffe882},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53563, value : 32'h119e0e0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53564, value : 32'hfacf0cc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53565, value : 32'h41c3e808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53566, value : 32'h301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53567, value : 32'hfbef096a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53568, value : 32'hf021d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53569, value : 32'hd80a732c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5356a, value : 32'hfbef095e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5356b, value : 32'h208ab918},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5356c, value : 32'h266f0204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5356d, value : 32'hb6001a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5356e, value : 32'h4142710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5356f, value : 32'h200a36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53570, value : 32'h40c342e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53571, value : 32'h9080000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53572, value : 32'h700cb600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53573, value : 32'ha264142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53574, value : 32'h42e10020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53575, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53576, value : 32'hb6008108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53577, value : 32'h2009ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53578, value : 32'h953d818},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53579, value : 32'hd80a227e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5357a, value : 32'h30241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5357b, value : 32'h91a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5357c, value : 32'h228afbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5357d, value : 32'hae62008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5357e, value : 32'h1000f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5357f, value : 32'h4010208f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53580, value : 32'hfc6f0a86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53581, value : 32'hbfe2730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53582, value : 32'h266f700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53583, value : 32'h20ca1a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53584, value : 32'h410203e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53585, value : 32'h2200c46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53586, value : 32'h14841e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53587, value : 32'hb809d841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53588, value : 32'hca0ab600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53589, value : 32'hfeae884},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5358a, value : 32'h8d00fbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5358b, value : 32'h20097a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5358c, value : 32'hca0ad809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5358d, value : 32'hd825e828},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5358e, value : 32'hb89f70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5358f, value : 32'h8820720e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53590, value : 32'h7e2588db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53591, value : 32'h13ee0e27},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53592, value : 32'hd0240e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53593, value : 32'h712cfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53594, value : 32'h42008d20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53595, value : 32'h43e1710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53596, value : 32'hfc2f09ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53597, value : 32'h8d204250},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53598, value : 32'h4242700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53599, value : 32'hfc2f09e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5359a, value : 32'h208d43e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5359b, value : 32'h71ed2bbf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5359c, value : 32'hfbef0f9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5359d, value : 32'h16008d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5359e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5359f, value : 32'hb8e50000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a0, value : 32'hfc4209bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a1, value : 32'hfecf0baa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a2, value : 32'h20500921},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a3, value : 32'h20448d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a4, value : 32'h9150c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a5, value : 32'h80b0c10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a6, value : 32'h700c017f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a7, value : 32'h710cf002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a8, value : 32'h2c00bda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535a9, value : 32'h1000e6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535aa, value : 32'h800cba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ab, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ac, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ad, value : 32'hc03c900f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ae, value : 32'h4c41800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535af, value : 32'h160087a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b0, value : 32'hdfa700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b1, value : 32'h41c30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b2, value : 32'h335},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b3, value : 32'hfbef083a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b4, value : 32'h9a6d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b5, value : 32'h700cfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b6, value : 32'h2a00f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b7, value : 32'h700cd807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b8, value : 32'hc420ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535b9, value : 32'hf0007fff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ba, value : 32'h2800c1a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535bb, value : 32'h4308c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535bc, value : 32'h730c71ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535bd, value : 32'h900f46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535be, value : 32'h80ec028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535bf, value : 32'hb6a0ff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c0, value : 32'h900847cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c1, value : 32'h97000288},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c2, value : 32'hb3db8a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c3, value : 32'hb7001031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c4, value : 32'h900f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c5, value : 32'h40c3c298},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c6, value : 32'h3fff0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c7, value : 32'h19e8b1a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c8, value : 32'h20508004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535c9, value : 32'h40c30341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ca, value : 32'hc2249007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535cb, value : 32'h1600b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535cc, value : 32'h80007082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535cd, value : 32'h2253000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ce, value : 32'hf205817e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535cf, value : 32'h51804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d0, value : 32'hb022f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d1, value : 32'hff2f0fc2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d2, value : 32'hd81fd80d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d3, value : 32'h135c1fac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d4, value : 32'hff2f0fb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d5, value : 32'h10051e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d6, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d7, value : 32'h4308c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d8, value : 32'hff2f0fa6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535d9, value : 32'h70add81f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535da, value : 32'h900846cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535db, value : 32'h740c03e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535dc, value : 32'hff2f0f96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535dd, value : 32'h1654b6a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535de, value : 32'h206c9700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535df, value : 32'hb8810040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e0, value : 32'h10300b0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e1, value : 32'h901c1e54},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e2, value : 32'h700cc6c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e3, value : 32'h900f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e4, value : 32'hb88cc280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e5, value : 32'h40c3b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e6, value : 32'hc2249007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e7, value : 32'hb0a2b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e8, value : 32'hc6c4b1ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535e9, value : 32'h4608c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ea, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535eb, value : 32'h128000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ec, value : 32'h8203208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ed, value : 32'h2ae0e24},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ee, value : 32'hef640c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ef, value : 32'he060040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f0, value : 32'hb22fecf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f1, value : 32'hca110080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f2, value : 32'h800145cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f3, value : 32'h25164fcc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f4, value : 32'h8721000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f5, value : 32'hb0c0fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f6, value : 32'h30821211},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f7, value : 32'ha5017d56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f8, value : 32'hc326a01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535f9, value : 32'h1a11faef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535fa, value : 32'hbfe3002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535fb, value : 32'hc6c40280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535fc, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535fd, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535fe, value : 32'h41583304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h535ff, value : 32'h4310c141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53600, value : 32'h702cc08e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53601, value : 32'hf96f08fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53602, value : 32'h708eda50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53603, value : 32'h35001c34},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53604, value : 32'h35001c30},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53605, value : 32'h35001c2c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53606, value : 32'hfbef0c76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53607, value : 32'h35001c28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53608, value : 32'h21350b27},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53609, value : 32'h2353c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5360a, value : 32'h730c20c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5360b, value : 32'h21787839},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5360c, value : 32'hb8c000db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5360d, value : 32'h202fc043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5360e, value : 32'h26f004c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5360f, value : 32'h80007000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53610, value : 32'hc04410cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53611, value : 32'h700cf007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53612, value : 32'hb890706f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53613, value : 32'h4063c044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53614, value : 32'h2350c043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53615, value : 32'h21842000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53616, value : 32'hc0473004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53617, value : 32'h46d3720c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53618, value : 32'h12298000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53619, value : 32'h800047d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5361a, value : 32'hc045c14c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5361b, value : 32'h458ad825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5361c, value : 32'h718eb89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5361d, value : 32'h881b8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5361e, value : 32'h2c007905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5361f, value : 32'hb8022340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53620, value : 32'h350200f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53621, value : 32'ha040200b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53622, value : 32'h210408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53623, value : 32'hffa730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53624, value : 32'h1e00fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53625, value : 32'hc0042342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53626, value : 32'hdc278a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53627, value : 32'hc04602a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53628, value : 32'hc8094110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53629, value : 32'h7825c106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5362a, value : 32'h208916b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5362b, value : 32'h20881602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5362c, value : 32'h8b2840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5362d, value : 32'h20811601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5362e, value : 32'h1064086d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5362f, value : 32'h96540a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53630, value : 32'h2940106e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53631, value : 32'h215a0380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53632, value : 32'h2005050c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53633, value : 32'hc78e02c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53634, value : 32'h7280244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53635, value : 32'hf832005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53636, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53637, value : 32'h679f700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53638, value : 32'h80020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53639, value : 32'h30310911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5363a, value : 32'h6822100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5363b, value : 32'h821220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5363c, value : 32'h80082f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5363d, value : 32'h30300b0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5363e, value : 32'h2422079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5363f, value : 32'h2078f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53640, value : 32'hea8f0242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53641, value : 32'h271080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53642, value : 32'h9340c68e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53643, value : 32'hf009b749},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53644, value : 32'h2822840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53645, value : 32'h7a65669e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53646, value : 32'h92407e14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53647, value : 32'h7104b640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53648, value : 32'hf1cc7124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53649, value : 32'h3005140c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5364a, value : 32'hc28c4162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5364b, value : 32'h708cc38a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5364c, value : 32'hfcaf0836},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5364d, value : 32'h40c370cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5364e, value : 32'h12e48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5364f, value : 32'h21798020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53650, value : 32'h40a13002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53651, value : 32'hca24340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53652, value : 32'h4250fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53653, value : 32'h30300b73},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53654, value : 32'h1407262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53655, value : 32'hfde710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53656, value : 32'h41c1fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53657, value : 32'h800a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53658, value : 32'h38812455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53659, value : 32'hda084022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5365a, value : 32'h44c14362},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5365b, value : 32'h3c052440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5365c, value : 32'h480260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5365d, value : 32'hd9671ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5365e, value : 32'h2455fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5365f, value : 32'hda23388f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53660, value : 32'hba0a40e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53661, value : 32'hf92f0f7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53662, value : 32'hc301702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53663, value : 32'h1408d808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53664, value : 32'h41623004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53665, value : 32'h2440704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53666, value : 32'h260a3c05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53667, value : 32'h70ec0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53668, value : 32'hfbaf094e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53669, value : 32'h2455c740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5366a, value : 32'hd263880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5366b, value : 32'h702cfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5366c, value : 32'hf82700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5366d, value : 32'h41c1fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5366e, value : 32'hc00e36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5366f, value : 32'h2455f029},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53670, value : 32'h40223881},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53671, value : 32'h4362da08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53672, value : 32'h244044c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53673, value : 32'h260a3c05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53674, value : 32'h71ec0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53675, value : 32'hfb6f0d36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53676, value : 32'h388f2455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53677, value : 32'h40e2da23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53678, value : 32'hf1eba0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53679, value : 32'h702cf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5367a, value : 32'hd808c301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5367b, value : 32'h30041408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5367c, value : 32'h704c4162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5367d, value : 32'h3c052440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5367e, value : 32'h480260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5367f, value : 32'h8f270ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53680, value : 32'hc740fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53681, value : 32'h38802455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53682, value : 32'hfb6f0cc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53683, value : 32'h1601702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53684, value : 32'h16022091},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53685, value : 32'h210c2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53686, value : 32'h25ca000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53687, value : 32'h40c3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53688, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53689, value : 32'h20118800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5368a, value : 32'h2468440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5368b, value : 32'h29400021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5368c, value : 32'hc0062315},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5368d, value : 32'h5402005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5368e, value : 32'hc049700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5368f, value : 32'h2280215a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53690, value : 32'h917c048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53691, value : 32'h21003031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53692, value : 32'h10202680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53693, value : 32'h200c0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53694, value : 32'h214a000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53695, value : 32'hb0d0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53696, value : 32'h20793030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53697, value : 32'hf0042240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53698, value : 32'h22402078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53699, value : 32'h2007014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5369a, value : 32'hc2080002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5369b, value : 32'h229a7202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5369c, value : 32'h2232000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5369d, value : 32'h80000f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5369e, value : 32'heb14c44c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5369f, value : 32'h700b2b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a0, value : 32'h5c02234},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a1, value : 32'hb1772e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a2, value : 32'h922100f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a3, value : 32'hde809282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a4, value : 32'h4e924913},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a5, value : 32'ha20b17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a6, value : 32'h42104291},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a7, value : 32'hf0074628},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a8, value : 32'h70cd704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536a9, value : 32'hde80f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536aa, value : 32'h215a4210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ab, value : 32'hc08e2501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ac, value : 32'hc007603a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ad, value : 32'h40f22f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ae, value : 32'hb1080f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536af, value : 32'hc08c4058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b0, value : 32'h44020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b1, value : 32'hd0ef00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b2, value : 32'h40e1fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b3, value : 32'hc08c4708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b4, value : 32'hfbaf0d02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b5, value : 32'h44020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b6, value : 32'h4f10661e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b7, value : 32'h20024ef1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b8, value : 32'h72760480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536b9, value : 32'h20ca4608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ba, value : 32'h26ca0045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536bb, value : 32'hb411046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536bc, value : 32'h12092030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536bd, value : 32'hbb73609},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536be, value : 32'h28402071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536bf, value : 32'h47cb220b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c0, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c1, value : 32'h154b2305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c2, value : 32'h124b2305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c3, value : 32'h1f812305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c4, value : 32'h6a0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c5, value : 32'hb90261b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c6, value : 32'h3c82105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c7, value : 32'h1f812305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c8, value : 32'h680001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536c9, value : 32'hb90261b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ca, value : 32'hf0787f25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536cb, value : 32'h220b2840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536cc, value : 32'h900042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536cd, value : 32'h23050000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ce, value : 32'h7bd0154b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536cf, value : 32'h124b2305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d0, value : 32'h23057810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d1, value : 32'h11f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d2, value : 32'h61b90068},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d3, value : 32'h7f4569f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d4, value : 32'h21099720},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d5, value : 32'h230500ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d6, value : 32'h11f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d7, value : 32'h61b9006a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d8, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536d9, value : 32'h10000088},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536da, value : 32'h21091101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536db, value : 32'h23050000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536dc, value : 32'hb9021341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536dd, value : 32'hf822105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536de, value : 32'h489004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536df, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e0, value : 32'h409004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e1, value : 32'h16009240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e2, value : 32'h80007083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e3, value : 32'hb8d00ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e4, value : 32'h91200030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e5, value : 32'hb9c6bac6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e6, value : 32'h21cc72d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e7, value : 32'h5e838d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e8, value : 32'ha59000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536e9, value : 32'h4a760065},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ea, value : 32'hb2df029},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536eb, value : 32'h210520b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ec, value : 32'h28401541},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ed, value : 32'h43c32202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ee, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ef, value : 32'h21057945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f0, value : 32'h10f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f1, value : 32'h62ba0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f2, value : 32'hf812105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f3, value : 32'h630001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f4, value : 32'hf00eba02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f5, value : 32'hf822105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f6, value : 32'h190001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f7, value : 32'h7ab4b981},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f8, value : 32'hba02b985},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536f9, value : 32'h43c3b990},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536fa, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536fb, value : 32'hb2c07a65},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536fc, value : 32'hb90261b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536fd, value : 32'hf0277965},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536fe, value : 32'h621c4976},
                          '{ step_type : REG_WRITE, reg_addr : 32'h536ff, value : 32'hf705e4fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53700, value : 32'he4ff611c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53701, value : 32'h90ff78a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53702, value : 32'h228700a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53703, value : 32'h4a700fc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53704, value : 32'h2187f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53705, value : 32'h49700fc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53706, value : 32'h1f812305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53707, value : 32'h6c0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53708, value : 32'h42c361b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53709, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5370a, value : 32'hb7c0b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5370b, value : 32'hb1c07945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5370c, value : 32'h1f812305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5370d, value : 32'h6e0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5370e, value : 32'h180061b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5370f, value : 32'hb9021004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53710, value : 32'hb1007945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53711, value : 32'h41c3c009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53712, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53713, value : 32'h340320f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53714, value : 32'h2402005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53715, value : 32'h2270080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53716, value : 32'h2840b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53717, value : 32'h78452282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53718, value : 32'hb0607825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53719, value : 32'h204c7106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5371a, value : 32'h5daa280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5371b, value : 32'h5a7ffc5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5371c, value : 32'h7126ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5371d, value : 32'h20110b1d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5371e, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5371f, value : 32'hc49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53720, value : 32'h2204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53721, value : 32'h900741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53722, value : 32'hb140c0c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53723, value : 32'hb100b8a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53724, value : 32'h7704c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53725, value : 32'h3d87014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53726, value : 32'hc045ffe2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53727, value : 32'h33042480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53728, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53729, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5372a, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5372b, value : 32'hd8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5372c, value : 32'h8002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5372d, value : 32'hb8257fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5372e, value : 32'hc1a4c3e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5372f, value : 32'h70cddd37},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53730, value : 32'h1501bd9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53731, value : 32'hc0621480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53732, value : 32'h14801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53733, value : 32'h30021c09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53734, value : 32'h14801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53735, value : 32'h30021c0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53736, value : 32'h14801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53737, value : 32'h30021c0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53738, value : 32'h14801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53739, value : 32'h1501c063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5373a, value : 32'h1c0d1480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5373b, value : 32'h15013002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5373c, value : 32'h1c0e1480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5373d, value : 32'h15143002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5373e, value : 32'h1c0f1480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5373f, value : 32'hc0823002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53740, value : 32'h22141c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53741, value : 32'h60cb0002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53742, value : 32'h9fe740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53743, value : 32'h42c1fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53744, value : 32'heef71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53745, value : 32'h15019214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53746, value : 32'hc0601480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53747, value : 32'h14801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53748, value : 32'h30021c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53749, value : 32'h14801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5374a, value : 32'h30021c02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5374b, value : 32'h14801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5374c, value : 32'h30021c03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5374d, value : 32'h14801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5374e, value : 32'h8d00c061},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5374f, value : 32'h30021c05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53750, value : 32'h1c068d01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53751, value : 32'h8d023002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53752, value : 32'h1c0770ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53753, value : 32'hc0803002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53754, value : 32'h22241c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53755, value : 32'h60ab0002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53756, value : 32'h9ae740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53757, value : 32'h42a1fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53758, value : 32'hdef71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53759, value : 32'hc7c49214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5375a, value : 32'h46cbc2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5375b, value : 32'h46a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5375c, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5375d, value : 32'h8131a28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5375e, value : 32'h470802ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5375f, value : 32'h20539600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53760, value : 32'hf41180be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53761, value : 32'h950af00d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53762, value : 32'hb50ab880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53763, value : 32'h20538e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53764, value : 32'hf20780be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53765, value : 32'ha503700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53766, value : 32'ha501a502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53767, value : 32'hcd6a500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53768, value : 32'h262ff98f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53769, value : 32'h8f3c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5376a, value : 32'hc6c60004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5376b, value : 32'h20538e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5376c, value : 32'hf20780be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5376d, value : 32'ha503700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5376e, value : 32'ha501a502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5376f, value : 32'hcb6a500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53770, value : 32'hc6c6f98f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53771, value : 32'h46a8c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53772, value : 32'h40704788},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53773, value : 32'h9d64548},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53774, value : 32'h4130fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53775, value : 32'h2281215f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53776, value : 32'h25cae589},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53777, value : 32'h60381221},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53778, value : 32'h229f7a0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53779, value : 32'h2200000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5377a, value : 32'h20000400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5377b, value : 32'h80000f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5377c, value : 32'h8960c44c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5377d, value : 32'hb1d710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5377e, value : 32'h78b800f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5377f, value : 32'h700b3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53780, value : 32'hb5178cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53781, value : 32'h78cb00b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53782, value : 32'h78cbeb83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53783, value : 32'hc6caf22c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53784, value : 32'hf3ff78cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53785, value : 32'h2180205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53786, value : 32'h40c3621a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53787, value : 32'hc14c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53788, value : 32'h9340621b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53789, value : 32'h78429301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5378a, value : 32'h93027c10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5378b, value : 32'h7a504f12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5378c, value : 32'h10850c1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5378d, value : 32'hb300b3e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5378e, value : 32'hf3ebf009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5378f, value : 32'h2180205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53790, value : 32'h70c36058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53791, value : 32'hc14e8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53792, value : 32'h1900b0e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53793, value : 32'hc6ca0083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53794, value : 32'h205ff5df},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53795, value : 32'h19002180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53796, value : 32'h605800c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53797, value : 32'h800070c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53798, value : 32'hf00ac150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53799, value : 32'h2180205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5379a, value : 32'h431900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5379b, value : 32'h70c36058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5379c, value : 32'hc14c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5379d, value : 32'hc6cab0e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5379e, value : 32'hc1a6c3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5379f, value : 32'h44104530},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a0, value : 32'hf2b27014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a1, value : 32'h230a70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a2, value : 32'h25142500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a3, value : 32'h244023d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a4, value : 32'h21143511},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a5, value : 32'h120023d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a6, value : 32'h20532100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a7, value : 32'h19010141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a8, value : 32'h702c2042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537a9, value : 32'h1900b826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537aa, value : 32'h8e62002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ab, value : 32'h4022feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ac, value : 32'h21001204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ad, value : 32'h34102440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ae, value : 32'h23d02014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537af, value : 32'h1412053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b0, value : 32'h20421801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b1, value : 32'hb826702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b2, value : 32'h20021800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b3, value : 32'hfeaf08c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b4, value : 32'h40224002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b5, value : 32'hdae4102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b6, value : 32'h724c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b7, value : 32'h2100120a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b8, value : 32'h7ef4c683},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537b9, value : 32'h1412053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ba, value : 32'h712cae21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537bb, value : 32'hae00b826},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537bc, value : 32'hfeaf089e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537bd, value : 32'h120e40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537be, value : 32'hc5822100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537bf, value : 32'h20537df4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c0, value : 32'had210141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c1, value : 32'hb826712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c2, value : 32'h886ad00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c3, value : 32'h40a1feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c4, value : 32'h41a140c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c5, value : 32'h600d6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c6, value : 32'h1101724c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c7, value : 32'he0c02080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c8, value : 32'hd940f704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537c9, value : 32'hf0044910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ca, value : 32'h3f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537cb, value : 32'h31812440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537cc, value : 32'ha90061f9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537cd, value : 32'h20801001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ce, value : 32'hf705e0c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537cf, value : 32'h4910d940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d0, value : 32'h2080f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d1, value : 32'hc181003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d2, value : 32'ha90061f9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d3, value : 32'he0c08e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d4, value : 32'hd940f704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d5, value : 32'hf0044910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d6, value : 32'h3f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d7, value : 32'h30812440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d8, value : 32'ha90061f9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537d9, value : 32'he0c08d01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537da, value : 32'hd940f704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537db, value : 32'hf0044910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537dc, value : 32'h3f2080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537dd, value : 32'h63f9c380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537de, value : 32'h238d71e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537df, value : 32'ha900227e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e0, value : 32'h7500240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e1, value : 32'h708d70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e2, value : 32'h704c706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e3, value : 32'h54020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e4, value : 32'h30802440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e5, value : 32'h22086088},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e6, value : 32'h13010001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e7, value : 32'h21080480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e8, value : 32'h24400002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537e9, value : 32'h60883180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ea, value : 32'h10012308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537eb, value : 32'h6088c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ec, value : 32'h21087185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ed, value : 32'h270a000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ee, value : 32'hc3830540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ef, value : 32'h32042440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f0, value : 32'h35052440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f1, value : 32'h34062440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f2, value : 32'h24147bb4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f3, value : 32'h25140344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f4, value : 32'h26140345},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f5, value : 32'h78af0346},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f6, value : 32'hfa2f0d36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f7, value : 32'h71a54161},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f8, value : 32'h95040ddb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537f9, value : 32'h78e0c7d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537fa, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537fb, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537fc, value : 32'h1c453b08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537fd, value : 32'h41183058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537fe, value : 32'h36001445},
                          '{ step_type : REG_WRITE, reg_addr : 32'h537ff, value : 32'h30981c46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53800, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53801, value : 32'h829122c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53802, value : 32'h1c470070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53803, value : 32'h144530d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53804, value : 32'he89f3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53805, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53806, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53807, value : 32'hc02078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53808, value : 32'h9b1200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53809, value : 32'hc0407104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5380a, value : 32'hf0118a01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5380b, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5380c, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5380d, value : 32'h412078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5380e, value : 32'h9b1202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5380f, value : 32'h7314c140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53810, value : 32'h20cac000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53811, value : 32'hc04000a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53812, value : 32'h1c438a03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53813, value : 32'hc3003018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53814, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53815, value : 32'h200ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53816, value : 32'hfb6f0eae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53817, value : 32'h70374223},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53818, value : 32'h2102f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53819, value : 32'h216fd920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5381a, value : 32'h89000bc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5381b, value : 32'h1a1e780a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5381c, value : 32'h8901301c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5381d, value : 32'h1a1f780a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5381e, value : 32'hc000301c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5381f, value : 32'h5327014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53820, value : 32'h70ee0021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53821, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53822, value : 32'h231f0a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53823, value : 32'h24003000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53824, value : 32'h3f98},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53825, value : 32'h24400124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53826, value : 32'h20803116},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53827, value : 32'h26803084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53828, value : 32'h702e2084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53829, value : 32'h800070c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5382a, value : 32'h1c441a44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5382b, value : 32'h1c483018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5382c, value : 32'h248a3018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5382d, value : 32'hc0817001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5382e, value : 32'hfc7218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5382f, value : 32'h34421a0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53830, value : 32'h14020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53831, value : 32'h1804b021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53832, value : 32'hd9ff0015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53833, value : 32'h7001248a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53834, value : 32'hfc7228a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53835, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53836, value : 32'h1240000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53837, value : 32'h27c31e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53838, value : 32'h35dc1c82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53839, value : 32'h305c1c84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5383a, value : 32'h14020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5383b, value : 32'h1804b041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5383c, value : 32'h456b0015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5383d, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5383e, value : 32'h2240000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5383f, value : 32'h37c31800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53840, value : 32'h51800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53841, value : 32'h1443b022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53842, value : 32'h8db3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53843, value : 32'hc0810364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53844, value : 32'h36001446},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53845, value : 32'ha0e79af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53846, value : 32'h1a0c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53847, value : 32'h45103358},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53848, value : 32'hdb9700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53849, value : 32'h251a240e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5384a, value : 32'h1f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5384b, value : 32'h211a0a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5384c, value : 32'h2f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5384d, value : 32'h1a0d28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5384e, value : 32'h661e3418},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5384f, value : 32'h209a4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53850, value : 32'h60d80184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53851, value : 32'h800070c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53852, value : 32'he661a44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53853, value : 32'h44100260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53854, value : 32'hf4f07014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53855, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53856, value : 32'h200c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53857, value : 32'hdaa42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53858, value : 32'h4302fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53859, value : 32'hfbe4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5385a, value : 32'h41a1fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5385b, value : 32'h24404210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5385c, value : 32'he8863113},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5385d, value : 32'h3f932400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5385e, value : 32'h1240000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5385f, value : 32'h2400d52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53860, value : 32'h42c3702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53861, value : 32'h1b468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53862, value : 32'ha0be812},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53863, value : 32'hc0812030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53864, value : 32'h2400f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53865, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53866, value : 32'h10820124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53867, value : 32'h40020701},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53868, value : 32'h184209a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53869, value : 32'h605860d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5386a, value : 32'h48319001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5386b, value : 32'h209a4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5386c, value : 32'h60d80184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5386d, value : 32'h20300a0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5386e, value : 32'h1600604a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5386f, value : 32'hf0042080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53870, value : 32'h30801000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53871, value : 32'h242f4a13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53872, value : 32'h40620046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53873, value : 32'ha4e4182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53874, value : 32'h4262faaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53875, value : 32'hf4ae7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53876, value : 32'h84b7106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53877, value : 32'h71a5a294},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53878, value : 32'hd06f193},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53879, value : 32'h41230060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5387a, value : 32'h704e7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5387b, value : 32'h2400f4a3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5387c, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5387d, value : 32'hcf20124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5387e, value : 32'h41230060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5387f, value : 32'hf49b7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53880, value : 32'h20821600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53881, value : 32'hc845cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53882, value : 32'h14840002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53883, value : 32'h740c3703},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53884, value : 32'hfb6f0cf6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53885, value : 32'h100041a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53886, value : 32'h254f3082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53887, value : 32'h24341401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53888, value : 32'h3f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53889, value : 32'hce20228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5388a, value : 32'h740cfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5388b, value : 32'h36001443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5388c, value : 32'h6e5080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5388d, value : 32'h1448714e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5388e, value : 32'hf07d3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5388f, value : 32'h360e1444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53890, value : 32'h1446476b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53891, value : 32'h79ef3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53892, value : 32'h12008da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53893, value : 32'h33d81a0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53894, value : 32'h2600c7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53895, value : 32'h45084410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53896, value : 32'heca4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53897, value : 32'h41e1fd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53898, value : 32'he808ed05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53899, value : 32'h208d1600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5389a, value : 32'he807f00d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5389b, value : 32'hf009c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5389c, value : 32'h308d1000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5389d, value : 32'h2400f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5389e, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5389f, value : 32'h10820124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a0, value : 32'h700e070d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a1, value : 32'hc6743d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a2, value : 32'h740c242e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a3, value : 32'hca41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a4, value : 32'h42e10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a5, value : 32'hc724302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a6, value : 32'h1a0dfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a7, value : 32'hc323418},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a8, value : 32'he8070240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538a9, value : 32'h88e4062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538aa, value : 32'h41a1fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ab, value : 32'h4062f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ac, value : 32'hfc6f0fa6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ad, value : 32'he8be41a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ae, value : 32'h84208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538af, value : 32'hcb41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b0, value : 32'h23320004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b1, value : 32'h740c2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b2, value : 32'h43e14222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b3, value : 32'hfb6f0c3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b4, value : 32'h400240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b5, value : 32'he80bca06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b6, value : 32'h36021445},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b7, value : 32'h14474062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b8, value : 32'h41233604},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538b9, value : 32'h3200b96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ba, value : 32'h71064322},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538bb, value : 32'ha2b4089b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538bc, value : 32'h21842380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538bd, value : 32'h2400bda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538be, value : 32'h1f82271a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538bf, value : 32'ha3c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c0, value : 32'h2f81211a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c1, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c2, value : 32'h40c37014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c3, value : 32'h1b468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c4, value : 32'hf2056159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c5, value : 32'ha8a06038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c6, value : 32'h6038f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c7, value : 32'h2695b0a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c8, value : 32'h144313ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538c9, value : 32'h77103600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ca, value : 32'hffe5071a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538cb, value : 32'hf18571e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538cc, value : 32'h7056704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538cd, value : 32'h210278},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ce, value : 32'h14447126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538cf, value : 32'h21963601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d0, value : 32'h1c440794},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d1, value : 32'hc1003058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d2, value : 32'ha040210c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d3, value : 32'hffc50562},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d4, value : 32'h25f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d5, value : 32'hb99f70ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d6, value : 32'h780a8900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d7, value : 32'h301c1a1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d8, value : 32'h780a8901},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538d9, value : 32'h301c1a1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538da, value : 32'h36001447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538db, value : 32'h936e806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538dc, value : 32'h70aefb8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538dd, value : 32'h71aee802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538de, value : 32'h44d3c781},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538df, value : 32'h1a448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e0, value : 32'h10842780},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e1, value : 32'h36001443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e2, value : 32'hb000230c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e3, value : 32'h2d0222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e4, value : 32'h144670ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e5, value : 32'h212f3600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e6, value : 32'hf8a06c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e7, value : 32'h1a0c00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e8, value : 32'h700e36d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538e9, value : 32'h30181c44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ea, value : 32'h36001444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538eb, value : 32'h84002011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ec, value : 32'h24c0270a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ed, value : 32'h248af2f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ee, value : 32'hc0817001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ef, value : 32'hfc7218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f0, value : 32'h1a0d702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f1, value : 32'h20a83418},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f2, value : 32'hb0210180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f3, value : 32'h151804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f4, value : 32'h1f00d8ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f5, value : 32'h1c8417c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f6, value : 32'hc000301c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f7, value : 32'h3008bd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f8, value : 32'h301d1c82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538f9, value : 32'h46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538fa, value : 32'h704e28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538fb, value : 32'h3380202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538fc, value : 32'h34421a0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538fd, value : 32'h211a45aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538fe, value : 32'h2e412380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h538ff, value : 32'h251f1096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53900, value : 32'h1a0e1601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53901, value : 32'h231a3358},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53902, value : 32'h61193596},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53903, value : 32'h209a4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53904, value : 32'h71c20184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53905, value : 32'h702c6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53906, value : 32'h600ace},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53907, value : 32'h47107082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53908, value : 32'hf4b87014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53909, value : 32'h71ad70b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5390a, value : 32'h7126f3e7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5390b, value : 32'h9c5c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5390c, value : 32'h70ada004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5390d, value : 32'h33421a0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5390e, value : 32'h2540210a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5390f, value : 32'h2600a92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53910, value : 32'h34581a0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53911, value : 32'h1382251a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53912, value : 32'h211f7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53913, value : 32'h43c32601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53914, value : 32'h1b468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53915, value : 32'h6159700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53916, value : 32'h229a4202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53917, value : 32'h71c20184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53918, value : 32'hf207623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53919, value : 32'h90216358},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5391a, value : 32'h37001484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5391b, value : 32'h22004910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5391c, value : 32'h626b0501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5391d, value : 32'h242f8f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5391e, value : 32'h7b420006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5391f, value : 32'hf9ec081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53920, value : 32'hc281fa6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53921, value : 32'h70144710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53922, value : 32'h7036f484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53923, value : 32'hf3d8712e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53924, value : 32'hc00071a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53925, value : 32'h90040da1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53926, value : 32'h740cd9bb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53927, value : 32'hfb6f0a6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53928, value : 32'h8f40b910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53929, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5392a, value : 32'h200bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5392b, value : 32'hfb6f0a5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5392c, value : 32'h37031484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5392d, value : 32'ha32c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5392e, value : 32'h702c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5392f, value : 32'h8d54710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53930, value : 32'h704e0031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53931, value : 32'h740c8f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53932, value : 32'hbd41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53933, value : 32'ha3a0002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53934, value : 32'h1484fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53935, value : 32'hd95f3703},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53936, value : 32'ha2e740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53937, value : 32'hb911fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53938, value : 32'h8adc000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53939, value : 32'h714e0030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5393a, value : 32'h220a702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5393b, value : 32'h1a0d2540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5393c, value : 32'h40c33442},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5393d, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5393e, value : 32'h211a791b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5393f, value : 32'h221f2002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53940, value : 32'hb8222041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53941, value : 32'h300d231a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53942, value : 32'h209a4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53943, value : 32'h61590184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53944, value : 32'h60b8653d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53945, value : 32'hf8e2000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53946, value : 32'h1a448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53947, value : 32'h26009b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53948, value : 32'h34981a0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53949, value : 32'h8f20e806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5394a, value : 32'hfc6f0e0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5394b, value : 32'hf00740c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5394c, value : 32'h37011484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5394d, value : 32'hfc6f0d22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5394e, value : 32'h471040c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5394f, value : 32'h4002e8a6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53950, value : 32'hbf41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53951, value : 32'h209a0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53952, value : 32'h42220184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53953, value : 32'h240a4363},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53954, value : 32'h60b80400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53955, value : 32'hf852032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53956, value : 32'h1b468000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53957, value : 32'hfb6f09aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53958, value : 32'hca06740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53959, value : 32'h1445e80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5395a, value : 32'h40c13602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5395b, value : 32'h36041447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5395c, value : 32'h90a702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5395d, value : 32'h43220320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5395e, value : 32'h714e7056},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5395f, value : 32'h7126f3bb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53960, value : 32'h96bc000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53961, value : 32'hf004a004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53962, value : 32'hf004704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53963, value : 32'h24c0270a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53964, value : 32'h20100a1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53965, value : 32'h204c7106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53966, value : 32'h610a280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53967, value : 32'h230affe5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53968, value : 32'h716725c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53969, value : 32'hffef05e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5396a, value : 32'h25c0230a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5396b, value : 32'h202f4710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5396c, value : 32'h248005c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5396d, value : 32'h14043b08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5396e, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5396f, value : 32'h1600c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53970, value : 32'h8000708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53971, value : 32'h40500008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53972, value : 32'hcd64130},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53973, value : 32'h4608f96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53974, value : 32'hd907706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53975, value : 32'hda284768},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53976, value : 32'h708cbf8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53977, value : 32'h70ac40e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53978, value : 32'hf9af0d02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53979, value : 32'hfaa70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5397a, value : 32'h700cf98f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5397b, value : 32'hda08d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5397c, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5397d, value : 32'hcee70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5397e, value : 32'h70ccf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5397f, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53980, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53981, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53982, value : 32'hf9af0cda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53983, value : 32'h6f1670cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53984, value : 32'h704c752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53985, value : 32'h4238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53986, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53987, value : 32'hf9af0cc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53988, value : 32'h257870cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53989, value : 32'h781b1080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5398a, value : 32'h20300845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5398b, value : 32'hd92b68a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5398c, value : 32'h10040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5398d, value : 32'h42a1000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5398e, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5398f, value : 32'h70cc45c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53990, value : 32'hf9af0ca2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53991, value : 32'h2f404010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53992, value : 32'hd92b1240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53993, value : 32'h706c42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53994, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53995, value : 32'hf9af0c8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53996, value : 32'h440260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53997, value : 32'hd92b4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53998, value : 32'h706c42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53999, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5399a, value : 32'hf00b70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5399b, value : 32'h12402f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5399c, value : 32'h42a1d92b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5399d, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5399e, value : 32'h260a45c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5399f, value : 32'hc660440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a0, value : 32'h700cf98f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a1, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a2, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a3, value : 32'hc5670ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a4, value : 32'h70ccf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a5, value : 32'hf98f0ee2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a6, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a7, value : 32'h706cda30},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a8, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539a9, value : 32'hf9af0c3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539aa, value : 32'hc6ca70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ab, value : 32'h1600c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ac, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ad, value : 32'h83f0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ae, value : 32'h45cb001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539af, value : 32'hc148900b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b0, value : 32'h10451d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b1, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b2, value : 32'h12ff0203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b3, value : 32'h8a008481},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b4, value : 32'hb810b918},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b5, value : 32'h12ff7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b6, value : 32'hb9088081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b7, value : 32'h12fe7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b8, value : 32'h20058080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539b9, value : 32'h8868040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ba, value : 32'h20cafeef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539bb, value : 32'h1d0002a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539bc, value : 32'hc6c21005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539bd, value : 32'h1600c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539be, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539bf, value : 32'h45cb001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c0, value : 32'hc40c900f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c1, value : 32'h510821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c2, value : 32'h900f40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c3, value : 32'h1d00c1e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c4, value : 32'h1d001045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c5, value : 32'h18001005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c6, value : 32'h18000185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c7, value : 32'hfea0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c8, value : 32'hd820feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539c9, value : 32'hfe2750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ca, value : 32'h1d00feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539cb, value : 32'hd8201045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539cc, value : 32'h900f46cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539cd, value : 32'hfd2c1e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ce, value : 32'h1e00feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539cf, value : 32'h1d001185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d0, value : 32'h1e001005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d1, value : 32'hc6c41005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d2, value : 32'hd841c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d3, value : 32'h900845cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d4, value : 32'hb50001e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d5, value : 32'hfeaf0fb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d6, value : 32'hd840750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d7, value : 32'hc6c2b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d8, value : 32'hc1a4c3f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539d9, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539da, value : 32'h15020150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539db, value : 32'hd93d1500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539dc, value : 32'hb2004283},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539dd, value : 32'h1502b911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539de, value : 32'hb2011500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539df, value : 32'h15001502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e0, value : 32'h1502b202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e1, value : 32'hb2031500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e2, value : 32'h15001502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e3, value : 32'h9500b204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e4, value : 32'h9501b205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e5, value : 32'h9502b206},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e6, value : 32'hf6eb207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e7, value : 32'h740cfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e8, value : 32'h908015d7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539e9, value : 32'h1210e804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ea, value : 32'hf0043092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539eb, value : 32'h3092120f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ec, value : 32'h710c702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ed, value : 32'he80872ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ee, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ef, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f0, value : 32'hf045e888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f1, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f2, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f3, value : 32'h100887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f4, value : 32'hc08070ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f5, value : 32'h78b5700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f6, value : 32'h70ed728e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f7, value : 32'h44020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f8, value : 32'h2005781b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539f9, value : 32'h40f93},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539fa, value : 32'ha571000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539fb, value : 32'h250a2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539fc, value : 32'h70cd2480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539fd, value : 32'h1b00255a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539fe, value : 32'h1f852632},
                          '{ step_type : REG_WRITE, reg_addr : 32'h539ff, value : 32'h4788000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a00, value : 32'h430242a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a01, value : 32'h440240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a02, value : 32'h201478d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a03, value : 32'h70020440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a04, value : 32'hf812000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a05, value : 32'h12308000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a06, value : 32'h706278ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a07, value : 32'hb89cb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a08, value : 32'h8000b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a09, value : 32'h262fa900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a0a, value : 32'h41c30007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a0b, value : 32'h5007b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a0c, value : 32'hfb2f0ed6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a0d, value : 32'h71c5740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a0e, value : 32'h27bf258d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a0f, value : 32'h248d71e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a10, value : 32'h710e25ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a11, value : 32'hd8f71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a12, value : 32'h700c9114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a13, value : 32'h2d7e268d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a14, value : 32'hc7d4712e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a15, value : 32'h4350c2f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a16, value : 32'h8854630},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a17, value : 32'h44100030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a18, value : 32'h20002678},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a19, value : 32'h220a70d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a1a, value : 32'h781b24c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a1b, value : 32'h202222ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a1c, value : 32'h70ae68e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a1d, value : 32'h250d255a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a1e, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a1f, value : 32'h652012e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a20, value : 32'hb89cb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a21, value : 32'hb53b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a22, value : 32'h10002030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a23, value : 32'h653d0118},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a24, value : 32'h8d29702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a25, value : 32'h20008d0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a26, value : 32'h40100497},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a27, value : 32'h44a222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a28, value : 32'h72624628},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a29, value : 32'hc264003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a2a, value : 32'h702cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a2b, value : 32'h412044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a2c, value : 32'h10400e17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a2d, value : 32'h20300e11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a2e, value : 32'h20402042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a2f, value : 32'h20402040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a30, value : 32'hf003ad0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a31, value : 32'h7126ad0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a32, value : 32'ha4e409d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a33, value : 32'h23d02000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a34, value : 32'h15c21d0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a35, value : 32'h248dad29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a36, value : 32'h71a6243f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a37, value : 32'h78e0c6d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a38, value : 32'h47cbc2ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a39, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a3a, value : 32'h42508fa0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a3b, value : 32'h1090251f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a3c, value : 32'h70911600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a3d, value : 32'h48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a3e, value : 32'h46084330},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a3f, value : 32'h20d12153},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a40, value : 32'h8a58f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a41, value : 32'he390344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a42, value : 32'ha99161f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a43, value : 32'h2d402030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a44, value : 32'h6e321380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a45, value : 32'h704c7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a46, value : 32'h408202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a47, value : 32'h20032314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a48, value : 32'hb80a784f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a49, value : 32'h78257144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a4a, value : 32'hb89cb892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a4b, value : 32'h9000b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a4c, value : 32'h784fb300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a4d, value : 32'h84a408e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a4e, value : 32'hf0347106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a4f, value : 32'h7e06c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a50, value : 32'h1f802604},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a51, value : 32'hfffe0fff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a52, value : 32'hfeff70c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a53, value : 32'h2843fff0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a54, value : 32'hf2118100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a55, value : 32'hd00823},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a56, value : 32'h900817},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a57, value : 32'h71081f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a58, value : 32'hfc240c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a59, value : 32'h41a1fd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a5a, value : 32'h710c7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a5b, value : 32'h720cf408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a5c, value : 32'h700cf006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a5d, value : 32'h730cf004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a5e, value : 32'h740cf002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a5f, value : 32'h2b01215f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a60, value : 32'h8f037915},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a61, value : 32'h340203c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a62, value : 32'h26447914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a63, value : 32'h60381040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a64, value : 32'h882660f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a65, value : 32'h408202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a66, value : 32'h20002314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a67, value : 32'hb0207106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a68, value : 32'hf1b071a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a69, value : 32'h78e0c6ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a6a, value : 32'h4410c2f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a6b, value : 32'h3952840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a6c, value : 32'h1600785b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a6d, value : 32'h80007096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a6e, value : 32'h2044008e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a6f, value : 32'hd8e40182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a70, value : 32'h2c407859},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a71, value : 32'hb8c12318},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a72, value : 32'h2f8e2505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a73, value : 32'h1c89004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a74, value : 32'hf112054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a75, value : 32'h40f2040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a76, value : 32'h1972140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a77, value : 32'h704e706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a78, value : 32'h700e70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a79, value : 32'h26012205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a7a, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a7b, value : 32'ha07e2653},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a7c, value : 32'h900441c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a7d, value : 32'hf20d0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a7e, value : 32'hb80278e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a7f, value : 32'h90007825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a80, value : 32'h1c120ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a81, value : 32'hb8647314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a82, value : 32'h2d20ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a83, value : 32'h2005f00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a84, value : 32'hb8020440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a85, value : 32'h218a7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a86, value : 32'h90000fbf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a87, value : 32'h770cb8e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a88, value : 32'h4120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a89, value : 32'h20022700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a8a, value : 32'he810ca07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a8b, value : 32'h2310811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a8c, value : 32'h37011222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a8d, value : 32'hf800915},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a8e, value : 32'h68150000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a8f, value : 32'h2510811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a90, value : 32'hf81090d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a91, value : 32'h71960000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a92, value : 32'hf003ba86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a93, value : 32'hd808ba87},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a94, value : 32'hfeaf0cb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a95, value : 32'h2505b640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a96, value : 32'h225624c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a97, value : 32'h20052812},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a98, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a99, value : 32'h900001cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a9a, value : 32'h20102380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a9b, value : 32'h2800b8c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a9c, value : 32'h71060400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a9d, value : 32'ha2740871},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a9e, value : 32'h78b07d05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53a9f, value : 32'hd7e4182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa0, value : 32'h1e00fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa1, value : 32'h780f1005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa2, value : 32'h78e0c6d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa3, value : 32'h2840c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa4, value : 32'h4708038e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa5, value : 32'h2605d889},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa6, value : 32'h90041f8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa7, value : 32'hb50001c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa8, value : 32'hfeaf0c66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aa9, value : 32'h244ad808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aaa, value : 32'h708d7240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aab, value : 32'h702c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aac, value : 32'h20a8706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aad, value : 32'h26050400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aae, value : 32'h22801080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aaf, value : 32'h20050010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab0, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab1, value : 32'h900001cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab2, value : 32'h7838b8c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab3, value : 32'h7b057124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab4, value : 32'h41e17870},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab5, value : 32'hfb2f0d26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab6, value : 32'h780fb580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab7, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab8, value : 32'h14422aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ab9, value : 32'h10421aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aba, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53abb, value : 32'ha04104b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53abc, value : 32'ha0207fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53abd, value : 32'h45cbc0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53abe, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53abf, value : 32'h46008d60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac0, value : 32'ha1b718d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac1, value : 32'h700c00b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac2, value : 32'h241235f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac3, value : 32'h710a13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac4, value : 32'he108de08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac5, value : 32'hd808dc09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac6, value : 32'h4160f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac7, value : 32'h150170cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac8, value : 32'h4e12108b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ac9, value : 32'h492240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aca, value : 32'hb377d6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53acb, value : 32'he2f1344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53acc, value : 32'hbd0e1024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53acd, value : 32'h7240240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ace, value : 32'h20a84008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53acf, value : 32'h7a2f0440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad0, value : 32'h26146199},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad1, value : 32'h2840008f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad2, value : 32'h7aa51282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad3, value : 32'h22057105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad4, value : 32'h90040f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad5, value : 32'h924001d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad6, value : 32'h7164b740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad7, value : 32'hc4c6f1e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad8, value : 32'h40c3c5e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ad9, value : 32'h4988000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ada, value : 32'he9ae8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53adb, value : 32'h431800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53adc, value : 32'he82aca00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53add, value : 32'h70ad712d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ade, value : 32'h800144cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53adf, value : 32'h2d404fa8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae0, value : 32'h244a1381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae1, value : 32'h42817240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae2, value : 32'h706d700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae3, value : 32'h5c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae4, value : 32'h2002105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae5, value : 32'h20057405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae6, value : 32'h90040f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae7, value : 32'h8a000200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae8, value : 32'h2900b300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ae9, value : 32'h120112c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aea, value : 32'h71650480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aeb, value : 32'h7825b80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aec, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aed, value : 32'h2f89004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aee, value : 32'h71a5b060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aef, value : 32'hdc3ca00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af0, value : 32'he4099024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af1, value : 32'h78e0c4c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af2, value : 32'hdc25c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af3, value : 32'h43c3bc9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af4, value : 32'h122c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af5, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af6, value : 32'h90070f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af7, value : 32'hcc24c408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af8, value : 32'h8c00b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53af9, value : 32'h8b01e818},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53afa, value : 32'h82d8b20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53afb, value : 32'h78220064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53afc, value : 32'h240a7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53afd, value : 32'h20a87000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53afe, value : 32'h40c30400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53aff, value : 32'h49c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b00, value : 32'h4220f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b01, value : 32'h3802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b02, value : 32'h20057124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b03, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b04, value : 32'hb040028c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b05, value : 32'h70148c1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b06, value : 32'h8b037ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b07, value : 32'h72108b42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b08, value : 32'h7cd20e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b09, value : 32'h71047842},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b0a, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b0b, value : 32'h3c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b0c, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b0d, value : 32'h20f4049c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b0e, value : 32'h2a400081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b0f, value : 32'h71440380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b10, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b11, value : 32'h28c9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b12, value : 32'h7ee0b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b13, value : 32'h21326038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b14, value : 32'h80000f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b15, value : 32'ha8401888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b16, value : 32'hf822132},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b17, value : 32'h18d38000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b18, value : 32'h82184b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b19, value : 32'hf822132},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b1a, value : 32'h191e8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b1b, value : 32'h821896},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b1c, value : 32'hf812132},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b1d, value : 32'h19698000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b1e, value : 32'h18e17fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b1f, value : 32'h78e00042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b20, value : 32'h4748c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b21, value : 32'h851101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b22, value : 32'h46288861},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b23, value : 32'h841100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b24, value : 32'h88404508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b25, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b26, value : 32'h500d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b27, value : 32'hfb2f0a6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b28, value : 32'h8e0046e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b29, value : 32'h71108d20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b2a, value : 32'hf7c7f233},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b2b, value : 32'h3e50915},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b2c, value : 32'had006909},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b2d, value : 32'h835f00f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b2e, value : 32'h770403c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b2f, value : 32'hf01fae00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b30, value : 32'hf1349f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b31, value : 32'had001070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b32, value : 32'h10900f1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b33, value : 32'h10c01501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b34, value : 32'h8d01f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b35, value : 32'h8002054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b36, value : 32'h262fad01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b37, value : 32'h32f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b38, value : 32'hd87f0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b39, value : 32'hf015ad01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b3a, value : 32'hf1378e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b3b, value : 32'hae001070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b3c, value : 32'h10900f1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b3d, value : 32'h10c01601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b3e, value : 32'h8e01f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b3f, value : 32'h8002054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b40, value : 32'h262fae01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b41, value : 32'haf005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b42, value : 32'hd87f0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b43, value : 32'h8e60ae01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b44, value : 32'hd541c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b45, value : 32'h8d400003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b46, value : 32'h8ce44e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b47, value : 32'h2238f8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b48, value : 32'hc6c600c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b49, value : 32'hd9c5c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b4a, value : 32'h9ded80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b4b, value : 32'hb912fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b4c, value : 32'hfeaf09d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b4d, value : 32'ha52d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b4e, value : 32'h41c3f9cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b4f, value : 32'h68008001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b50, value : 32'hfa2f0d36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b51, value : 32'h43206f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b52, value : 32'h41c3e887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b53, value : 32'h315},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b54, value : 32'hfb2f09b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b55, value : 32'hc12d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b56, value : 32'h4200fc4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b57, value : 32'h41c34320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b58, value : 32'h10316},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b59, value : 32'hfb2f09a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b5a, value : 32'ha1ed80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b5b, value : 32'h46cbf9cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b5c, value : 32'h32740000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b5d, value : 32'h45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b5e, value : 32'he37332c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b5f, value : 32'hd80a1365},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b60, value : 32'h31741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b61, value : 32'h9820001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b62, value : 32'h42a1fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b63, value : 32'hda2700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b64, value : 32'h41a1fa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b65, value : 32'h4608d963},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b66, value : 32'h96eb913},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b67, value : 32'hd80afb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b68, value : 32'h40a1d941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b69, value : 32'hfa2f0cd2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b6a, value : 32'h60ddb90a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b6b, value : 32'h41c3f018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b6c, value : 32'h10319},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b6d, value : 32'hfb2f0952},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b6e, value : 32'h700c42c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b6f, value : 32'hfa2f0cba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b70, value : 32'h450841c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b71, value : 32'h31a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b72, value : 32'h93e0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b73, value : 32'hd80afb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b74, value : 32'h40c1d941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b75, value : 32'hfa2f0d5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b76, value : 32'h651db90a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b77, value : 32'h41c3ed87},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b78, value : 32'h31b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b79, value : 32'hfb2f0922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b7a, value : 32'hb7ed80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b7b, value : 32'h45cbfc4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b7c, value : 32'h4508000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b7d, value : 32'h223d8540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b7e, value : 32'h85410003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b7f, value : 32'h40223d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b80, value : 32'h20ca7150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b81, value : 32'he88600c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b82, value : 32'hfc4f0b5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b83, value : 32'ha500a521},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b84, value : 32'hfc4f0b56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b85, value : 32'h43204200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b86, value : 32'h31c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b87, value : 32'h8ea0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b88, value : 32'hd80afb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b89, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b8a, value : 32'h48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b8b, value : 32'h15e082f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b8c, value : 32'h85208501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b8d, value : 32'h213c7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b8e, value : 32'h10f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b8f, value : 32'h79c0f42c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b90, value : 32'h41c3e98d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b91, value : 32'h31d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b92, value : 32'hfb2f08be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b93, value : 32'h41c3d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b94, value : 32'h31e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b95, value : 32'hf8af0f92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b96, value : 32'hc6c4700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b97, value : 32'h4010c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b98, value : 32'hd86d80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b99, value : 32'hd90ffa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b9a, value : 32'hc2ad80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b9b, value : 32'h712cf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b9c, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b9d, value : 32'h8ea0122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b9e, value : 32'h1280255f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53b9f, value : 32'hf8f2000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba0, value : 32'h4e048001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba1, value : 32'h85f8e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba2, value : 32'h40c30344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba3, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba4, value : 32'h84d8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba5, value : 32'h79af036e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba6, value : 32'ha00c8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba7, value : 32'h2d404002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba8, value : 32'h244a138b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ba9, value : 32'h708d7280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53baa, value : 32'h20a8706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bab, value : 32'h82b0680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bac, value : 32'h240500ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bad, value : 32'h210512c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bae, value : 32'h90040f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53baf, value : 32'h210502dc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb0, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb1, value : 32'h924002e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb2, value : 32'h213d9120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb3, value : 32'h793b0081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb4, value : 32'h67796949},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb5, value : 32'h2480a940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb6, value : 32'h71641010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb7, value : 32'h71a5e70a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb8, value : 32'hc6c8f1d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bb9, value : 32'hfeac2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bba, value : 32'h450801e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bbb, value : 32'h1600e888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bbc, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bbd, value : 32'h811000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bbe, value : 32'h40a100bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bbf, value : 32'h22008b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc0, value : 32'hc6c240a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc1, value : 32'hfd2f0ab6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc2, value : 32'hc6c2702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc3, value : 32'h1600c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc4, value : 32'h8000708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc5, value : 32'h47280008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc6, value : 32'hf92f0b86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc7, value : 32'h700c4508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc8, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bc9, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bca, value : 32'hbba70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bcb, value : 32'h70ccf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bcc, value : 32'h10802678},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bcd, value : 32'he5a781b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bce, value : 32'h68c2f96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bcf, value : 32'h700cef11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd0, value : 32'h724cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd1, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd2, value : 32'hb9a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd3, value : 32'h74ccf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd4, value : 32'h752c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd5, value : 32'h238a4040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd6, value : 32'hb8950004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd7, value : 32'h704cf01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd8, value : 32'h4040752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bd9, value : 32'h4238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bda, value : 32'h708cb895},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bdb, value : 32'hb7645a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bdc, value : 32'h70ccf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bdd, value : 32'hd92b74ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bde, value : 32'h42c1bf98},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bdf, value : 32'h706c40e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be0, value : 32'h45a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be1, value : 32'hf96f0b5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be2, value : 32'h40e170cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be3, value : 32'h42c1d92b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be4, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be5, value : 32'hb4e45a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be6, value : 32'h70ccf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be7, value : 32'hd92bd841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be8, value : 32'h42c1b812},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53be9, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bea, value : 32'hb3a45a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53beb, value : 32'h70ccf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bec, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bed, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bee, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bef, value : 32'hf96f0b26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf0, value : 32'h280264a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf1, value : 32'hd907706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf2, value : 32'h744c4060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf3, value : 32'h708cb88f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf4, value : 32'hb1270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf5, value : 32'h70ccf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf6, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf7, value : 32'h706cda08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf8, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bf9, value : 32'hf96f0afe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bfa, value : 32'hd8e70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bfb, value : 32'h700cf94f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bfc, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bfd, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bfe, value : 32'haea70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53bff, value : 32'h70ccf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c00, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c01, value : 32'h2482c3f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c02, value : 32'h42103403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c03, value : 32'h38002455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c04, value : 32'h702c4330},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c05, value : 32'hf8af08ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c06, value : 32'h40c3da50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c07, value : 32'hf0b00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c08, value : 32'hb415448b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c09, value : 32'h73044899},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c0a, value : 32'hb409b42f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c0b, value : 32'ha812057},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c0c, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c0d, value : 32'h1c66ff74},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c0e, value : 32'h21573004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c0f, value : 32'h1c5a09c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c10, value : 32'hb86e3004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c11, value : 32'h30041c42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c12, value : 32'hb41bb863},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c13, value : 32'h140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c14, value : 32'hda07f0ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c15, value : 32'h1c5c686e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c16, value : 32'h71ad3084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c17, value : 32'h30841c44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c18, value : 32'h2342b45c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c19, value : 32'hc0490342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c1a, value : 32'h140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c1b, value : 32'hc043ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c1c, value : 32'h3392080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c1d, value : 32'hda40c240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c1e, value : 32'h30841c6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c1f, value : 32'h8022040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c20, value : 32'hc258c05b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c21, value : 32'h77046843},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c22, value : 32'hc04fb423},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c23, value : 32'h41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c24, value : 32'h1600fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c25, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c26, value : 32'h20790008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c27, value : 32'h1c4e0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c28, value : 32'h1c403044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c29, value : 32'h702c3004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c2a, value : 32'hb802b41d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c2b, value : 32'h42c3c255},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c2c, value : 32'hf0040007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c2d, value : 32'hc809b417},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c2e, value : 32'hb42bb42e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c2f, value : 32'h1c70b425},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c30, value : 32'h1c643044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c31, value : 32'h1c5e3044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c32, value : 32'h1c583044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c33, value : 32'h1c523044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c34, value : 32'h1c4c3044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c35, value : 32'hc2523044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c36, value : 32'h1c466b4b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c37, value : 32'hb43a3044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c38, value : 32'hf812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c39, value : 32'hf00b000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c3a, value : 32'h2254c15e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c3b, value : 32'h78250941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c3c, value : 32'h1c72c346},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c3d, value : 32'hb8303004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c3e, value : 32'h702cc24c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c3f, value : 32'h30041c74},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c40, value : 32'h704c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c41, value : 32'hb4b6706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c42, value : 32'hb4aab4b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c43, value : 32'h1c68b4a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c44, value : 32'h1c503344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c45, value : 32'hb4b43344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c46, value : 32'hb4a8b4b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c47, value : 32'h30851c04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c48, value : 32'h30851c7c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c49, value : 32'hfcef0d7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c4a, value : 32'h33441c76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c4b, value : 32'h42c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c4c, value : 32'h700c5555},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c4d, value : 32'h4340722c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c4e, value : 32'hcde4440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c4f, value : 32'h4540fcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c50, value : 32'h98ac080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c51, value : 32'hd97e0260},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c52, value : 32'ha9ed80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c53, value : 32'hd90ffa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c54, value : 32'h900741d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c55, value : 32'h1900f804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c56, value : 32'h47cb2105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c57, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c58, value : 32'h6832c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c59, value : 32'h2105d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c5a, value : 32'h90070f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c5b, value : 32'hb200fc48},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c5c, value : 32'hf822105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c5d, value : 32'hfc4c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c5e, value : 32'h2105b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c5f, value : 32'h90070f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c60, value : 32'hb200fc40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c61, value : 32'hf822105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c62, value : 32'hfc449007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c63, value : 32'h2d00b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c64, value : 32'hb8021480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c65, value : 32'h200f8f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c66, value : 32'h8f01048e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c67, value : 32'ha4082b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c68, value : 32'hba0e7842},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c69, value : 32'h240a7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c6a, value : 32'h20a87000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c6b, value : 32'h210503c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c6c, value : 32'h72c30080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c6d, value : 32'h40000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c6e, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c6f, value : 32'h57c9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c70, value : 32'hbb8a9060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c71, value : 32'h8a6b060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c72, value : 32'h9defc4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c73, value : 32'h242f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c74, value : 32'hd8552387},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c75, value : 32'h704cd955},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c76, value : 32'he02706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c77, value : 32'h240a0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c78, value : 32'h40820500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c79, value : 32'hffef0d2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c7a, value : 32'hd860702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c7b, value : 32'hf96f08a6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c7c, value : 32'h208a712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c7d, value : 32'h40d30fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c7e, value : 32'hc2cc9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c7f, value : 32'h20041800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c80, value : 32'h20041804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c81, value : 32'h71001600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c82, value : 32'h2c09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c83, value : 32'hc002045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c84, value : 32'ha00418f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c85, value : 32'ha34418f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c86, value : 32'h8f008f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c87, value : 32'h10240c43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c88, value : 32'h2840d9ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c89, value : 32'h244a0388},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c8a, value : 32'h706d7240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c8b, value : 32'h20a8704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c8c, value : 32'hb1305c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c8d, value : 32'h20002031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c8e, value : 32'h11200681},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c8f, value : 32'ha190081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c90, value : 32'h20050040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c91, value : 32'h210512c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c92, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c93, value : 32'h916001d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c94, value : 32'hb160e320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c95, value : 32'h10102380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c96, value : 32'h71047144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c97, value : 32'h46cbf1e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c98, value : 32'h1068000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c99, value : 32'hd8538e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c9a, value : 32'hd724340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c9b, value : 32'h240a0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c9c, value : 32'h8e000500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c9d, value : 32'h8fa0e81c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c9e, value : 32'h8258f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53c9f, value : 32'h8e000344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca0, value : 32'ha008a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca1, value : 32'h2d4079af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca2, value : 32'h21051381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca3, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca4, value : 32'hb1003830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca5, value : 32'h75108f01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca6, value : 32'hf7b371a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca7, value : 32'hfc7218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca8, value : 32'h900740c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ca9, value : 32'h1800f834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53caa, value : 32'hb0220005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cab, value : 32'hc624082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cac, value : 32'h712cffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cad, value : 32'h42c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cae, value : 32'h700cac53},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53caf, value : 32'h4340722c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb0, value : 32'hb564440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb1, value : 32'h4540fcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb2, value : 32'h91ed80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb3, value : 32'hd90ffa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb4, value : 32'hdd2870cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb5, value : 32'hfbed808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb6, value : 32'h712cf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb7, value : 32'h108b1701},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb8, value : 32'hb578f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cb9, value : 32'hd90f1024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cba, value : 32'h3892840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cbb, value : 32'h7240244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cbc, value : 32'h708d700d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cbd, value : 32'h7c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cbe, value : 32'h20310b11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cbf, value : 32'h6812000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc0, value : 32'h811120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc1, value : 32'h10400c29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc2, value : 32'h12412005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc3, value : 32'h210570cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc4, value : 32'h90040f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc5, value : 32'h210502dc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc6, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc7, value : 32'h924001d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc8, value : 32'hea069160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cc9, value : 32'h8032354},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cca, value : 32'hb1604648},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ccb, value : 32'h10102080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ccc, value : 32'h71047185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ccd, value : 32'h8b2f1d7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cce, value : 32'hd80ffa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ccf, value : 32'h133f258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd0, value : 32'h10002678},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd1, value : 32'h2de41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd2, value : 32'ha9e0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd3, value : 32'h4242f8af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd4, value : 32'h38002455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd5, value : 32'hfa2712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd6, value : 32'h704cffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd7, value : 32'hfee4042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd8, value : 32'h712cfa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cd9, value : 32'hf002054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cda, value : 32'h38012455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cdb, value : 32'h706c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cdc, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cdd, value : 32'h260085a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cde, value : 32'h40c34588},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cdf, value : 32'hf8309007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce0, value : 32'h73441e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce1, value : 32'hc29c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce2, value : 32'ha34418f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce3, value : 32'h73441e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce4, value : 32'h4901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce5, value : 32'h23441900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce6, value : 32'hb0a2b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce7, value : 32'h20080a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce8, value : 32'hc7d0b0a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ce9, value : 32'hd820c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cea, value : 32'h900b45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ceb, value : 32'hb5ac280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cec, value : 32'h1d00fe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ced, value : 32'h1d001045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cee, value : 32'hc6c21005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cef, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf0, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf1, value : 32'h41db3202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf2, value : 32'hc17c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf3, value : 32'h901c43d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf4, value : 32'h190004a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf5, value : 32'h42103005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf6, value : 32'h20551b5c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf7, value : 32'hc8094338},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf8, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cf9, value : 32'hda7204b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cfa, value : 32'h71ad702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cfb, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cfc, value : 32'h180004c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cfd, value : 32'hcf20045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cfe, value : 32'hc085f86f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53cff, value : 32'h702c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d00, value : 32'ha9e704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d01, value : 32'h706cfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d02, value : 32'h722c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d03, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d04, value : 32'ha06708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d05, value : 32'h70acfcef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d06, value : 32'heb2c085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d07, value : 32'hd9720220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d08, value : 32'hfacf0fc2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d09, value : 32'hfc2d80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d0a, value : 32'hd90ff9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d0b, value : 32'hff8f0b1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d0c, value : 32'h40c3d90a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d0d, value : 32'h4e7c8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d0e, value : 32'h200e8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d0f, value : 32'h40024010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d10, value : 32'hedad90a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d11, value : 32'h704cf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d12, value : 32'hd90a4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d13, value : 32'hfdef0dba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d14, value : 32'h4002da59},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d15, value : 32'h200e6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d16, value : 32'h4002d92e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d17, value : 32'hebed92e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d18, value : 32'h704cf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d19, value : 32'he5e4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d1a, value : 32'hd9120020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d1b, value : 32'hd9124002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d1c, value : 32'hf96f0eaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d1d, value : 32'hcc2daef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d1e, value : 32'hc0810060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d1f, value : 32'hd16c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d20, value : 32'hd90afb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d21, value : 32'hd0ec081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d22, value : 32'hd92efb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d23, value : 32'hd06c081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d24, value : 32'hd912fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d25, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d26, value : 32'h41421228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d27, value : 32'h219f8f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d28, value : 32'h704c02c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d29, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d2a, value : 32'h708cc381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d2b, value : 32'h2d006119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d2c, value : 32'hb8021480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d2d, value : 32'h200f7102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d2e, value : 32'h6d12048d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d2f, value : 32'h7e0f78a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d30, value : 32'h81640c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d31, value : 32'h40d90220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d32, value : 32'hf864002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d33, value : 32'hd90affaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d34, value : 32'hf7e4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d35, value : 32'hd912ffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d36, value : 32'hf764002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d37, value : 32'hd92effaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d38, value : 32'h700c7daf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d39, value : 32'h704c702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d3a, value : 32'haf2706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d3b, value : 32'h44a10060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d3c, value : 32'h92e710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d3d, value : 32'h712c0060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d3e, value : 32'hc4e40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d3f, value : 32'h702c01e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d40, value : 32'h740cd9b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d41, value : 32'hfaef0a02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d42, value : 32'hd860b912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d43, value : 32'hf92f0d86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d44, value : 32'he6e712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d45, value : 32'h8f03fc8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d46, value : 32'h82b8f22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d47, value : 32'h78220064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d48, value : 32'h29406841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d49, value : 32'h240a0380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d4a, value : 32'h20a87080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d4b, value : 32'h20050340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d4c, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d4d, value : 32'h914001d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d4e, value : 32'h70c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d4f, value : 32'hbac54000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d50, value : 32'h700cb140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d51, value : 32'hd4e712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d52, value : 32'h1c00f92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d53, value : 32'hd80f3fc1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d54, value : 32'hf9ef0e96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d55, value : 32'h40a1d90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d56, value : 32'h1e00bee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d57, value : 32'h208a712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d58, value : 32'h46cb0fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d59, value : 32'hc2cc9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d5a, value : 32'h41c3b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d5b, value : 32'h2d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d5c, value : 32'hd881b602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d5d, value : 32'h90041ef8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d5e, value : 32'h1ef4d830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d5f, value : 32'h98a9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d60, value : 32'h740cfaef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d61, value : 32'h40a1ddff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d62, value : 32'h461045b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d63, value : 32'h700c44b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d64, value : 32'hf92f0d02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d65, value : 32'h8f03712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d66, value : 32'h8618f22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d67, value : 32'h70ee0064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d68, value : 32'h29407822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d69, value : 32'h7104038c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d6a, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d6b, value : 32'h7c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d6c, value : 32'h2405c280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d6d, value : 32'h90041f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d6e, value : 32'h900002dc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d6f, value : 32'h2079623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d70, value : 32'h8a000003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d71, value : 32'h7865781b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d72, value : 32'h2053aa00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d73, value : 32'h240580be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d74, value : 32'h90041f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d75, value : 32'h904001d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d76, value : 32'h2254f205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d77, value : 32'h71ee0802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d78, value : 32'h7124b040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d79, value : 32'h74c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d7a, value : 32'h14034000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d7b, value : 32'hc5203096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d7c, value : 32'h30951402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d7d, value : 32'h30941401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d7e, value : 32'hdeed80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d7f, value : 32'hd90ff9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d80, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d81, value : 32'h402d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d82, value : 32'h438242a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d83, value : 32'h540240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d84, value : 32'hfaef08f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d85, value : 32'h580250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d86, value : 32'h90b7126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d87, value : 32'hf732e15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d88, value : 32'hdd5ba011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d89, value : 32'h20002778},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d8a, value : 32'hfbebd13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d8b, value : 32'h41a1f86f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d8c, value : 32'h1401254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d8d, value : 32'hfaef08d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d8e, value : 32'h8f03740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d8f, value : 32'h82d8f22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d90, value : 32'h78220064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d91, value : 32'h29406841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d92, value : 32'h240a0380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d93, value : 32'h20a87080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d94, value : 32'h20050380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d95, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d96, value : 32'h914001d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d97, value : 32'h70c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d98, value : 32'h22554000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d99, value : 32'hb1400802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d9a, value : 32'hb6a070ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d9b, value : 32'hd12b6a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d9c, value : 32'h1ef4fcaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d9d, value : 32'h700c9344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d9e, value : 32'h200d42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53d9f, value : 32'hd881712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da0, value : 32'h2da41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da1, value : 32'h1ef80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da2, value : 32'h87e9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da3, value : 32'h740cfaef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da4, value : 32'hc02d840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da5, value : 32'h712cf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da6, value : 32'h712c4063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da7, value : 32'hffaf0c5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da8, value : 32'h8f23724c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53da9, value : 32'h9238f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53daa, value : 32'h79020024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dab, value : 32'h240a7124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dac, value : 32'h20a87040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dad, value : 32'h23f402c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dae, value : 32'h23143001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53daf, value : 32'h21803002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db0, value : 32'h7104003e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db1, value : 32'h4042b220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db2, value : 32'hfa2f0c82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db3, value : 32'h48c8712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db4, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db5, value : 32'h714c4163},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db6, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db7, value : 32'h2200cf2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db8, value : 32'hd92071ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53db9, value : 32'h900740c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dba, value : 32'hb0a0c29c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dbb, value : 32'h22c1229f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dbc, value : 32'h804418ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dbd, value : 32'h834418ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dbe, value : 32'h73441e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dbf, value : 32'hc164900b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc0, value : 32'h93441ef8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc1, value : 32'h30451900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc2, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc3, value : 32'h4c12005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc4, value : 32'hffef0c96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc5, value : 32'h8f00b1a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc6, value : 32'h209f704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc7, value : 32'hc3810582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc8, value : 32'h7042708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dc9, value : 32'h4012000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dca, value : 32'h1e00dae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dcb, value : 32'hca004003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dcc, value : 32'h10250d31},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dcd, value : 32'h138c2d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dce, value : 32'h7240244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dcf, value : 32'h702c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd0, value : 32'h38020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd1, value : 32'h2405716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd2, value : 32'h7b381080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd3, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd4, value : 32'h2f89004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd5, value : 32'h102280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd6, value : 32'hb0607124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd7, value : 32'hf1e971a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd8, value : 32'h32022480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dd9, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dda, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ddb, value : 32'h4408c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ddc, value : 32'h2084880b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ddd, value : 32'hac0b01c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dde, value : 32'hb8a38c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ddf, value : 32'h1600ac01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de0, value : 32'h800070c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de1, value : 32'h80f000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de2, value : 32'h8c130012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de3, value : 32'h3002046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de4, value : 32'h94aac13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de5, value : 32'he808f8cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de6, value : 32'hb8858c0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de7, value : 32'h8c03ac0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de8, value : 32'hac03b887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53de9, value : 32'hf9cf0a7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dea, value : 32'h8c15e807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53deb, value : 32'hac15b8a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dec, value : 32'hb8868c03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ded, value : 32'hd840ac03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dee, value : 32'h10831c14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53def, value : 32'h8c0dac10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df0, value : 32'hac0db8a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df1, value : 32'h20458c11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df2, value : 32'hac110e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df3, value : 32'h206c8c12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df4, value : 32'hac120080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df5, value : 32'h20448c1c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df6, value : 32'hac1c0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df7, value : 32'h10801429},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df8, value : 32'hc0d1b8c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53df9, value : 32'h1c297fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dfa, value : 32'h78e01002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dfb, value : 32'h40c3c5e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dfc, value : 32'h4988000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dfd, value : 32'he9328820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dfe, value : 32'ha840704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53dff, value : 32'ha5dca00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e00, value : 32'h2a400025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e01, value : 32'h244a0381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e02, value : 32'h706c7240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e03, value : 32'h90020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e04, value : 32'h802216},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e05, value : 32'h20006078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e06, value : 32'h80010f8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e07, value : 32'h6b124fa8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e08, value : 32'h20057825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e09, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e0a, value : 32'h90800200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e0b, value : 32'hb13ad80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e0c, value : 32'hb0600231},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e0d, value : 32'h22008d80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e0e, value : 32'h18200680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e0f, value : 32'h2b400302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e10, value : 32'h718d0280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e11, value : 32'h7c787825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e12, value : 32'h20057164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e13, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e14, value : 32'hb08002f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e15, value : 32'hf1d47144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e16, value : 32'h78e0c4c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e17, value : 32'hc1a2c3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e18, value : 32'h900042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e19, value : 32'h92800184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e1a, value : 32'h903841c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e1b, value : 32'h246c0184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e1c, value : 32'h91601140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e1d, value : 32'h236cb200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e1e, value : 32'hb1000140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e1f, value : 32'h9202722d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e20, value : 32'hb8c891a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e21, value : 32'h704cb280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e22, value : 32'h44cbbdc8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e23, value : 32'h5ac8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e24, value : 32'hc241b160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e25, value : 32'hb1014183},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e26, value : 32'hc809b1a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e27, value : 32'h10832415},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e28, value : 32'h30062440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e29, value : 32'h70ad720d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e2a, value : 32'hf41c7aab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e2b, value : 32'h13412415},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e2c, value : 32'h7e0583c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e2d, value : 32'h79c58123},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e2e, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e2f, value : 32'h90030f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e30, value : 32'hb99cc000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e31, value : 32'h91e0b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e32, value : 32'h134124f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e33, value : 32'hc1817f26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e34, value : 32'h34b21f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e35, value : 32'h8126f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e36, value : 32'h2c12900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e37, value : 32'hb62079e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e38, value : 32'h193f208d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e39, value : 32'h218d71ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e3a, value : 32'h714c16ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e3b, value : 32'h2042c805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e3c, value : 32'hf20e803c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e3d, value : 32'hd99c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e3e, value : 32'h28020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e3f, value : 32'hf822005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e40, value : 32'h3649004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e41, value : 32'h70c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e42, value : 32'hb2204000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e43, value : 32'h9661468b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e44, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e45, value : 32'h20070},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e46, value : 32'hdee96a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e47, value : 32'h42a1faaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e48, value : 32'hdc7fc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e49, value : 32'h2553bc09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e4a, value : 32'h68321202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e4b, value : 32'hf832105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e4c, value : 32'h20289024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e4d, value : 32'h21059300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e4e, value : 32'h90240f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e4f, value : 32'h7884202c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e50, value : 32'h8d2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e51, value : 32'h78849100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e52, value : 32'h7845b3a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e53, value : 32'h740cb100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e54, value : 32'h7141c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e55, value : 32'hdb20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e56, value : 32'h9640faaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e57, value : 32'h78e0c7c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e58, value : 32'hdc25c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e59, value : 32'h43c3bc9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e5a, value : 32'h122c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e5b, value : 32'h21056832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e5c, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e5d, value : 32'h2105c408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e5e, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e5f, value : 32'h91200408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e60, value : 32'h305c1a24},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e61, value : 32'hf812104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e62, value : 32'hff9f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e63, value : 32'h8c00b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e64, value : 32'h8b01e818},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e65, value : 32'h82d8b20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e66, value : 32'h78220064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e67, value : 32'h240a7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e68, value : 32'h20a87000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e69, value : 32'h29400400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e6a, value : 32'h26140380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e6b, value : 32'h80007042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e6c, value : 32'h2005049c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e6d, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e6e, value : 32'h9000028c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e6f, value : 32'hb2007124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e70, value : 32'h70148c1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e71, value : 32'h8b037ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e72, value : 32'h71108b22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e73, value : 32'h7cd20e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e74, value : 32'h71047822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e75, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e76, value : 32'h3c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e77, value : 32'h3802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e78, value : 32'h70422614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e79, value : 32'h49c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e7a, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e7b, value : 32'h28c9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e7c, value : 32'h71249000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e7d, value : 32'h7ee0b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e7e, value : 32'h45cbc2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e7f, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e80, value : 32'h40108dc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e81, value : 32'h85b8d01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e82, value : 32'h40c30384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e83, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e84, value : 32'h84b8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e85, value : 32'h79cf03ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e86, value : 32'h60090a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e87, value : 32'h44084002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e88, value : 32'h2e40c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e89, value : 32'h244a1382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e8a, value : 32'h68327280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e8b, value : 32'h702c7a25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e8c, value : 32'h54020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e8d, value : 32'h104e0c25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e8e, value : 32'h1500265a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e8f, value : 32'h20007834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e90, value : 32'h80010f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e91, value : 32'h29404e2c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e92, value : 32'h78450280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e93, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e94, value : 32'h3209004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e95, value : 32'hb3009000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e96, value : 32'h71c57124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e97, value : 32'hc6c8f1d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e98, value : 32'h706cc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e99, value : 32'h6852726d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e9a, value : 32'he808710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e9b, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e9c, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e9d, value : 32'hf020e888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e9e, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53e9f, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea0, value : 32'h7ce07014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea1, value : 32'h7180244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea2, value : 32'h58020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea3, value : 32'h3802b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea4, value : 32'h800044cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea5, value : 32'h784519b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea6, value : 32'h20057c74},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea7, value : 32'h90000f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea8, value : 32'h912001c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ea9, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eaa, value : 32'h1b49000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eab, value : 32'h7164b420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eac, value : 32'hb40e9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ead, value : 32'h238ddb07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eae, value : 32'h700c16ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eaf, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb0, value : 32'h21006038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb1, value : 32'h80000f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb2, value : 32'h88401888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb3, value : 32'h2100ab40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb4, value : 32'h80000f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb5, value : 32'h104b18d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb6, value : 32'hab400082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb7, value : 32'hf832100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb8, value : 32'h191e8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eb9, value : 32'h821096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eba, value : 32'h800071c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ebb, value : 32'hab401969},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ebc, value : 32'h8010e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ebd, value : 32'ha9007fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ebe, value : 32'h2142ea1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ebf, value : 32'h7ce0803c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec0, value : 32'h64020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec1, value : 32'h4831001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec2, value : 32'h4811001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec3, value : 32'h4821001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec4, value : 32'h7b25b908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec5, value : 32'h4811001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec6, value : 32'h7945b908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec7, value : 32'h7965b910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec8, value : 32'hb99cb902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ec9, value : 32'h9120b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eca, value : 32'h521801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ecb, value : 32'h1801b928},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ecc, value : 32'hf0200052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ecd, value : 32'h803c2142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ece, value : 32'h72220e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ecf, value : 32'h4831001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed0, value : 32'h4811001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed1, value : 32'h4821001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed2, value : 32'h7b25b908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed3, value : 32'h4811001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed4, value : 32'h7945b908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed5, value : 32'h4821001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed6, value : 32'h7965b910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed7, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed8, value : 32'h90030f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ed9, value : 32'h1001c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eda, value : 32'hb9080481},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53edb, value : 32'hb3207945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53edc, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53edd, value : 32'h7915793b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ede, value : 32'hf802100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53edf, value : 32'h4608000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee0, value : 32'hb0407fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee1, value : 32'h40c34100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee2, value : 32'h12e28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee3, value : 32'he8898800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee4, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee5, value : 32'h88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee6, value : 32'h1110807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee7, value : 32'h7fe0793b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee8, value : 32'h78e07830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ee9, value : 32'he0c04100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eea, value : 32'hd840f704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eeb, value : 32'hf0044831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eec, value : 32'h3f2180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eed, value : 32'h782f7fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eee, value : 32'h24056892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eef, value : 32'h90071f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef0, value : 32'h1800c2d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef1, value : 32'h40c30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef2, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef3, value : 32'h88608841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef4, value : 32'h20e07350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef5, value : 32'h4a7007cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef6, value : 32'h7104bb0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef7, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef8, value : 32'h30020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ef9, value : 32'h10c02405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53efa, value : 32'h73c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53efb, value : 32'h20054000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53efc, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53efd, value : 32'hb02002d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53efe, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53eff, value : 32'h443206f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f00, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f01, value : 32'h88201226},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f02, value : 32'h703219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f03, value : 32'h810010fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f04, value : 32'h1031a01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f05, value : 32'h77046038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f06, value : 32'h402805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f07, value : 32'haa007fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f08, value : 32'h70cdc0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f09, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f0a, value : 32'h1e00122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f0b, value : 32'h90077384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f0c, value : 32'h8ae1fed4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f0d, value : 32'h1047232f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f0e, value : 32'hf638a60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f0f, value : 32'h2b4010e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f10, value : 32'h238c038d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f11, value : 32'hf4169fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f12, value : 32'h1f822505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f13, value : 32'h3ed49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f14, value : 32'h23f091d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f15, value : 32'h2300b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f16, value : 32'h12200682},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f17, value : 32'hba0a0082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f18, value : 32'h25057d45},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f19, value : 32'h90041f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f1a, value : 32'hb2c002d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f1b, value : 32'hf1e77164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f1c, value : 32'h4028702d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f1d, value : 32'h8f9704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f1e, value : 32'haf59010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f1f, value : 32'h202f8275},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f20, value : 32'hf7499202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f21, value : 32'h124c2505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f22, value : 32'h1f8c2405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f23, value : 32'h2d49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f24, value : 32'h2180b400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f25, value : 32'h71441010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f26, value : 32'hc4c6f1ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f27, value : 32'hd32c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f28, value : 32'h4408f96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f29, value : 32'h1843256f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f2a, value : 32'h9679520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f2b, value : 32'h41c30050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f2c, value : 32'h12298000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f2d, value : 32'h800043c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f2e, value : 32'hc1b0460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f2f, value : 32'h894010f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f30, value : 32'h15307b55},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f31, value : 32'h93401081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f32, value : 32'h9321e909},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f33, value : 32'h422208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f34, value : 32'h2450f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f35, value : 32'h79551001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f36, value : 32'h621b6172},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f37, value : 32'h6852c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f38, value : 32'hf802205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f39, value : 32'h34901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f3a, value : 32'hc805b060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f3b, value : 32'h803c2042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f3c, value : 32'h700cf20d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f3d, value : 32'h2c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f3e, value : 32'h12205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f3f, value : 32'h70c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f40, value : 32'hb9924000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f41, value : 32'hb99fb99c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f42, value : 32'he9eb160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f43, value : 32'hc6c2ff8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f44, value : 32'hc809c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f45, value : 32'h120570ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f46, value : 32'h706c3608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f47, value : 32'h1202212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f48, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f49, value : 32'h68920460},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f4a, value : 32'h2250b51},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f4b, value : 32'h233dd940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f4c, value : 32'hb99f024b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f4d, value : 32'h20798900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f4e, value : 32'h23040002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f4f, value : 32'h26f4908f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f50, value : 32'hf20613c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f51, value : 32'hd10817},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f52, value : 32'hf0079623},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f53, value : 32'h808111e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f54, value : 32'hd1090b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f55, value : 32'h22089622},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f56, value : 32'h26140042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f57, value : 32'h716413c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f58, value : 32'hb142b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f59, value : 32'h13412405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f5a, value : 32'h75c3b992},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f5b, value : 32'h40000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f5c, value : 32'hb99fb99c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f5d, value : 32'hf1dab140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f5e, value : 32'h96219600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f5f, value : 32'hf96f0c52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f60, value : 32'hc2108},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f61, value : 32'h60985021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f62, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f63, value : 32'h901c0f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f64, value : 32'hb1000034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f65, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f66, value : 32'hc1a4c3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f67, value : 32'hc0804708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f68, value : 32'h200b96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f69, value : 32'hc0804528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f6a, value : 32'hfb2f0bea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f6b, value : 32'h46cbd918},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f6c, value : 32'h4e7c8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f6d, value : 32'hd91840c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f6e, value : 32'h20096a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f6f, value : 32'h78bd42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f70, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f71, value : 32'hb8c01228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f72, value : 32'h209f8920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f73, value : 32'h704c02c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f74, value : 32'h582219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f75, value : 32'h708cc380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f76, value : 32'h6d126119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f77, value : 32'h61d978a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f78, value : 32'h1a00ef6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f79, value : 32'hc7c6780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f7a, value : 32'h4528c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f7b, value : 32'hf8af0cb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f7c, value : 32'h700c4608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f7d, value : 32'h724c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f7e, value : 32'h244a43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f7f, value : 32'h45a10780},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f80, value : 32'hf8ef0ce2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f81, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f82, value : 32'hfced922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f83, value : 32'h704cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f84, value : 32'hc82700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f85, value : 32'h712cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f86, value : 32'h78e0c6c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f87, value : 32'h900742c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f88, value : 32'hb200c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f89, value : 32'hb2227fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f8a, value : 32'hc1a4c3e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f8b, value : 32'hc0804010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f8c, value : 32'hb064548},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f8d, value : 32'h47280020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f8e, value : 32'hafc3208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f8f, value : 32'h800146cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f90, value : 32'hf20c4e7c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f91, value : 32'h28c02054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f92, value : 32'hc080790f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f93, value : 32'hfb2f0b46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f94, value : 32'h40c14030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f95, value : 32'hf02c4102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f96, value : 32'hb3ac080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f97, value : 32'hd946fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f98, value : 32'hb32c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f99, value : 32'hd947fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f9a, value : 32'hb2ac080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f9b, value : 32'hd948fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f9c, value : 32'hb22c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f9d, value : 32'hd949fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f9e, value : 32'hb1ac080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53f9f, value : 32'hd94afb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa0, value : 32'hd94640c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa1, value : 32'h20089e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa2, value : 32'h40c142e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa3, value : 32'h896d947},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa4, value : 32'h42e10020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa5, value : 32'hd94840c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa6, value : 32'h20088a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa7, value : 32'h40c142e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa8, value : 32'h882d949},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fa9, value : 32'h42e10020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53faa, value : 32'hd94a40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fab, value : 32'h200876},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fac, value : 32'h79bd42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fad, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fae, value : 32'h88001228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53faf, value : 32'h209fb9c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb0, value : 32'h704c0582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb1, value : 32'h2c1219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb2, value : 32'h708cc380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb3, value : 32'h6d126119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb4, value : 32'h61d978a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb5, value : 32'h1a00e02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb6, value : 32'hc7c8780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb7, value : 32'hdb1fc0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb8, value : 32'hc8094100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fb9, value : 32'h2085bb0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fba, value : 32'hda0b08c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fbb, value : 32'hece708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fbc, value : 32'h4128fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fbd, value : 32'hc8094600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fbe, value : 32'h9012085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fbf, value : 32'hda0b4121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc0, value : 32'hfc2f0eba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc1, value : 32'hc0d1718c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc2, value : 32'h40c07fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc3, value : 32'hc8094100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc4, value : 32'h8c12085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc5, value : 32'h238ada09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc6, value : 32'h6a10008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc7, value : 32'h708cfc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc8, value : 32'h184b6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fc9, value : 32'ha8400082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fca, value : 32'h821896},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fcb, value : 32'h18e17fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fcc, value : 32'h78e00082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fcd, value : 32'h45cbc2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fce, value : 32'h4608000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fcf, value : 32'hfa2e806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd0, value : 32'h700cffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd1, value : 32'hc6c2b504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd2, value : 32'hffef0f96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd3, value : 32'hc6c29504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd4, value : 32'h4528c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd5, value : 32'hf8af0b4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd6, value : 32'h700c4608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd7, value : 32'h724c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd8, value : 32'h248a43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fd9, value : 32'h45a10141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fda, value : 32'hf8ef0b7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fdb, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fdc, value : 32'he66d922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fdd, value : 32'h704cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fde, value : 32'hb1a700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fdf, value : 32'h712cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe0, value : 32'h78e0c6c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe1, value : 32'hdd25c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe2, value : 32'h901c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe3, value : 32'hbd9f01c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe4, value : 32'h1480151b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe5, value : 32'h15c6b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe6, value : 32'hc329480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe7, value : 32'hb102ff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe8, value : 32'h8359500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fe9, value : 32'hf84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fea, value : 32'hc8090c81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53feb, value : 32'h40c36852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fec, value : 32'hc50902c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fed, value : 32'h22059020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fee, value : 32'h90240f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fef, value : 32'h9062201c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff0, value : 32'h71046917},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff1, value : 32'hb4006b37},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff2, value : 32'hf802205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff3, value : 32'h20209024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff4, value : 32'hb0207124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff5, value : 32'h78e0c6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff6, value : 32'h4588c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff7, value : 32'h47484668},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff8, value : 32'habe4030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ff9, value : 32'h4110f8af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ffa, value : 32'h800140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ffb, value : 32'h88604e90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ffc, value : 32'hbbc5700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ffd, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53ffe, value : 32'h500244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h53fff, value : 32'hae645a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54000, value : 32'h70ccf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54001, value : 32'h762c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54002, value : 32'h4322da22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54003, value : 32'h840244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54004, value : 32'had245a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54005, value : 32'h70ccf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54006, value : 32'h700cda22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54007, value : 32'h4302762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54008, value : 32'h45a14440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54009, value : 32'hf8ef0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5400a, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5400b, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5400c, value : 32'h244a43e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5400d, value : 32'h45a107c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5400e, value : 32'hf8ef0aaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5400f, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54010, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54011, value : 32'h244a43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54012, value : 32'h45a10800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54013, value : 32'hf8ef0a96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54014, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54015, value : 32'hf8ef0a3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54016, value : 32'hc6ca712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54017, value : 32'hd925c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54018, value : 32'h8900b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54019, value : 32'h7f0589fb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5401a, value : 32'h540c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5401b, value : 32'hf36cc60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5401c, value : 32'h752cfdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5401d, value : 32'hfe2f0d7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5401e, value : 32'ha264608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5401f, value : 32'hbfc1f88f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54020, value : 32'hd90c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54021, value : 32'h706cda20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54022, value : 32'h45e1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54023, value : 32'hf8ef0a56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54024, value : 32'h40c370cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54025, value : 32'h1d4c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54026, value : 32'hfdef0f0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54027, value : 32'h60dd722c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54028, value : 32'h262f700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54029, value : 32'hd9070347},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5402a, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5402b, value : 32'ha36708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5402c, value : 32'h70acf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5402d, value : 32'h920d2d41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5402e, value : 32'h700cf20d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5402f, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54030, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54031, value : 32'ha1e70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54032, value : 32'h268af8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54033, value : 32'h258c0fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54034, value : 32'h700c1dff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54035, value : 32'h744cd910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54036, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54037, value : 32'ha0645e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54038, value : 32'h70ccf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54039, value : 32'h387262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5403a, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5403b, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5403c, value : 32'h9f2708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5403d, value : 32'h70acf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5403e, value : 32'h920d2e41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5403f, value : 32'h700cf20d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54040, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54041, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54042, value : 32'h9da70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54043, value : 32'h268af8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54044, value : 32'h258c0fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54045, value : 32'hd8801dff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54046, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54047, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54048, value : 32'h9c270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54049, value : 32'h70ccf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5404a, value : 32'h96a700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5404b, value : 32'h712cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5404c, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5404d, value : 32'ha023772c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5404e, value : 32'ha021a022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5404f, value : 32'ha0207fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54050, value : 32'h4628c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54051, value : 32'h21534508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54052, value : 32'h710c0142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54053, value : 32'hf82f0b52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54054, value : 32'hbe23702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54055, value : 32'h16022644},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54056, value : 32'h8540655d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54057, value : 32'ha5007845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54058, value : 32'h78258501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54059, value : 32'hc6c4a501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5405a, value : 32'h700cc0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5405b, value : 32'hc6ad910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5405c, value : 32'h714cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5405d, value : 32'h702cd810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5405e, value : 32'hf8ef0c5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5405f, value : 32'h700c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54060, value : 32'hc56d90a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54061, value : 32'h714cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54062, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54063, value : 32'h752c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54064, value : 32'hf8ef0445},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54065, value : 32'h78e0714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54066, value : 32'hd8ac0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54067, value : 32'h208af8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54068, value : 32'h40c30b04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54069, value : 32'h4888000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5406a, value : 32'hf8ef0d8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5406b, value : 32'h710c9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5406c, value : 32'h1e00702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5406d, value : 32'h901c7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5406e, value : 32'h90204c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5406f, value : 32'h700cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54070, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54071, value : 32'hdcec350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54072, value : 32'hd90ffdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54073, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54074, value : 32'h901c41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54075, value : 32'h190004c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54076, value : 32'h11c00005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54077, value : 32'he87f8100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54078, value : 32'h800519bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54079, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5407a, value : 32'h5a91388},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5407b, value : 32'h702cfdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5407c, value : 32'h4030c2f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5407d, value : 32'h41004508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5407e, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5407f, value : 32'h88c01228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54080, value : 32'h2c1219f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54081, value : 32'h47cb40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54082, value : 32'h4e7d8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54083, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54084, value : 32'h67386119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54085, value : 32'h710c882f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54086, value : 32'h80f78b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54087, value : 32'hb8022030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54088, value : 32'hd4216c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54089, value : 32'h2145f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5408a, value : 32'h8760154},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5408b, value : 32'h200ff8af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5408c, value : 32'h87b0351},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5408d, value : 32'h40822030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5408e, value : 32'h12c1259f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5408f, value : 32'h1582269f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54090, value : 32'h1012085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54091, value : 32'h2447222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54092, value : 32'h700c7b0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54093, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54094, value : 32'h400244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54095, value : 32'h250a65dd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54096, value : 32'h67be0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54097, value : 32'h13d32532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54098, value : 32'h10901613},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54099, value : 32'hf8ef087e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5409a, value : 32'h234470cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5409b, value : 32'hf20ca213},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5409c, value : 32'h700c65eb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5409d, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5409e, value : 32'h250a718c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5409f, value : 32'h8660480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a0, value : 32'h70ccf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a1, value : 32'h20d02053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a2, value : 32'h20b1080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a3, value : 32'h8107076},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a4, value : 32'hf00df881},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a5, value : 32'h700c8e73},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a6, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a7, value : 32'h500244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a8, value : 32'h480250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540a9, value : 32'hf8ef083e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540aa, value : 32'h244f70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ab, value : 32'h252f2183},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ac, value : 32'h7b6f0447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ad, value : 32'h762cd880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ae, value : 32'h244ada22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540af, value : 32'h8260400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b0, value : 32'h70ccf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b1, value : 32'hfce700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b2, value : 32'h712cf8af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b3, value : 32'h340c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b4, value : 32'hcc2d090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b5, value : 32'h702cfdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b6, value : 32'h78e0c6d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b7, value : 32'h88945021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b8, value : 32'h69528801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540b9, value : 32'hf812205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ba, value : 32'hc054900f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540bb, value : 32'hc0206d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540bc, value : 32'hf832205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540bd, value : 32'hc02c903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540be, value : 32'h2205b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540bf, value : 32'h90070f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c0, value : 32'h2444c1f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c1, value : 32'hbcc11300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c2, value : 32'h2478b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c3, value : 32'h783b1001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c4, value : 32'h2205b300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c5, value : 32'h90070f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c6, value : 32'h7fe0c3ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c7, value : 32'h78e0b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c8, value : 32'h215fc0e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540c9, value : 32'h44cb0a03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ca, value : 32'h11428000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540cb, value : 32'h647970cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540cc, value : 32'h63959141},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540cd, value : 32'he237d04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ce, value : 32'h231510a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540cf, value : 32'h61990381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d0, value : 32'h8139123},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d1, value : 32'h79db006e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d2, value : 32'h412314},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d3, value : 32'h91226199},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d4, value : 32'h71c57d25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d5, value : 32'h40a1f1f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d6, value : 32'h78e0c4c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d7, value : 32'h901c44cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d8, value : 32'h16000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540d9, value : 32'h90047102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540da, value : 32'h94203804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540db, value : 32'h900743c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540dc, value : 32'hbaa0f804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540dd, value : 32'h7a05b9a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540de, value : 32'hb3407825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540df, value : 32'h7fe0b400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e0, value : 32'h51b04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e1, value : 32'he81fc2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e2, value : 32'h2fd41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e3, value : 32'hb7a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e4, value : 32'h740cfa6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e5, value : 32'h72ad700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e6, value : 32'hb99fd925},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e7, value : 32'h893b8940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e8, value : 32'h712c7a25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540e9, value : 32'hb9027918},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ea, value : 32'h1210f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540eb, value : 32'hf207794b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ec, value : 32'hf9af0f9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ed, value : 32'hdd2712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ee, value : 32'h258dfb8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ef, value : 32'h710c1c3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f0, value : 32'hd9bfc6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f1, value : 32'hb42d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f2, value : 32'hb912fa6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f3, value : 32'h1a43256f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f4, value : 32'hfc6f09ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f5, value : 32'h14051d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f6, value : 32'h81ed807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f7, value : 32'h1a060020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f8, value : 32'hd8103043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540f9, value : 32'h30031a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540fa, value : 32'hb500b88f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540fb, value : 32'hfeaf0bba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540fc, value : 32'hc6c2740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540fd, value : 32'hc1b6c3f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540fe, value : 32'hd8404608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h540ff, value : 32'h1000b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54100, value : 32'hace0095},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54101, value : 32'h10e50160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54102, value : 32'h70148092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54103, value : 32'h20cad80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54104, value : 32'h267c01a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54105, value : 32'h1a0b1393},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54106, value : 32'h2e013002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54107, value : 32'h7380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54108, value : 32'h20443279},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54109, value : 32'he150051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5410a, value : 32'h230411f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5410b, value : 32'h16002453},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5410c, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5410d, value : 32'he88d0161},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5410e, value : 32'h73146e0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5410f, value : 32'hd0214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54110, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54111, value : 32'h1608000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54112, value : 32'h2087014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54113, value : 32'hb5a0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54114, value : 32'h712cf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54115, value : 32'hb0f4708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54116, value : 32'he0b2011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54117, value : 32'he151290},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54118, value : 32'hc7a11d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54119, value : 32'he806f84f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5411a, value : 32'h1fc7258a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5411b, value : 32'hf004718e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5411c, value : 32'h708eddff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5411d, value : 32'hfaef0c12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5411e, value : 32'h6e0b730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5411f, value : 32'h1350831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54120, value : 32'h11412679},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54121, value : 32'h10c02679},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54122, value : 32'h502004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54123, value : 32'h82f6e0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54124, value : 32'h702c00b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54125, value : 32'h14009b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54126, value : 32'h16007014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54127, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54128, value : 32'h742c0181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54129, value : 32'h1e221ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5412a, value : 32'hf010e88e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5412b, value : 32'hf2e6e687},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5412c, value : 32'hb30e68c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5412d, value : 32'h40a100e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5412e, value : 32'h1600f00d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5412f, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54130, value : 32'he8040182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54131, value : 32'h30021a0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54132, value : 32'h42a178f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54133, value : 32'hd3a4302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54134, value : 32'h267dfd8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54135, value : 32'h21781381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54136, value : 32'h25052000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54137, value : 32'h21052495},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54138, value : 32'h70ad0012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54139, value : 32'h40d370ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5413a, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5413b, value : 32'h12672f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5413c, value : 32'h25110026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5413d, value : 32'hf28ca5c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5413e, value : 32'h416240e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5413f, value : 32'hf9af0e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54140, value : 32'h23421801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54141, value : 32'hfbaf0d66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54142, value : 32'hc0824610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54143, value : 32'hbf2702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54144, value : 32'hda50f7ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54145, value : 32'hfaef0b72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54146, value : 32'hed5730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54147, value : 32'h20251395},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54148, value : 32'hf01a0380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54149, value : 32'hf028f023},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5414a, value : 32'hf062f062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5414b, value : 32'hf060f060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5414c, value : 32'hf026f05e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5414d, value : 32'hf005f036},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5414e, value : 32'hf05af041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5414f, value : 32'h78aff001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54150, value : 32'h428279f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54151, value : 32'h200ade},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54152, value : 32'he9d43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54153, value : 32'he8d1350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54154, value : 32'hf04e12d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54155, value : 32'he6a78af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54156, value : 32'hc182ff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54157, value : 32'hb22700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54158, value : 32'h712cf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54159, value : 32'h712c710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5415a, value : 32'h78aff026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5415b, value : 32'h1e0099a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5415c, value : 32'hf03ec182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5415d, value : 32'h1e0098e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5415e, value : 32'hf03a78af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5415f, value : 32'hc18078af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54160, value : 32'h706c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54161, value : 32'hfbaf0fce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54162, value : 32'h40224110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54163, value : 32'h714cc180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54164, value : 32'h1c04716c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54165, value : 32'hfbe3001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54166, value : 32'h1c00fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54167, value : 32'hf0283001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54168, value : 32'ha6678af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54169, value : 32'h4182ff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5416a, value : 32'had6700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5416b, value : 32'h702cf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5416c, value : 32'h702c710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5416d, value : 32'hf90f0aca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5416e, value : 32'h1600f01a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5416f, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54170, value : 32'hb8e30009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54171, value : 32'hf40578af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54172, value : 32'h400cda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54173, value : 32'h79f0f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54174, value : 32'ha524282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54175, value : 32'hdb0b0020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54176, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54177, value : 32'h17c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54178, value : 32'h1e080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54179, value : 32'h7104cc23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5417a, value : 32'h301c1a23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5417b, value : 32'ha9a730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5417c, value : 32'h1800faef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5417d, value : 32'hca0a2003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5417e, value : 32'h1600e88a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5417f, value : 32'h80007081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54180, value : 32'h7baf0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54181, value : 32'ha424042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54182, value : 32'h42c2faaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54183, value : 32'h71e671a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54184, value : 32'he0df16e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54185, value : 32'he1512d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54186, value : 32'hf00f1350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54187, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54188, value : 32'h17c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54189, value : 32'h1e0813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5418a, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5418b, value : 32'h18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5418c, value : 32'h808b8e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5418d, value : 32'h1600f902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5418e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5418f, value : 32'hb8e60001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54190, value : 32'hf8e20f0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54191, value : 32'h1e0040c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54192, value : 32'h80007003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54193, value : 32'hc7d6000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54194, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54195, value : 32'h1638000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54196, value : 32'he68de806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54197, value : 32'he68af202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54198, value : 32'hffc105ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54199, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5419a, value : 32'h18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5419b, value : 32'h70edb8e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5419c, value : 32'hffef05e7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5419d, value : 32'h13e127ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5419e, value : 32'hf94f0bee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5419f, value : 32'h2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a0, value : 32'h2562840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a1, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a2, value : 32'h1838000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a3, value : 32'h1a0be803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a4, value : 32'h26053002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a5, value : 32'hddf42356},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a6, value : 32'h8d00bd9f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a7, value : 32'h5f082f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a8, value : 32'h1400866},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541a9, value : 32'hd917e813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541aa, value : 32'h85e740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ab, value : 32'hb915fa6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ac, value : 32'h10901500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ad, value : 32'h204f702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ae, value : 32'h42c22040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541af, value : 32'h78f0ad00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b0, value : 32'hfdaf0b46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b1, value : 32'h1d00726c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b2, value : 32'h78f01402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b3, value : 32'h42c2702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b4, value : 32'hffef05ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b5, value : 32'h78e0726c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b6, value : 32'hc1a1c3f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b7, value : 32'h43304550},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b8, value : 32'hfaef0ba6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541b9, value : 32'h70cd4210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ba, value : 32'h800040d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541bb, value : 32'h22531140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541bc, value : 32'h708e204d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541bd, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541be, value : 32'hb351228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541bf, value : 32'h18002030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c0, value : 32'h16002382},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c1, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c2, value : 32'h825001b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c3, value : 32'h708e007e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c4, value : 32'hfcef0e76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c5, value : 32'h8f404042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c6, value : 32'h750c4410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c7, value : 32'h17841c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c8, value : 32'h43420003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541c9, value : 32'hfa2f0fe2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ca, value : 32'h500240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541cb, value : 32'h41624042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541cc, value : 32'h87a704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541cd, value : 32'h2578fd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ce, value : 32'h71561096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541cf, value : 32'h341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d0, value : 32'hc80908d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d1, value : 32'h82221d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d2, value : 32'h8f207825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d3, value : 32'h7825b90c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d4, value : 32'h16009de},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d5, value : 32'h7dd0d940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d6, value : 32'he5ff708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d7, value : 32'h2d0096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d8, value : 32'h11c0234a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541d9, value : 32'h2005c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541da, value : 32'h8f000301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541db, value : 32'h7825b80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541dc, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541dd, value : 32'hd80003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541de, value : 32'h16009b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541df, value : 32'h238d41a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e0, value : 32'h24561d3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e1, value : 32'hf72180c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e2, value : 32'h40c2fecf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e3, value : 32'h734cc180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e4, value : 32'h708c4362},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e5, value : 32'hf7ef0f7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e6, value : 32'h1400702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e7, value : 32'h244a300b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e8, value : 32'h20a871c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541e9, value : 32'h2b0108c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ea, value : 32'h29401440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541eb, value : 32'h20442203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ec, value : 32'h8f000042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ed, value : 32'h1c209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ee, value : 32'h607870a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ef, value : 32'h882060b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f0, value : 32'ha8207945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f1, value : 32'h22002140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f2, value : 32'h10002b01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f3, value : 32'h20447126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f4, value : 32'h8f000041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f5, value : 32'h1c209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f6, value : 32'h607870a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f7, value : 32'h108060b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f8, value : 32'h79450282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541f9, value : 32'h40c3a820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541fa, value : 32'h4848000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541fb, value : 32'h661e8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541fc, value : 32'hc809f1b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541fd, value : 32'h20057885},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541fe, value : 32'h30f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h541ff, value : 32'h932f0d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54200, value : 32'h702c0160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54201, value : 32'h1dff238d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54202, value : 32'h180c2456},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54203, value : 32'hfecf0eea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54204, value : 32'h702c4042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54205, value : 32'hfb2f0d02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54206, value : 32'h20431800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54207, value : 32'hc7d44082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54208, value : 32'h2482c3fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54209, value : 32'h1cd43617},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5420a, value : 32'h41303080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5420b, value : 32'h24004710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5420c, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5420d, value : 32'h702c0380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5420e, value : 32'h8c6da78},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5420f, value : 32'h4178f7ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54210, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54211, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54212, value : 32'h8b60308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54213, value : 32'hda78f7ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54214, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54215, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54216, value : 32'h8a60290},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54217, value : 32'hda78f7ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54218, value : 32'h919704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54219, value : 32'h700f32b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5421a, value : 32'h70981600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5421b, value : 32'hc8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5421c, value : 32'h30012084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5421d, value : 32'h31982841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5421e, value : 32'h300414d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5421f, value : 32'h42e2740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54220, value : 32'h1d741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54221, value : 32'h43220005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54222, value : 32'h640250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54223, value : 32'hfa2f0e7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54224, value : 32'h600260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54225, value : 32'h702c710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54226, value : 32'h5d32800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54227, value : 32'hf9af0aae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54228, value : 32'h84b40e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54229, value : 32'h1cd83031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5422a, value : 32'hc0823000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5422b, value : 32'hfc2f0b4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5422c, value : 32'h14c841e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5422d, value : 32'h42c33101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5422e, value : 32'h9038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5422f, value : 32'h7905c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54230, value : 32'h7945b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54231, value : 32'h216d9120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54232, value : 32'h14ca0a10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54233, value : 32'h78253101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54234, value : 32'h1d841c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54235, value : 32'hb8020002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54236, value : 32'h42027845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54237, value : 32'h206d9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54238, value : 32'h740c0a0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54239, value : 32'hfa2f0e22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5423a, value : 32'h2b4043a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5423b, value : 32'hba22093},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5423c, value : 32'h2179fa6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5423d, value : 32'h1c5a334e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5423e, value : 32'h16003018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5423f, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54240, value : 32'h206d0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54241, value : 32'h70140940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54242, value : 32'h30001ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54243, value : 32'h6120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54244, value : 32'h33710919},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54245, value : 32'h30001ce0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54246, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54247, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54248, value : 32'hc234903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54249, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5424a, value : 32'hd327fdb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5424b, value : 32'h230f0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5424c, value : 32'h1cdc25d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5424d, value : 32'h24003000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5424e, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5424f, value : 32'h702c0218},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54250, value : 32'hf7af0fbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54251, value : 32'h46d3da78},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54252, value : 32'hea48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54253, value : 32'h800045d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54254, value : 32'h8b7122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54255, value : 32'h26403030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54256, value : 32'h1e0023c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54257, value : 32'h90077484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54258, value : 32'h1e00c17c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54259, value : 32'h901c7045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5425a, value : 32'hc80904a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5425b, value : 32'hb802da60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5425c, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5425d, value : 32'h504901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5425e, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5425f, value : 32'h70c51e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54260, value : 32'hc164900b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54261, value : 32'hf7af0f62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54262, value : 32'h3e402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54263, value : 32'h3e402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54264, value : 32'h1a0093a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54265, value : 32'h710cd960},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54266, value : 32'hffaf0c86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54267, value : 32'h242f712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54268, value : 32'h700c0507},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54269, value : 32'h704c702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5426a, value : 32'hffaf0e32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5426b, value : 32'h1501706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5426c, value : 32'h15002080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5426d, value : 32'h8c52082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5426e, value : 32'h784200a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5426f, value : 32'h280c2740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54270, value : 32'hc8096821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54271, value : 32'h7040240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54272, value : 32'h78020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54273, value : 32'h3012a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54274, value : 32'h3f832400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54275, value : 32'h2100000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54276, value : 32'h7b546199},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54277, value : 32'hb9027905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54278, value : 32'hb99cb992},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54279, value : 32'h9120b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5427a, value : 32'h218cb320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5427b, value : 32'h238a8005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5427c, value : 32'h21c0003c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5427d, value : 32'h240000cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5427e, value : 32'h3f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5427f, value : 32'h7b540208},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54280, value : 32'hb3207144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54281, value : 32'h14d1f03a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54282, value : 32'h232f3087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54283, value : 32'h14cc2507},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54284, value : 32'h24553083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54285, value : 32'h14d43e41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54286, value : 32'h240a3006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54287, value : 32'h14cf04c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54288, value : 32'h24403082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54289, value : 32'hce63205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5428a, value : 32'h14dcf9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5428b, value : 32'h14d13000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5428c, value : 32'h24003087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5428d, value : 32'h3f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5428e, value : 32'h14cd0184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5428f, value : 32'h240a3083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54290, value : 32'h14d404c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54291, value : 32'h24403006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54292, value : 32'h14cf3405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54293, value : 32'hd4e3082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54294, value : 32'h14dcf9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54295, value : 32'h14403000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54296, value : 32'h1c683600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54297, value : 32'h14e93018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54298, value : 32'he80c3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54299, value : 32'h1cec710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5429a, value : 32'hb8903480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5429b, value : 32'h34981c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5429c, value : 32'h30001cf0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5429d, value : 32'h30181c64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5429e, value : 32'h6e06bd08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5429f, value : 32'h212fe70d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a0, value : 32'h1c5b2447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a1, value : 32'h28403358},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a2, value : 32'h70ad2210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a3, value : 32'h30181c5d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a4, value : 32'h33d81c5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a5, value : 32'h34181c5c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a6, value : 32'h3600145e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a7, value : 32'h4907510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a8, value : 32'h145d0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542a9, value : 32'h78a23600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542aa, value : 32'h14e0790e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ab, value : 32'h29083000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ac, value : 32'h262f0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ad, value : 32'hf4aaf048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ae, value : 32'hf2aa7017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542af, value : 32'h15802532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b0, value : 32'h1507262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b1, value : 32'h78256834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b2, value : 32'hc8a41c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b3, value : 32'h780fffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b4, value : 32'he7640c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b5, value : 32'h702c0120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b6, value : 32'h20811501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b7, value : 32'h34981c60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b8, value : 32'h20801500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542b9, value : 32'h240933},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ba, value : 32'h34981c5f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542bb, value : 32'h71247902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542bc, value : 32'h7040240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542bd, value : 32'h44020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542be, value : 32'h3812840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542bf, value : 32'hf822105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c0, value : 32'h3dd09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c1, value : 32'h3f812400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c2, value : 32'h2080000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c3, value : 32'h121f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c4, value : 32'he1207104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c5, value : 32'hc36b220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c6, value : 32'hd80ffecf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c7, value : 32'hf96f08ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c8, value : 32'h208ad90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542c9, value : 32'h46cb0086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ca, value : 32'hc2c49007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542cb, value : 32'hd840b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542cc, value : 32'hf86f0f62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542cd, value : 32'h1501712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ce, value : 32'h15002081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542cf, value : 32'h9332080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d0, value : 32'h79020024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d1, value : 32'h240a7124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d2, value : 32'h20a87040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d3, value : 32'h284004c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d4, value : 32'h24000381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d5, value : 32'h3f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d6, value : 32'h7b14017c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d7, value : 32'hf822105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d8, value : 32'h1d09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542d9, value : 32'h71049220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542da, value : 32'he120b320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542db, value : 32'hbdeb220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542dc, value : 32'hd80ffecf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542dd, value : 32'hf96f0872},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542de, value : 32'hd882d90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542df, value : 32'hb600712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e0, value : 32'hf86f0f12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e1, value : 32'h1500d840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e2, value : 32'h1501208e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e3, value : 32'h8792080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e4, value : 32'h78af03a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e5, value : 32'hfa0f0b4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e6, value : 32'h2e404010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e7, value : 32'h20051380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e8, value : 32'h90040f8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542e9, value : 32'h240001d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ea, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542eb, value : 32'h9720017c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ec, value : 32'h38020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ed, value : 32'h20547822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ee, value : 32'h108801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ef, value : 32'h44200023},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f0, value : 32'h70012602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f1, value : 32'hffc00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f2, value : 32'h42c1d840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f3, value : 32'h24004831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f4, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f5, value : 32'h78b60218},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f6, value : 32'h78d44302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f7, value : 32'h41c3b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f8, value : 32'h301dd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542f9, value : 32'hfa2f0b22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542fa, value : 32'h2400740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542fb, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542fc, value : 32'h20f40210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542fd, value : 32'hb7000380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542fe, value : 32'h20801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h542ff, value : 32'h79e7610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54300, value : 32'h71c5ffe5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54301, value : 32'hfecf0b46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54302, value : 32'hf14871a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54303, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54304, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54305, value : 32'hcea0588},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54306, value : 32'hda50f7af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54307, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54308, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54309, value : 32'hcda0538},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5430a, value : 32'hda50f7af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5430b, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5430c, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5430d, value : 32'hcca04e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5430e, value : 32'hda50f7af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5430f, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54310, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54311, value : 32'hcba0498},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54312, value : 32'hda50f7af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54313, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54314, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54315, value : 32'hcaa0448},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54316, value : 32'hda50f7af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54317, value : 32'h2400702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54318, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54319, value : 32'hc9a03f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5431a, value : 32'hda50f7af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5431b, value : 32'h33710975},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5431c, value : 32'h145b6d34},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5431d, value : 32'h79053600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5431e, value : 32'h1300254e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5431f, value : 32'h4b2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54320, value : 32'h3601145c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54321, value : 32'h79a57810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54322, value : 32'h1209b804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54323, value : 32'h78253609},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54324, value : 32'h20811500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54325, value : 32'h710d7e3b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54326, value : 32'h903843c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54327, value : 32'h29400000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54328, value : 32'h1501034f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54329, value : 32'h20142081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5432a, value : 32'h8511048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5432b, value : 32'h270513a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5432c, value : 32'h14c8124c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5432d, value : 32'h27963102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5432e, value : 32'h71c51008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5432f, value : 32'h300114d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54330, value : 32'h79856159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54331, value : 32'h7965b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54332, value : 32'h14cab100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54333, value : 32'h14d83102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54334, value : 32'h61593001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54335, value : 32'hb9027985},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54336, value : 32'h19007965},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54337, value : 32'hf1e702c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54338, value : 32'h15802532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54339, value : 32'h78256834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5433a, value : 32'h507212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5433b, value : 32'h32b10917},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5433c, value : 32'ha62780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5433d, value : 32'hf004ff8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5433e, value : 32'hfb4f0d72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5433f, value : 32'h1fc7268a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54340, value : 32'h8eaf004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54341, value : 32'hde7fff8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54342, value : 32'h308114cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54343, value : 32'h3e402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54344, value : 32'h906c282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54345, value : 32'h2455f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54346, value : 32'h14dc3e4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54347, value : 32'he8263000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54348, value : 32'h308114cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54349, value : 32'h14d442e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5434a, value : 32'hc3823005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5434b, value : 32'h308014cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5434c, value : 32'h36042440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5434d, value : 32'h70ec70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5434e, value : 32'h922c741},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5434f, value : 32'hc640fbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54350, value : 32'h3e402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54351, value : 32'h704c41e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54352, value : 32'h3f842400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54353, value : 32'h5880000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54354, value : 32'h3f852400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54355, value : 32'h5380000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54356, value : 32'h3f862400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54357, value : 32'h4e80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54358, value : 32'hfbef0d62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54359, value : 32'hf025c386},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5435a, value : 32'h20008ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5435b, value : 32'h308714d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5435c, value : 32'h507222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5435d, value : 32'h308114cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5435e, value : 32'h145a4322},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5435f, value : 32'h24403604},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54360, value : 32'h14cf3205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54361, value : 32'h14d43080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54362, value : 32'hd663006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54363, value : 32'hc740f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54364, value : 32'h3f812400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54365, value : 32'h5880000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54366, value : 32'h3f822400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54367, value : 32'h5380000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54368, value : 32'h3f832400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54369, value : 32'h4e80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5436a, value : 32'hfb6f094e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5436b, value : 32'h14cdc086},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5436c, value : 32'h24003081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5436d, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5436e, value : 32'h24000184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5436f, value : 32'h3f8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54370, value : 32'h8560184},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54371, value : 32'hc284f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54372, value : 32'h300014dc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54373, value : 32'h14cde827},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54374, value : 32'h42e23081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54375, value : 32'h300514d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54376, value : 32'h14cfc384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54377, value : 32'h24403080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54378, value : 32'h70cc3804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54379, value : 32'hc74171ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5437a, value : 32'hfbef0872},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5437b, value : 32'h41e2c640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5437c, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5437d, value : 32'h1840000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5437e, value : 32'h2400714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5437f, value : 32'h3f84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54380, value : 32'h24000498},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54381, value : 32'h3f85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54382, value : 32'h24000448},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54383, value : 32'h3f86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54384, value : 32'hcb203f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54385, value : 32'hc388fbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54386, value : 32'h83ef024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54387, value : 32'h14d00200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54388, value : 32'h222f3087},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54389, value : 32'h14cd0507},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5438a, value : 32'h43223081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5438b, value : 32'h3604145a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5438c, value : 32'h34052440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5438d, value : 32'h308014cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5438e, value : 32'h300614d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5438f, value : 32'hf9ef0cb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54390, value : 32'h2400c740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54391, value : 32'h3f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54392, value : 32'h24000498},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54393, value : 32'h3f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54394, value : 32'h24000448},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54395, value : 32'h3f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54396, value : 32'h89e03f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54397, value : 32'hc088fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54398, value : 32'h20861501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54399, value : 32'h308714ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5439a, value : 32'h208c1500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5439b, value : 32'h59c74d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5439c, value : 32'h706dffed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5439d, value : 32'h1284245a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5439e, value : 32'h3f8f2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5439f, value : 32'h3080000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a0, value : 32'h3f8e2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a1, value : 32'h3800000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a2, value : 32'h7eb67fb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a3, value : 32'h7e947f94},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a4, value : 32'h1fc1218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a5, value : 32'hb71d97f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a6, value : 32'h210c11e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a7, value : 32'h14d49040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a8, value : 32'he8883000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543a9, value : 32'h16802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543aa, value : 32'h801020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ab, value : 32'h10000b55},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ac, value : 32'h11082300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ad, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ae, value : 32'h5380000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543af, value : 32'h20220f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b0, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b1, value : 32'h4e80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b2, value : 32'h20020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b3, value : 32'h96004853},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b4, value : 32'hb6006078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b5, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b6, value : 32'h4480000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b7, value : 32'h20220f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b8, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543b9, value : 32'h3f80000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ba, value : 32'h20020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543bb, value : 32'h97407842},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543bc, value : 32'h7810621a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543bd, value : 32'h2492009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543be, value : 32'h20097870},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543bf, value : 32'hb7400041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c0, value : 32'hf1cb7165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c1, value : 32'h9700f745},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c2, value : 32'h4121b600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c3, value : 32'hf407f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c4, value : 32'h96209700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c5, value : 32'h804408f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c6, value : 32'h2400f1f9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c7, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c8, value : 32'h78b60290},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543c9, value : 32'h71857894},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ca, value : 32'hf1a2b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543cb, value : 32'h30300847},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543cc, value : 32'h3e402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543cd, value : 32'h74841e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ce, value : 32'hc164900b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543cf, value : 32'h6832c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d0, value : 32'h901c40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d1, value : 32'h79050504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d2, value : 32'h4841900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d3, value : 32'h18a4d920},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d4, value : 32'h40c38484},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d5, value : 32'hc17c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d6, value : 32'h451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d7, value : 32'h74841e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d8, value : 32'hfed49007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543d9, value : 32'h5c1886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543da, value : 32'hff2f0c3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543db, value : 32'h49c1886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543dc, value : 32'hf5ef005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543dd, value : 32'h14ccf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543de, value : 32'h15003081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543df, value : 32'h40c3208f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e0, value : 32'h7070707},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e1, value : 32'h30181c5f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e2, value : 32'h20801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e3, value : 32'h3f8e2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e4, value : 32'h17c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e5, value : 32'h24a7710},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e6, value : 32'h41e2002d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e7, value : 32'h70ad66fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e8, value : 32'h708e714e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543e9, value : 32'h70ce706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ea, value : 32'h3600145d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543eb, value : 32'h790e78a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ec, value : 32'h300014e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ed, value : 32'h12908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ee, value : 32'hf048262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ef, value : 32'h81df434},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f0, value : 32'h42e13030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f1, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f2, value : 32'h2180000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f3, value : 32'h20f478b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f4, value : 32'h210a03d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f5, value : 32'hf01b2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f6, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f7, value : 32'h3800000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f8, value : 32'h41c378b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543f9, value : 32'h401e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543fa, value : 32'h20f443a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543fb, value : 32'h240003d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543fc, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543fd, value : 32'h78b60290},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543fe, value : 32'h440250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h543ff, value : 32'h3d020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54400, value : 32'hf06740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54401, value : 32'h240af9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54402, value : 32'h200c0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54403, value : 32'hf705a580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54404, value : 32'hb21f410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54405, value : 32'haea02445},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54406, value : 32'h260a718e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54407, value : 32'h230a2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54408, value : 32'h714e2440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54409, value : 32'h145e71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5440a, value : 32'hd813600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5440b, value : 32'hf00d9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5440c, value : 32'h20300c13},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5440d, value : 32'ha580200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5440e, value : 32'ha4c121cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5440f, value : 32'h206122c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54410, value : 32'h708ef3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54411, value : 32'h202ff1f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54412, value : 32'h214c0487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54413, value : 32'h6829b340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54414, value : 32'h300014e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54415, value : 32'h8e00790c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54416, value : 32'h783d7914},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54417, value : 32'hae007d0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54418, value : 32'h740cf489},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54419, value : 32'h1e741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5441a, value : 32'h42e10003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5441b, value : 32'he9a43a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5441c, value : 32'h240af9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5441d, value : 32'h740c04c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5441e, value : 32'h1e841c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5441f, value : 32'h42e10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54420, value : 32'hf9ef0e86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54421, value : 32'h122343a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54422, value : 32'h41c33704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54423, value : 32'h301e9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54424, value : 32'h100202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54425, value : 32'h78f642e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54426, value : 32'h70c343a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54427, value : 32'h4d4c8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54428, value : 32'he66b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54429, value : 32'h740cf9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5442a, value : 32'h310114c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5442b, value : 32'h13482f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5442c, value : 32'h360b1209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5442d, value : 32'h1306254e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5442e, value : 32'h300014d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5442f, value : 32'h120c2305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54430, value : 32'h145c6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54431, value : 32'h78853601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54432, value : 32'h903843c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54433, value : 32'hb8020000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54434, value : 32'h2e4079a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54435, value : 32'h78650102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54436, value : 32'h20007a25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54437, value : 32'h1f89},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54438, value : 32'hb0401000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54439, value : 32'h124e2305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5443a, value : 32'h310014c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5443b, value : 32'h300114d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5443c, value : 32'h78c56038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5443d, value : 32'h7865b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5443e, value : 32'h14cab040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5443f, value : 32'h14d83100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54440, value : 32'h60383001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54441, value : 32'h78856d34},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54442, value : 32'h360c145b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54443, value : 32'h2405b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54444, value : 32'h7865118c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54445, value : 32'hb0807c25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54446, value : 32'h310114ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54447, value : 32'h300014d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54448, value : 32'h78c56038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54449, value : 32'h7865b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5444a, value : 32'h1600b080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5444b, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5444c, value : 32'h8a9017c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5444d, value : 32'h1600001f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5444e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5444f, value : 32'h89d0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54450, value : 32'h2305013f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54451, value : 32'h40c315cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54452, value : 32'h15409038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54453, value : 32'h12032305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54454, value : 32'h2305bb02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54455, value : 32'hb1400001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54456, value : 32'h12412305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54457, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54458, value : 32'h2054000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54459, value : 32'h7b050800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5445a, value : 32'hb5407825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5445b, value : 32'hb080b380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5445c, value : 32'hd6ef034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5445d, value : 32'h40a1f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5445e, value : 32'h32b1091f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5445f, value : 32'h8394608},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54460, value : 32'hd8403030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54461, value : 32'h1ea41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54462, value : 32'h20020003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54463, value : 32'h740c04c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54464, value : 32'h43a142e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54465, value : 32'h740cf018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54466, value : 32'h1ed41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54467, value : 32'h42e10003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54468, value : 32'hd6643a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54469, value : 32'h240af9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5446a, value : 32'h740c04c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5446b, value : 32'h1ee41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5446c, value : 32'hf0100002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5446d, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5446e, value : 32'h301eb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5446f, value : 32'h43a142e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54470, value : 32'h4c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54471, value : 32'hf9cf0d42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54472, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54473, value : 32'h201ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54474, value : 32'hd3642e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54475, value : 32'h43c1f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54476, value : 32'hffef05b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54477, value : 32'h240071e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54478, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54479, value : 32'habe017c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5447a, value : 32'h42230160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5447b, value : 32'h30310893},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5447c, value : 32'h95a40e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5447d, value : 32'h702cf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5447e, value : 32'h4210d9e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5447f, value : 32'hd0ab911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54480, value : 32'h740cf9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54481, value : 32'h20901500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54482, value : 32'h24132240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54483, value : 32'h24922240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54484, value : 32'h1407272f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54485, value : 32'h20801501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54486, value : 32'h3e40863},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54487, value : 32'h13112f40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54488, value : 32'h275f70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54489, value : 32'hc0821501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5448a, value : 32'h43a142e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5448b, value : 32'h740c603e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5448c, value : 32'h41c37eb4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5448d, value : 32'h401cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5448e, value : 32'h11051620},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5448f, value : 32'hf9ef0cca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54490, value : 32'h11041670},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54491, value : 32'h12012d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54492, value : 32'h2105c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54493, value : 32'h43c30441},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54494, value : 32'h9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54495, value : 32'h71a57825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54496, value : 32'h4812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54497, value : 32'h4c02005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54498, value : 32'h96306952},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54499, value : 32'hb8027a65},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5449a, value : 32'h7865b220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5449b, value : 32'h11011670},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5449c, value : 32'h92740db3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5449d, value : 32'h7106b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5449e, value : 32'hd76f1cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5449f, value : 32'h1600ff0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a0, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a1, value : 32'h8190009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a2, value : 32'h218a00bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a3, value : 32'h14d40fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a4, value : 32'h70143000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a5, value : 32'he1ad8ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a6, value : 32'h703cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a7, value : 32'h78e0c7da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a8, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544a9, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544aa, value : 32'h40103d06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ab, value : 32'hda78702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ac, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ad, value : 32'h13c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ae, value : 32'hc1504528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544af, value : 32'hc14ec14f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b0, value : 32'hc14cc14d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b1, value : 32'hc14ac14b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b2, value : 32'hf76f0e36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b3, value : 32'h2455c149},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b4, value : 32'h702c3c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b5, value : 32'hf76f0e2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b6, value : 32'h2455da78},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b7, value : 32'h702c3880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b8, value : 32'hc548da3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544b9, value : 32'hf76f0e1a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ba, value : 32'hc093c547},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544bb, value : 32'he12702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544bc, value : 32'hda3cf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544bd, value : 32'hc552712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544be, value : 32'h70441e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544bf, value : 32'h4a8901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c0, value : 32'hc546c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c1, value : 32'h6852c545},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c2, value : 32'hf802205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c3, value : 32'h504901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c4, value : 32'h2205b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c5, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c6, value : 32'h90000090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c7, value : 32'hf832205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c8, value : 32'hc0909007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544c9, value : 32'hb888c042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ca, value : 32'h1600b300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544cb, value : 32'h80007083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544cc, value : 32'h16000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544cd, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ce, value : 32'h811017c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544cf, value : 32'h2205001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d0, value : 32'h903b0f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d1, value : 32'hb020c234},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d2, value : 32'h40e2900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d3, value : 32'h7fcfbbc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d4, value : 32'h40e1752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d5, value : 32'hfa2f0a12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d6, value : 32'h44d3c343},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d7, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d8, value : 32'h208d1400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544d9, value : 32'h35112440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544da, value : 32'h20801401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544db, value : 32'h3640841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544dc, value : 32'h160040e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544dd, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544de, value : 32'h83112e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544df, value : 32'h4002036e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e0, value : 32'hfbef0da2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e1, value : 32'he81241a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e2, value : 32'h742c78af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e3, value : 32'hfeaf0e1e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e4, value : 32'h42004202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e5, value : 32'h23402114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e6, value : 32'h41c343a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e7, value : 32'h201a9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e8, value : 32'hb66b040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544e9, value : 32'h750cf9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ea, value : 32'hf1e071a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544eb, value : 32'hfa2f09ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ec, value : 32'h1400762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ed, value : 32'h706f208d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ee, value : 32'h20801401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ef, value : 32'h364084d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f0, value : 32'h16006e12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f1, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f2, value : 32'h83d12e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f3, value : 32'h4002036e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f4, value : 32'hfbef0d52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f5, value : 32'he81841a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f6, value : 32'h20f4c085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f7, value : 32'h8290340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f8, value : 32'h78af0071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544f9, value : 32'hdc6742c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544fa, value : 32'h4202feaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544fb, value : 32'h750c4708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544fc, value : 32'h41c342e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544fd, value : 32'h201aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544fe, value : 32'hf9ef0b0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h544ff, value : 32'hf0943a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54500, value : 32'h716f11d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54501, value : 32'hf1da71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54502, value : 32'h78cf7e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54503, value : 32'hf82f093e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54504, value : 32'hc044c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54505, value : 32'h60640c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54506, value : 32'hc0510606},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54507, value : 32'h2005c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54508, value : 32'h14b70400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54509, value : 32'hb8022097},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5450a, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5450b, value : 32'h15409038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5450c, value : 32'h1181000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5450d, value : 32'h1401d80d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5450e, value : 32'h2084208f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5450f, value : 32'hc041300c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54510, value : 32'h20831400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54511, value : 32'h35c7212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54512, value : 32'hdec0c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54513, value : 32'h40b2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54514, value : 32'h10c40f9b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54515, value : 32'h30ee0993},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54516, value : 32'h2b40c591},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54517, value : 32'h65690342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54518, value : 32'h6002105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54519, value : 32'h4e31b904},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5451a, value : 32'h22057905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5451b, value : 32'h284002c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5451c, value : 32'h22960088},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5451d, value : 32'h20050008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5451e, value : 32'h90381f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5451f, value : 32'hb0201540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54520, value : 32'h20056568},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54521, value : 32'hb8040601},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54522, value : 32'h79054e10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54523, value : 32'h2c02205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54524, value : 32'h42c36892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54525, value : 32'h15809038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54526, value : 32'h1f802405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54527, value : 32'h15409038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54528, value : 32'h6568b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54529, value : 32'h6012005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5452a, value : 32'h4e10b804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5452b, value : 32'h20057905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5452c, value : 32'hb0201080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5452d, value : 32'h65687a85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5452e, value : 32'h6012005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5452f, value : 32'h4e10b804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54530, value : 32'h702c7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54531, value : 32'hc08db200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54532, value : 32'hb0207874},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54533, value : 32'h7874c08f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54534, value : 32'hc08bb020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54535, value : 32'hb0207874},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54536, value : 32'h7874c089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54537, value : 32'h30300b0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54538, value : 32'h1800b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54539, value : 32'h71640045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5453a, value : 32'h70cdf1b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5453b, value : 32'h1f802632},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5453c, value : 32'hea48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5453d, value : 32'h78256834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5453e, value : 32'h8f2c100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5453f, value : 32'h780fff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54540, value : 32'hf86f0a22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54541, value : 32'ha2ed8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54542, value : 32'hc004f86f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54543, value : 32'hdae700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54544, value : 32'h712cf82f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54545, value : 32'h8d6c100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54546, value : 32'h700cff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54547, value : 32'h84ac000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54548, value : 32'hd91afa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54549, value : 32'h704e72ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5454a, value : 32'h20100a0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5454b, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5454c, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5454d, value : 32'h212fe827},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5454e, value : 32'h40020480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5454f, value : 32'hfbef0be6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54550, value : 32'h46104130},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54551, value : 32'h20532140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54552, value : 32'h41227014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54553, value : 32'h4c121ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54554, value : 32'h742c782f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54555, value : 32'hfeaf0c56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54556, value : 32'hc5924202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54557, value : 32'h75224708},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54558, value : 32'hb5004102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54559, value : 32'hfc6f0886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5455a, value : 32'he80d4042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5455b, value : 32'h23ca70d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5455c, value : 32'h202f2441},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5455d, value : 32'h742c04c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5455e, value : 32'hfeaf0c32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5455f, value : 32'h78e54202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54560, value : 32'h258db500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54561, value : 32'h714e253f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54562, value : 32'hf9ef0956},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54563, value : 32'h140078cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54564, value : 32'h4110208d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54565, value : 32'h20801401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54566, value : 32'h1347510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54567, value : 32'h2111002d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54568, value : 32'hf294b340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54569, value : 32'h208f1403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5456a, value : 32'hb7a4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5456b, value : 32'h41a1fbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5456c, value : 32'h1342273c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5456d, value : 32'h21f4c192},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5456e, value : 32'h2078008c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5456f, value : 32'h781b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54570, value : 32'h38822455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54571, value : 32'h73046862},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54572, value : 32'h10c12c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54573, value : 32'h21447c19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54574, value : 32'h255a0043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54575, value : 32'hc09313c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54576, value : 32'h6119623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54577, value : 32'h61d862da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54578, value : 32'h2444aa60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54579, value : 32'ha8401042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5457a, value : 32'h78b4c08b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5457b, value : 32'h9299020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5457c, value : 32'h438900e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5457d, value : 32'hc08fb060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5457e, value : 32'h902078b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5457f, value : 32'hb0806981},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54580, value : 32'h178c255a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54581, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54582, value : 32'h13c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54583, value : 32'h78346098},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54584, value : 32'h4441800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54585, value : 32'h78b4c089},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54586, value : 32'h9239020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54587, value : 32'hb0400080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54588, value : 32'h78b4c08d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54589, value : 32'h69819020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5458a, value : 32'h255ab080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5458b, value : 32'h2455178c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5458c, value : 32'h60983c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5458d, value : 32'h18007834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5458e, value : 32'he910444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5458f, value : 32'hc18f13b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54590, value : 32'h910079b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54591, value : 32'h50083d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54592, value : 32'h7074e88f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54593, value : 32'h1783255a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54594, value : 32'he7f208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54595, value : 32'h3f812400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54596, value : 32'h13c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54597, value : 32'h1e120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54598, value : 32'hb1006179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54599, value : 32'heb8ef00e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5459a, value : 32'hb1606861},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5459b, value : 32'h1783255a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5459c, value : 32'h3f812400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5459d, value : 32'h13c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5459e, value : 32'h79146179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5459f, value : 32'h1c51900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a0, value : 32'h78b4c08d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a1, value : 32'he9179020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a2, value : 32'h32c22305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a3, value : 32'h16cb2304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a4, value : 32'h10032378},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a5, value : 32'hf41a7a6b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a6, value : 32'h700931},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a7, value : 32'hb0406941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a8, value : 32'h1782255a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545a9, value : 32'h3c402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545aa, value : 32'h78346058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ab, value : 32'h1c51800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ac, value : 32'h7054f00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ad, value : 32'h1782255a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ae, value : 32'he7f208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545af, value : 32'h3c412455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b0, value : 32'h1e120ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b1, value : 32'hb1006159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b2, value : 32'hf16671a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b3, value : 32'he68f71c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b4, value : 32'hffc5061c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b5, value : 32'h41c3750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b6, value : 32'h101b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b7, value : 32'hf9ef082a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b8, value : 32'h41c34202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545b9, value : 32'h1b7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ba, value : 32'hf9ef081e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545bb, value : 32'h70ad740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545bc, value : 32'hfeede0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545bd, value : 32'h78aff9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545be, value : 32'h41c34200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545bf, value : 32'h101b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c0, value : 32'hf9ef0806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c1, value : 32'h268d740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c2, value : 32'h71a51dff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c3, value : 32'h1b941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c4, value : 32'hff60000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c5, value : 32'h740cf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c6, value : 32'h20911400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c7, value : 32'h215fc693},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c8, value : 32'h245523cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545c9, value : 32'h66be3880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ca, value : 32'h1401651d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545cb, value : 32'hf71208f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545cc, value : 32'h740c1464},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545cd, value : 32'h1ba41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ce, value : 32'hfce0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545cf, value : 32'h4222f9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d0, value : 32'h42b1df0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d1, value : 32'h24821201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d2, value : 32'h1bb41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d3, value : 32'hfba0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d4, value : 32'h740cf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d5, value : 32'h1e3f278c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d6, value : 32'h740cd96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d7, value : 32'hf9af0faa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d8, value : 32'h740cb912},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545d9, value : 32'h1bd41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545da, value : 32'hf9e0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545db, value : 32'h4222f9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545dc, value : 32'h42d1df0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545dd, value : 32'h24821201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545de, value : 32'h1be41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545df, value : 32'hf8a0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e0, value : 32'h740cf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e1, value : 32'h1e3f278d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e2, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e3, value : 32'h1bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e4, value : 32'hf98f0f76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e5, value : 32'he50fe60f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e6, value : 32'hf1c97126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e7, value : 32'h208d1400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e8, value : 32'h13640fab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545e9, value : 32'h42a14fb0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ea, value : 32'h240a7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545eb, value : 32'h20a87000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ec, value : 32'h96d0e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ed, value : 32'hc08f30ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ee, value : 32'h8120f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ef, value : 32'hb40925},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f0, value : 32'h783225a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f1, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f2, value : 32'h13c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f3, value : 32'h20146078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f4, value : 32'h98800041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f5, value : 32'h814111fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f6, value : 32'h2c44643c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f7, value : 32'hb0201081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f8, value : 32'h20f4c08d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545f9, value : 32'h2455008c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545fa, value : 32'h60783c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545fb, value : 32'h10b40c17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545fc, value : 32'h20149820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545fd, value : 32'h14fe030c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545fe, value : 32'h6199914c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h545ff, value : 32'h812944},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54600, value : 32'h2400b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54601, value : 32'h3f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54602, value : 32'hc087013c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54603, value : 32'h10c32435},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54604, value : 32'h7854792e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54605, value : 32'h2b44633b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54606, value : 32'hb0200081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54607, value : 32'hc6877144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54608, value : 32'h91f7eb4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54609, value : 32'h740c336e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5460a, value : 32'h11441600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5460b, value : 32'h41c34202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5460c, value : 32'h301c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5460d, value : 32'hf9af0ed2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5460e, value : 32'h140143a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5460f, value : 32'h72c5208f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54610, value : 32'h71a575f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54611, value : 32'h1400f7af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54612, value : 32'hf99208d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54613, value : 32'hc1871364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54614, value : 32'h79b44fb0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54615, value : 32'h240a7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54616, value : 32'h42a17000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54617, value : 32'h34020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54618, value : 32'h308e0913},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54619, value : 32'h80b9900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5461a, value : 32'hb8830052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5461b, value : 32'h7813f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5461c, value : 32'h7224b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5461d, value : 32'hf0367144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5461e, value : 32'h270479b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5461f, value : 32'h262f2040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54620, value : 32'hf22df007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54621, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54622, value : 32'h17c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54623, value : 32'hc08fe809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54624, value : 32'h34020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54625, value : 32'hc08de808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54626, value : 32'h34020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54627, value : 32'h2706e804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54628, value : 32'hf01d2057},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54629, value : 32'hc287c191},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5462a, value : 32'h22f561b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5462b, value : 32'ha190342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5462c, value : 32'h890001f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5462d, value : 32'h3310815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5462e, value : 32'h700c7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5462f, value : 32'h1c441c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54630, value : 32'hf00a0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54631, value : 32'h7704e804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54632, value : 32'hf009a900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54633, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54634, value : 32'h101c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54635, value : 32'hf76f0d12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54636, value : 32'h140142a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54637, value : 32'h71a5208f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54638, value : 32'h93650f99},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54639, value : 32'hc001712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5463a, value : 32'h262f7704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5463b, value : 32'hc041f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5463c, value : 32'h262ff205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5463d, value : 32'h34cf5c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5463e, value : 32'h1600ffc2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5463f, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54640, value : 32'h895017c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54641, value : 32'h1400001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54642, value : 32'hf8d2081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54643, value : 32'hc8091044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54644, value : 32'h903841cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54645, value : 32'h160015c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54646, value : 32'h80007088},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54647, value : 32'h200512e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54648, value : 32'h4f30040b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54649, value : 32'h240a7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5464a, value : 32'h20a87000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5464b, value : 32'h8670d80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5464c, value : 32'hc491106e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5464d, value : 32'h34d2940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5464e, value : 32'h2205642a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5464f, value : 32'h6a740600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54650, value : 32'h4a76dac0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54651, value : 32'h25057e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54652, value : 32'h687212c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54653, value : 32'h10082596},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54654, value : 32'h2402305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54655, value : 32'h6428b0c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54656, value : 32'h60e2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54657, value : 32'h4a10b804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54658, value : 32'h25057e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54659, value : 32'h68b212c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5465a, value : 32'h12402505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5465b, value : 32'h6428b0c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5465c, value : 32'h60e2005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5465d, value : 32'h4a10b804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5465e, value : 32'h21547e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5465f, value : 32'h7b051800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54660, value : 32'hb3c078a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54661, value : 32'h2305642b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54662, value : 32'hbb04060c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54663, value : 32'h7a857a62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54664, value : 32'h7124b040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54665, value : 32'h716e70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54666, value : 32'hef08724e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54667, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54668, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54669, value : 32'h100879},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5466a, value : 32'h40027efb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5466b, value : 32'hfbaf0f76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5466c, value : 32'hc18741c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5466d, value : 32'h894079d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5466e, value : 32'he8058922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5466f, value : 32'h7d4569b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54670, value : 32'h6ab4f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54671, value : 32'h710c7d25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54672, value : 32'hebe78f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54673, value : 32'h780ffa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54674, value : 32'h2347212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54675, value : 32'h4202750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54676, value : 32'h1c741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54677, value : 32'h43e10003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54678, value : 32'hf9af0d26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54679, value : 32'h440240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5467a, value : 32'hc02c100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5467b, value : 32'h4022ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5467c, value : 32'h205fc003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5467d, value : 32'h60d80b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5467e, value : 32'h70827002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5467f, value : 32'h20300815},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54680, value : 32'hb27a8b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54681, value : 32'h1e002010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54682, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54683, value : 32'hf00800f7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54684, value : 32'h20100b21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54685, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54686, value : 32'hf28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54687, value : 32'h228d71ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54688, value : 32'h706e2ffe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54689, value : 32'h1e00f00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5468a, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5468b, value : 32'hf0060101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5468c, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5468d, value : 32'hfc8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5468e, value : 32'hfa2f0e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5468f, value : 32'hc809730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54690, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54691, value : 32'h90070f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54692, value : 32'hc002c090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54693, value : 32'h2480b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54694, value : 32'h14043d06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54695, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54696, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54697, value : 32'hc1a5b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54698, value : 32'h702cc140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54699, value : 32'h9eec044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5469a, value : 32'hc000f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5469b, value : 32'h1443256f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5469c, value : 32'h8d00c043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5469d, value : 32'h900747cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5469e, value : 32'h2078c2c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5469f, value : 32'hd90f0100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a0, value : 32'he030b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a1, value : 32'h962b700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a2, value : 32'hd80ff8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a3, value : 32'h71aed9ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a4, value : 32'h208a700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a5, value : 32'hb7320fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a6, value : 32'h15441f28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a7, value : 32'h94041fdc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a8, value : 32'hb708b706},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546a9, value : 32'h15441f04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546aa, value : 32'h7054c200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ab, value : 32'h976711c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ac, value : 32'h710cff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ad, value : 32'hfacf0fb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ae, value : 32'h1097150e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546af, value : 32'h720c776e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b0, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b1, value : 32'h46d31228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b2, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b3, value : 32'h34041c0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b4, value : 32'h34041c08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b5, value : 32'h8e00c041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b6, value : 32'hd840e803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b7, value : 32'hd825f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b8, value : 32'h2d00b89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546b9, value : 32'hb9022401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ba, value : 32'h40d210f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546bb, value : 32'h7d0b8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546bc, value : 32'h40c3f2a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546bd, value : 32'h12e48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546be, value : 32'h40028020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546bf, value : 32'haeac200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c0, value : 32'hc300fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c1, value : 32'h7dafc203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c2, value : 32'he0a700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c3, value : 32'h41a1f96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c4, value : 32'hf78f0f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c5, value : 32'h702c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c6, value : 32'hf96f094a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c7, value : 32'h450842a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c8, value : 32'hf82f0c02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546c9, value : 32'hc0ed8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ca, value : 32'h78b0f82f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546cb, value : 32'h329b2440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546cc, value : 32'h32192440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546cd, value : 32'h341b2300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ce, value : 32'h34192100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546cf, value : 32'h70ad700f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d0, value : 32'h6892c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d1, value : 32'h1f802405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d2, value : 32'hc034901f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d3, value : 32'h8e23b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d4, value : 32'h9338e02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d5, value : 32'h79020024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d6, value : 32'h20831600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d7, value : 32'h28406941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d8, value : 32'h240a0381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546d9, value : 32'h20a87080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546da, value : 32'hb1303c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546db, value : 32'h2405002e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546dc, value : 32'hba921042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546dd, value : 32'hba9fba9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546de, value : 32'h7104b2a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546df, value : 32'h71c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e0, value : 32'hb864000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e1, value : 32'hd814fd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e2, value : 32'hfecf081e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e3, value : 32'h712cc004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e4, value : 32'hf7ef0f02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e5, value : 32'h8e027810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e6, value : 32'h4110704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e7, value : 32'h3942840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e8, value : 32'h83f8e03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546e9, value : 32'hd80f0464},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ea, value : 32'h20801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546eb, value : 32'h44e0827},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ec, value : 32'h2f802405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ed, value : 32'h2f49004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ee, value : 32'h22059000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ef, value : 32'he88b2012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f0, value : 32'h41c3740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f1, value : 32'h3024b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f2, value : 32'h43224202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f3, value : 32'hf9af0b3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f4, value : 32'h712644a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f5, value : 32'h2f942400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f6, value : 32'h40000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f7, value : 32'h80af1e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f8, value : 32'hd90ff8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546f9, value : 32'h3011082d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546fa, value : 32'h20310a33},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546fb, value : 32'h15c02500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546fc, value : 32'h7a10702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546fd, value : 32'hf824002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546fe, value : 32'h4150feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h546ff, value : 32'h712c4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54700, value : 32'hfeef0f76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54701, value : 32'h1b004222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54702, value : 32'h23083342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54703, value : 32'hf0062353},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54704, value : 32'h20110a0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54705, value : 32'h33421900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54706, value : 32'h71a5710f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54707, value : 32'h98d40d25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54708, value : 32'h41c34003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54709, value : 32'h10250},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5470a, value : 32'hf76f09be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5470b, value : 32'hcae4202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5470c, value : 32'hc001f94f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5470d, value : 32'h7704710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5470e, value : 32'hc0417014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5470f, value : 32'h202ff54d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54710, value : 32'h41c304ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54711, value : 32'h252},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54712, value : 32'hf76f099e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54713, value : 32'h202fb83f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54714, value : 32'h43c304c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54715, value : 32'h1328000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54716, value : 32'h140b70e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54717, value : 32'h2049308d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54718, value : 32'hc0220881},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54719, value : 32'h140a4832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5471a, value : 32'h49103080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5471b, value : 32'h802009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5471c, value : 32'hab02ab00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5471d, value : 32'h6852c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5471e, value : 32'h30801409},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5471f, value : 32'hf8c2205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54720, value : 32'hc034901f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54721, value : 32'h4834b420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54722, value : 32'h200949b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54723, value : 32'hab010300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54724, value : 32'h8e03ab03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54725, value : 32'h8378e62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54726, value : 32'h786200e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54727, value : 32'h38d2b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54728, value : 32'h40c36881},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54729, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5472a, value : 32'h240a88c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5472b, value : 32'h20a87300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5472c, value : 32'he1303c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5472d, value : 32'h220510ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5472e, value : 32'hb8920340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5472f, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54730, value : 32'h7164b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54731, value : 32'h75c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54732, value : 32'hede4000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54733, value : 32'h700cfe8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54734, value : 32'hb708b706},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54735, value : 32'hc0a5b702},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54736, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54737, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54738, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54739, value : 32'hc1bbb6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5473a, value : 32'h710c4018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5473b, value : 32'h1402800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5473c, value : 32'h2140250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5473d, value : 32'h160068b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5473e, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5473f, value : 32'h260a0162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54740, value : 32'h44702100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54741, value : 32'h47304158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54742, value : 32'hb203208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54743, value : 32'h31801c68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54744, value : 32'he899f403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54745, value : 32'he809f009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54746, value : 32'hbd41208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54747, value : 32'hbf8220cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54748, value : 32'h700000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54749, value : 32'h2050f20f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5474a, value : 32'h204a3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5474b, value : 32'h208c21c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5474c, value : 32'hf40d8802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5474d, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5474e, value : 32'h1648000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5474f, value : 32'h80802053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54750, value : 32'ha66f205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54751, value : 32'h712cf86f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54752, value : 32'h26424010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54753, value : 32'h250f20c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54754, value : 32'h212f1553},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54755, value : 32'h8232007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54756, value : 32'h706f0135},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54757, value : 32'h40c3790d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54758, value : 32'hfa88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54759, value : 32'h2022040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5475a, value : 32'h4d20f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5475b, value : 32'h5222f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5475c, value : 32'hbb8e736c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5475d, value : 32'h736cf006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5475e, value : 32'h45cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5475f, value : 32'h704effff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54760, value : 32'h44cb710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54761, value : 32'hfe030000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54762, value : 32'hb60a468b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54763, value : 32'h41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54764, value : 32'hb604f0b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54765, value : 32'h1c5c6943},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54766, value : 32'h276f3004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54767, value : 32'h1c441443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54768, value : 32'hb61c3004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54769, value : 32'h6c0ab610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5476a, value : 32'h40c3b60f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5476b, value : 32'hffb50001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5476c, value : 32'hb969b629},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5476d, value : 32'h2258b643},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5476e, value : 32'hc0400b02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5476f, value : 32'h140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54770, value : 32'h1c4efe04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54771, value : 32'h24403084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54772, value : 32'hb63b1282},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54773, value : 32'hb662489a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54774, value : 32'h743c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54775, value : 32'hc058f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54776, value : 32'h1c42b864},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54777, value : 32'h42c33084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54778, value : 32'hf0b40001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54779, value : 32'h6b0bc04c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5477a, value : 32'h6a0bc049},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5477b, value : 32'h8f00c046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5477c, value : 32'h1002078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5477d, value : 32'hb61ac152},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5477e, value : 32'hb617b962},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5477f, value : 32'he030b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54780, value : 32'hb60bc14f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54781, value : 32'hd966c080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54782, value : 32'h33041c5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54783, value : 32'h31c51c50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54784, value : 32'h31c51c2c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54785, value : 32'h36c41c2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54786, value : 32'h36c41c10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54787, value : 32'h1c0ac243},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54788, value : 32'h1c6436c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54789, value : 32'h1c5e36c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5478a, value : 32'h1c5836c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5478b, value : 32'hc35536c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5478c, value : 32'h36c41c52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5478d, value : 32'h36c41c4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5478e, value : 32'h36c41c46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5478f, value : 32'h36c41c40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54790, value : 32'h36c41c3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54791, value : 32'h31851c28},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54792, value : 32'h30851c22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54793, value : 32'he00c7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54794, value : 32'h30c51c1c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54795, value : 32'h4142d80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54796, value : 32'h43424242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54797, value : 32'hfb6f0f62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54798, value : 32'h480240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54799, value : 32'h722c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5479a, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5479b, value : 32'hfaa44a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5479c, value : 32'h45a1fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5479d, value : 32'h14c7262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5479e, value : 32'h12012d41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5479f, value : 32'h704c78af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a0, value : 32'h95a706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a1, value : 32'h44c1ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a2, value : 32'h2102217d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a3, value : 32'h407212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a4, value : 32'hfe2f0f2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a5, value : 32'h40c240c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a6, value : 32'hf8ef08d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a7, value : 32'h45cb41a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a8, value : 32'h4db48001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547a9, value : 32'hb2b43b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547aa, value : 32'h212f3135},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ab, value : 32'hc7606c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ac, value : 32'h4082ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ad, value : 32'h7280244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ae, value : 32'h20a8702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547af, value : 32'h80b0240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b0, value : 32'h1d00004e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b1, value : 32'h72a515c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b2, value : 32'h71677124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b3, value : 32'hf9ff1ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b4, value : 32'h46ea2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b5, value : 32'hb203208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b6, value : 32'h4082f406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b7, value : 32'he00d52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b8, value : 32'hf010702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547b9, value : 32'hbc01208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ba, value : 32'h40c2f406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547bb, value : 32'h1600916},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547bc, value : 32'hf0084182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547bd, value : 32'h410340a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547be, value : 32'h99e4223},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547bf, value : 32'h706c0160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c0, value : 32'hbc01208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c1, value : 32'h76f2f205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c2, value : 32'hfe610f54},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c3, value : 32'hf524082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c4, value : 32'h4082fe6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c5, value : 32'h2a102354},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c6, value : 32'h2382222f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c7, value : 32'h456a702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c8, value : 32'h21350945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547c9, value : 32'h447212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ca, value : 32'hff2f0bfa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547cb, value : 32'h704c4082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547cc, value : 32'h2950a2d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547cd, value : 32'h8e081d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ce, value : 32'h20832033},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547cf, value : 32'he90dc11a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d0, value : 32'h520b0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d1, value : 32'h79c29520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d2, value : 32'h9520b520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d3, value : 32'hb5207142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d4, value : 32'h714472a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d5, value : 32'hbf7f1ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d6, value : 32'hf1f68013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d7, value : 32'h22902040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d8, value : 32'hf1e07126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547d9, value : 32'ha0310a71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547da, value : 32'h208c464a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547db, value : 32'hf407b203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547dc, value : 32'hcbe4082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547dd, value : 32'h702c00e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547de, value : 32'h208cf00f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547df, value : 32'hf407bc01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e0, value : 32'h88240c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e1, value : 32'h41820160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e2, value : 32'h40a2f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e3, value : 32'h42234103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e4, value : 32'h1600906},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e5, value : 32'h704c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e6, value : 32'h900741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e7, value : 32'h1924c29c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e8, value : 32'h706c0015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547e9, value : 32'h70841e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ea, value : 32'hfed49007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547eb, value : 32'h708c8f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ec, value : 32'h1002078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ed, value : 32'h1904b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ee, value : 32'hd80f0014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ef, value : 32'hb144b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f0, value : 32'h1e00b146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f1, value : 32'h90077084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f2, value : 32'h1e00f804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f3, value : 32'h901f7084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f4, value : 32'hdeec004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f5, value : 32'h702cfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f6, value : 32'h1404c0bb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f7, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f8, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547f9, value : 32'hc1bab6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547fa, value : 32'h41c34510},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547fb, value : 32'h3d9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547fc, value : 32'hf96f0f16},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547fd, value : 32'h730c740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547fe, value : 32'h900741db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h547ff, value : 32'h70eec17c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54800, value : 32'hfa2f0886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54801, value : 32'h30051900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54802, value : 32'hfeef09f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54803, value : 32'h8fe40a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54804, value : 32'h710cfa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54805, value : 32'h45cbd840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54806, value : 32'h4e7c8001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54807, value : 32'hd90bb89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54808, value : 32'h10e588e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54809, value : 32'ha9e8090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5480a, value : 32'h40a1feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5480b, value : 32'ha9640a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5480c, value : 32'hd911feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5480d, value : 32'hd90bc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5480e, value : 32'hb802daf7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5480f, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54810, value : 32'hb89038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54811, value : 32'hc0409000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54812, value : 32'hf82f0ad2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54813, value : 32'h40a140a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54814, value : 32'hacad911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54815, value : 32'hdaf8f82f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54816, value : 32'hd91140a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54817, value : 32'hfcaf09aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54818, value : 32'h8d6724c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54819, value : 32'hc096ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5481a, value : 32'h92ac096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5481b, value : 32'hd90bfa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5481c, value : 32'h922c096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5481d, value : 32'hd911fa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5481e, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5481f, value : 32'h8e001228},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54820, value : 32'h209f704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54821, value : 32'hc3960582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54822, value : 32'h60b9708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54823, value : 32'ha00c4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54824, value : 32'h2705750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54825, value : 32'h40db141b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54826, value : 32'h4ec78001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54827, value : 32'h30f10b1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54828, value : 32'h30cf2378},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54829, value : 32'h704c8e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5482a, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5482b, value : 32'h708cc396},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5482c, value : 32'h6012000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5482d, value : 32'ha00c22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5482e, value : 32'h6f01d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5482f, value : 32'h903b46d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54830, value : 32'hc041c0b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54831, value : 32'h42c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54832, value : 32'hc809b5bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54833, value : 32'h718c43a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54834, value : 32'h70cc70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54835, value : 32'h68324350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54836, value : 32'h2105d870},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54837, value : 32'hb1000581},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54838, value : 32'hc02d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54839, value : 32'h218affef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5483a, value : 32'h44d30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5483b, value : 32'h4db48001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5483c, value : 32'h32112440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5483d, value : 32'h800047cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5483e, value : 32'h220a12e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5483f, value : 32'h24402500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54840, value : 32'hf413210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54841, value : 32'hd8c82135},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54842, value : 32'h82d8f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54843, value : 32'h212f05ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54844, value : 32'ha1205c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54845, value : 32'h40a2ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54846, value : 32'h7280244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54847, value : 32'h4342708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54848, value : 32'h20a84202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54849, value : 32'h80b0280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5484a, value : 32'h9320030e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5484b, value : 32'h7264b220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5484c, value : 32'h71857244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5484d, value : 32'h25122240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5484e, value : 32'h25102040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5484f, value : 32'hf1e371e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54850, value : 32'h4218a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54851, value : 32'h43a24262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54852, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54853, value : 32'hb9670cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54854, value : 32'h704effef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54855, value : 32'h2500200a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54856, value : 32'h21350a45},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54857, value : 32'h8f0040a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54858, value : 32'h4ae0831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54859, value : 32'h487212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5485a, value : 32'hff2f09ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5485b, value : 32'h244a40a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5485c, value : 32'h706d7280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5485d, value : 32'h442a4302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5485e, value : 32'h30020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5485f, value : 32'h2ce080f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54860, value : 32'h94209340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54861, value : 32'h793d6159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54862, value : 32'h7264b320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54863, value : 32'h71657285},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54864, value : 32'h25102040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54865, value : 32'h25112140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54866, value : 32'hf1e07146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54867, value : 32'he00a92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54868, value : 32'h1600702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54869, value : 32'h90387100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5486a, value : 32'hd9100034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5486b, value : 32'h42c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5486c, value : 32'h43a22798},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5486d, value : 32'h70ac718c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5486e, value : 32'hb88070cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5486f, value : 32'h1e004050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54870, value : 32'h903b7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54871, value : 32'hb1ec034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54872, value : 32'hd870ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54873, value : 32'hd910d870},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54874, value : 32'h43a24202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54875, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54876, value : 32'hffef0b0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54877, value : 32'hc80970cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54878, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54879, value : 32'hc0000581},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5487a, value : 32'h40a1b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5487b, value : 32'hfe6f0a62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5487c, value : 32'h40a1d90b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5487d, value : 32'hfe6f0a5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5487e, value : 32'hf3ed911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5487f, value : 32'hc096feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54880, value : 32'hf92c096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54881, value : 32'hd90bf9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54882, value : 32'hf8ac096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54883, value : 32'hd911f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54884, value : 32'h704c8e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54885, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54886, value : 32'h708cc396},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54887, value : 32'haba60b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54888, value : 32'h750c00a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54889, value : 32'h30f10b1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5488a, value : 32'h8e00704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5488b, value : 32'h582209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5488c, value : 32'h708cc396},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5488d, value : 32'h6012000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5488e, value : 32'ha00a9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5488f, value : 32'h70cdd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54890, value : 32'h800045cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54891, value : 32'hc001bf6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54892, value : 32'h10250e5f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54893, value : 32'h387252f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54894, value : 32'h218ad8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54895, value : 32'h42620004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54896, value : 32'h728c43a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54897, value : 32'hffef0a86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54898, value : 32'h200a70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54899, value : 32'h702e2500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5489a, value : 32'h2115093b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5489b, value : 32'h82d8f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5489c, value : 32'h212f046e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5489d, value : 32'h8ae0447},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5489e, value : 32'h40a2ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5489f, value : 32'h7280244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a0, value : 32'h4302708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a1, value : 32'h20a841a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a2, value : 32'h80b0280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a3, value : 32'h9340030e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a4, value : 32'h7264b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a5, value : 32'h71857224},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a6, value : 32'h25102040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a7, value : 32'h7126e514},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a8, value : 32'h71c5f1e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548a9, value : 32'h40a2f1d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548aa, value : 32'he00986},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ab, value : 32'he5e712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ac, value : 32'h700cf9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ad, value : 32'h30451900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ae, value : 32'h1404c0ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548af, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b0, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b1, value : 32'h2494b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b2, value : 32'hc1443ea9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b3, value : 32'hc049702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b4, value : 32'he2ec08d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b5, value : 32'hda28f6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b6, value : 32'ha8e750c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b7, value : 32'hd918f9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b8, value : 32'h800041db},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548b9, value : 32'h1100122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ba, value : 32'he3a3081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548bb, value : 32'h700cfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548bc, value : 32'h12052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548bd, value : 32'h30801100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548be, value : 32'h742c6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548bf, value : 32'h704c7e0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c0, value : 32'hfe2f0eaa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c1, value : 32'h206d40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c2, value : 32'h740c01cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c3, value : 32'h41c342a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c4, value : 32'h20338},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c5, value : 32'hf96f0bf2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c6, value : 32'hed8a43c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c7, value : 32'h33a41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c8, value : 32'hbe60000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548c9, value : 32'hd80af96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ca, value : 32'h7cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548cb, value : 32'h1243266f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548cc, value : 32'hf86f0f36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548cd, value : 32'h148f16f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ce, value : 32'h750cc04c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548cf, value : 32'hf9af0a2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d0, value : 32'h1100702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d1, value : 32'hdde3081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d2, value : 32'h700cfb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d3, value : 32'h12052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d4, value : 32'h30801100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d5, value : 32'h742c6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d6, value : 32'h704c7d0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d7, value : 32'hfe2f0e4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d8, value : 32'h206d40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548d9, value : 32'h41c301c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548da, value : 32'h20339},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548db, value : 32'hc04243a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548dc, value : 32'hb96740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548dd, value : 32'hc202f96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548de, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548df, value : 32'hf812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e0, value : 32'hc0909007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e1, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e2, value : 32'h909004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e3, value : 32'hb8899000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e4, value : 32'hc004b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e5, value : 32'h2079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e6, value : 32'hc045e008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e7, value : 32'h7014c00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e8, value : 32'h20cac005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548e9, value : 32'hc04502a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ea, value : 32'hc0438e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548eb, value : 32'h10801639},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ec, value : 32'h730c7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ed, value : 32'hf219c046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ee, value : 32'hc003c102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ef, value : 32'h700c790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f0, value : 32'h20cac047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f1, value : 32'hc04700e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f2, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f3, value : 32'h17b8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f4, value : 32'h1e081b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f5, value : 32'hc003c102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f6, value : 32'hd807790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f7, value : 32'h20cac046},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f8, value : 32'hc0460122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548f9, value : 32'h700cf003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548fa, value : 32'hc004c047},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548fb, value : 32'h2fc3268a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548fc, value : 32'h208a7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548fd, value : 32'hde250fc7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548fe, value : 32'h200226ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h548ff, value : 32'hbe9fc006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54900, value : 32'h301b141c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54901, value : 32'h2300bfc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54902, value : 32'h702e301b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54903, value : 32'hc74a700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54904, value : 32'ha6c0200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54905, value : 32'h2d0212},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54906, value : 32'hc10272ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54907, value : 32'h2400220a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54908, value : 32'h790bc003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54909, value : 32'hf20e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5490a, value : 32'h220ac006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5490b, value : 32'h200c2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5490c, value : 32'h700ca000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5490d, value : 32'h1418f7c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5490e, value : 32'hc0063012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5490f, value : 32'h400200e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54910, value : 32'h21012a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54911, value : 32'h22056852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54912, value : 32'h7a052052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54913, value : 32'h68b66834},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54914, value : 32'h728e7945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54915, value : 32'h706e7d25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54916, value : 32'h8e204262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54917, value : 32'h716e8e1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54918, value : 32'h2b007825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54919, value : 32'hb9022081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5491a, value : 32'h81210f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5491b, value : 32'hf211790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5491c, value : 32'h202f7f2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5491d, value : 32'h9260487},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5491e, value : 32'h41e1feef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5491f, value : 32'hc003c102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54920, value : 32'hf207790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54921, value : 32'hd8ff79af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54922, value : 32'hfeef09a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54923, value : 32'h248c42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54924, value : 32'h160029bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54925, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54926, value : 32'h8130001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54927, value : 32'h244a00bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54928, value : 32'h16000fc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54929, value : 32'h80007084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5492a, value : 32'hc0090120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5492b, value : 32'h42c2702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5492c, value : 32'h70ac726c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5492d, value : 32'hf8af0ed2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5492e, value : 32'h720f70ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5492f, value : 32'h25c0230a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54930, value : 32'h8e1b8e20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54931, value : 32'h790571ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54932, value : 32'h24c02f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54933, value : 32'h200fb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54934, value : 32'h782b04c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54935, value : 32'h45d3f2a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54936, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54937, value : 32'h2540231f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54938, value : 32'h308d1102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54939, value : 32'h20952d41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5493a, value : 32'h154f251f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5493b, value : 32'h1105671f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5493c, value : 32'h83b3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5493d, value : 32'h704e0364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5493e, value : 32'h800044d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5493f, value : 32'hc0051a44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54940, value : 32'h20050a25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54941, value : 32'he888c004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54942, value : 32'h16802500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54943, value : 32'h801020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54944, value : 32'h20000a0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54945, value : 32'h600a9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54946, value : 32'h23c02400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54947, value : 32'h21842480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54948, value : 32'hf1ef7146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54949, value : 32'h71a577a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5494a, value : 32'hc202f1e3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5494b, value : 32'h7a2bc103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5494c, value : 32'h1102f239},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5494d, value : 32'h8e9308d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5494e, value : 32'h25440364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5494f, value : 32'h11031052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54950, value : 32'h203c3080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54951, value : 32'h70ed0354},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54952, value : 32'hf53c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54953, value : 32'hc0041005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54954, value : 32'h2500e887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54955, value : 32'h10201680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54956, value : 32'hf3f0080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54957, value : 32'h14101000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54958, value : 32'h79b03006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54959, value : 32'h40627bf0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5495a, value : 32'h718c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5495b, value : 32'hf7ef0dd6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5495c, value : 32'h410271ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5495d, value : 32'h219a4262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5495e, value : 32'hc3970005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5495f, value : 32'h802229f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54960, value : 32'h623a6179},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54961, value : 32'h219f4182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54962, value : 32'h623a0401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54963, value : 32'h2a01225f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54964, value : 32'h7af5623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54965, value : 32'h71e5a200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54966, value : 32'h1105f1d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54967, value : 32'h71a53080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54968, value : 32'h708ef1cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54969, value : 32'h20950c79},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5496a, value : 32'h20100c09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5496b, value : 32'hf0038e1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5496c, value : 32'he8348e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5496d, value : 32'h20100c0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5496e, value : 32'h30921104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5496f, value : 32'h1102f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54970, value : 32'h24783092},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54971, value : 32'he8852000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54972, value : 32'h308f1105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54973, value : 32'h1103f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54974, value : 32'hc305308f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54975, value : 32'h14104062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54976, value : 32'h41423006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54977, value : 32'h718c42e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54978, value : 32'hf7ef0d62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54979, value : 32'h410270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5497a, value : 32'h219a4262},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5497b, value : 32'h458a0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5497c, value : 32'h802229f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5497d, value : 32'h259ac397},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5497e, value : 32'h14101401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5497f, value : 32'h728c3006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54980, value : 32'h617970ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54981, value : 32'h623ac305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54982, value : 32'h655d4142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54983, value : 32'ha50042e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54984, value : 32'hf7ef0d32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54985, value : 32'ha50a4062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54986, value : 32'hf1c67186},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54987, value : 32'h343d208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54988, value : 32'hffef05f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54989, value : 32'h40a27106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5498a, value : 32'h1600c04b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5498b, value : 32'h80007081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5498c, value : 32'h16000025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5498d, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5498e, value : 32'h79050040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5498f, value : 32'h2800710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54990, value : 32'hb8020440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54991, value : 32'h440200f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54992, value : 32'hf2b9782b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54993, value : 32'h7116700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54994, value : 32'hd016a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54995, value : 32'h2010080f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54996, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54997, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54998, value : 32'h1600f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54999, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5499a, value : 32'h70140025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5499b, value : 32'h704ef2a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5499c, value : 32'h240e2214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5499d, value : 32'h1427156},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5499e, value : 32'hc005000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5499f, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a0, value : 32'h20a8c08d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a1, value : 32'h18040140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a2, value : 32'h24000011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a3, value : 32'h3f94},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a4, value : 32'h24160afc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a5, value : 32'h706e2454},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a6, value : 32'h24142415},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a7, value : 32'h24942414},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a8, value : 32'hc003c102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549a9, value : 32'hf23e790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549aa, value : 32'h79cf70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ab, value : 32'h8f67aaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ac, value : 32'h710cf96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ad, value : 32'he988c104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ae, value : 32'h16812600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549af, value : 32'h811120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b0, value : 32'h10400d57},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b1, value : 32'h42224162},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b2, value : 32'h5219a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b3, value : 32'h229fc397},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b4, value : 32'h61790802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b5, value : 32'h4102623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b6, value : 32'h401219a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b7, value : 32'h225a623a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b8, value : 32'h61592a01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549b9, value : 32'hc08d4901},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ba, value : 32'h804078b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549bb, value : 32'h450a2b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549bc, value : 32'h211fa020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549bd, value : 32'h2f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549be, value : 32'h24000050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549bf, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c0, value : 32'h60380a5c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c1, value : 32'h2a01205a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c2, value : 32'h225a6119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c3, value : 32'h61192500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c4, value : 32'h190079b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c5, value : 32'h71a504c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c6, value : 32'hd93c005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c7, value : 32'hf0189004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c8, value : 32'h41224062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549c9, value : 32'h5209a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ca, value : 32'h219fc297},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549cb, value : 32'h60580802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549cc, value : 32'h40026119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549cd, value : 32'h401209a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ce, value : 32'h225a6119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549cf, value : 32'h61002a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d0, value : 32'h90dc10d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d1, value : 32'h1c000005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d2, value : 32'hc04d24c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d3, value : 32'ha6c0230c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d4, value : 32'hffe50750},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d5, value : 32'hc1027166},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d6, value : 32'h790bc003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d7, value : 32'h70adf21e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d8, value : 32'hc004c78d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549d9, value : 32'h2600e887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549da, value : 32'h10201680},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549db, value : 32'hd210080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549dc, value : 32'h87001000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549dd, value : 32'h700ce88c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549de, value : 32'h34041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549df, value : 32'h42220004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e0, value : 32'h240a4302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e1, value : 32'he620480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e2, value : 32'h45a1f6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e3, value : 32'hc00571a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e4, value : 32'h90240dd3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e5, value : 32'hf00e74e5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e6, value : 32'he88cc00d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e7, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e8, value : 32'h30341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549e9, value : 32'h43024222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ea, value : 32'hf6ef0e3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549eb, value : 32'h480240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ec, value : 32'h71c57146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ed, value : 32'h7106f160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ee, value : 32'h258df14b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ef, value : 32'h712e2e7c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f0, value : 32'h710c704e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f1, value : 32'h1600c048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f2, value : 32'h80007081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f3, value : 32'h16000025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f4, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f5, value : 32'h79050040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f6, value : 32'h2800710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f7, value : 32'hb8020480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f8, value : 32'h49b200f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549f9, value : 32'hb040230b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549fa, value : 32'h2102f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549fb, value : 32'hd9504042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549fc, value : 32'hf76f0932},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549fd, value : 32'h200a734c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549fe, value : 32'h24003480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h549ff, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a00, value : 32'h209f0a5c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a01, value : 32'h70ae3401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a02, value : 32'h30182000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a03, value : 32'h2d271b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a04, value : 32'hd11000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a05, value : 32'h16002010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a06, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a07, value : 32'hf0060040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a08, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a09, value : 32'h258000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a0a, value : 32'h2ac7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a0b, value : 32'h710c0021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a0c, value : 32'h5402800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a0d, value : 32'hf9ef0852},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a0e, value : 32'h252f780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a0f, value : 32'h40421540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a10, value : 32'hfb6f08e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a11, value : 32'h471041a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a12, value : 32'hc003c102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a13, value : 32'hf2c0790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a14, value : 32'h20002752},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a15, value : 32'h700e708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a16, value : 32'h23512200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a17, value : 32'h8fbc049},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a18, value : 32'hdb0820b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a19, value : 32'h2007c009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a1a, value : 32'h790f0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a1b, value : 32'h215f700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a1c, value : 32'h653e0502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a1d, value : 32'h43484330},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a1e, value : 32'h82bc105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a1f, value : 32'h796f0065},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a20, value : 32'he988c104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a21, value : 32'h16812600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a22, value : 32'h811120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a23, value : 32'h400811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a24, value : 32'h30812034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a25, value : 32'h71917c6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a26, value : 32'h4523ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a27, value : 32'h71047244},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a28, value : 32'hc006f1ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a29, value : 32'h708dc207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a2a, value : 32'h32109},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a2b, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a2c, value : 32'hafc0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a2d, value : 32'h4802016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a2e, value : 32'h5402015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a2f, value : 32'h4c02014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a30, value : 32'hc005b060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a31, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a32, value : 32'h50020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a33, value : 32'he888c004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a34, value : 32'h16802600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a35, value : 32'h801020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a36, value : 32'h10000c15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a37, value : 32'h32c02000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a38, value : 32'h79629020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a39, value : 32'h820907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a3a, value : 32'hb020c107},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a3b, value : 32'h71857265},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a3c, value : 32'h72ce70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a3d, value : 32'h244a6f72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a3e, value : 32'h702c7100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a3f, value : 32'h20a870cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a40, value : 32'h40420640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a41, value : 32'h3f822400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a42, value : 32'ha5c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a43, value : 32'h401209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a44, value : 32'h255a6058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a45, value : 32'h621a2a02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a46, value : 32'h2500235f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a47, value : 32'h20f46058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a48, value : 32'h783b00c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a49, value : 32'h71647124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a4a, value : 32'h2a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a4b, value : 32'h27147e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a4c, value : 32'h79cf140f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a4d, value : 32'hcf678ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a4e, value : 32'h222ffeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a4f, value : 32'hc00a06c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a50, value : 32'hb00205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a51, value : 32'h71ed78f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a52, value : 32'h70237022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a53, value : 32'h253f268d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a54, value : 32'h7106a8de},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a55, value : 32'h4042f185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a56, value : 32'h2a02255a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a57, value : 32'h401209f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a58, value : 32'h3f812400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a59, value : 32'ha5c0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a5a, value : 32'h621a6038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a5b, value : 32'he886c004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a5c, value : 32'h5041a24},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a5d, value : 32'h5041a10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a5e, value : 32'he886c00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a5f, value : 32'h5041a26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a60, value : 32'h5041a12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a61, value : 32'hf1b8a30},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a62, value : 32'h12242030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a63, value : 32'hb8020080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a64, value : 32'h8a127905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a65, value : 32'h7825b804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a66, value : 32'h811226},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a67, value : 32'hb902f008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a68, value : 32'h12267905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a69, value : 32'hb8040080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a6a, value : 32'h8a327825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a6b, value : 32'h222f69d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a6c, value : 32'h7e0506c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a6d, value : 32'hc76740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a6e, value : 32'h79cffeaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a6f, value : 32'h205fc00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a70, value : 32'h60b80b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a71, value : 32'h70237042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a72, value : 32'h382182e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a73, value : 32'h3f802400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a74, value : 32'hafc0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a75, value : 32'h4802016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a76, value : 32'h5402015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a77, value : 32'h20300f0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a78, value : 32'h880290e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a79, value : 32'hf004b804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a7a, value : 32'hbf049001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a7b, value : 32'h212f7f05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a7c, value : 32'h78ef06c7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a7d, value : 32'hfeaf0ba6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a7e, value : 32'hc00a4410},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a7f, value : 32'h38902140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a80, value : 32'hb00205f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a81, value : 32'h39912140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a82, value : 32'h3b932140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a83, value : 32'h434242a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a84, value : 32'h500240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a85, value : 32'h7542651d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a86, value : 32'h334e2100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a87, value : 32'h23462032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a88, value : 32'h2140aef2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a89, value : 32'h161e3a8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a8a, value : 32'h21321085},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a8b, value : 32'h67a92347},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a8c, value : 32'h23402332},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a8d, value : 32'h41c3c140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a8e, value : 32'h80342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a8f, value : 32'hccac041},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a90, value : 32'h740cf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a91, value : 32'h20300d25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a92, value : 32'hc0088e32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a93, value : 32'hc003e81d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a94, value : 32'h70421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a95, value : 32'hfb8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a96, value : 32'h790bc102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a97, value : 32'h8e3ef23c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a98, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a99, value : 32'hf02a0171},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a9a, value : 32'he81cc008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a9b, value : 32'h1e00c003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a9c, value : 32'h80007042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a9d, value : 32'hc10200f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a9e, value : 32'hf22e790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54a9f, value : 32'h40c38e3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa0, value : 32'h1678000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa1, value : 32'hc003f01a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa2, value : 32'h70421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa3, value : 32'h1008000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa4, value : 32'h790bc102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa5, value : 32'h8e3ef220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa6, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa7, value : 32'hf00e0176},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa8, value : 32'h1e00c003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aa9, value : 32'h80007042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aaa, value : 32'hc10200f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aab, value : 32'hf214790b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aac, value : 32'h40c38e3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aad, value : 32'h16c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aae, value : 32'h521801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aaf, value : 32'h23412032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab0, value : 32'h521801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab1, value : 32'h23412132},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab2, value : 32'h67a9a820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab3, value : 32'h2332a821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab4, value : 32'ha8222341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab5, value : 32'h3a182040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab6, value : 32'hffef0535},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab7, value : 32'hc00b71a6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab8, value : 32'h7704714e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ab9, value : 32'h7014c04b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aba, value : 32'h4de700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54abb, value : 32'hc048ffe2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54abc, value : 32'hf9af0d96},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54abd, value : 32'h2494730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54abe, value : 32'h14043196},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54abf, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac0, value : 32'hd76c2e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac1, value : 32'h710cf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac2, value : 32'h30641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac3, value : 32'hbfa0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac4, value : 32'hd80af92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac5, value : 32'h30741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac6, value : 32'h42c30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac7, value : 32'h24080000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac8, value : 32'hf92f0be6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ac9, value : 32'h45cbd80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aca, value : 32'h40308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54acb, value : 32'h41a1740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54acc, value : 32'h726c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54acd, value : 32'hbd2738c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ace, value : 32'h74acf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54acf, value : 32'h1401254f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad0, value : 32'h704c740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad1, value : 32'h123444c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad2, value : 32'h45c3abcd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad3, value : 32'hef12abcd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad4, value : 32'hf92f0bb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad5, value : 32'hd22db07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad6, value : 32'h700cf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad7, value : 32'h200a7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad8, value : 32'h700cd807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ad9, value : 32'hc420ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ada, value : 32'hf0007fff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54adb, value : 32'h2079c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54adc, value : 32'h4708000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54add, value : 32'h256f4e18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ade, value : 32'hb5001a43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54adf, value : 32'h10002752},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae0, value : 32'hf82f0ed6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae1, value : 32'h30021a06},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae2, value : 32'h41c3e808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae3, value : 32'h2f7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae4, value : 32'hf92f0b76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae5, value : 32'hf019d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae6, value : 32'hef06d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae7, value : 32'h2f541c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae8, value : 32'hf0050000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ae9, value : 32'h2f641c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aea, value : 32'hb5e0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aeb, value : 32'h8f6f90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aec, value : 32'he803f94f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aed, value : 32'h78dbef85},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aee, value : 32'hfeef083e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aef, value : 32'h78db7404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af0, value : 32'hfeef0836},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af1, value : 32'h70f57304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af2, value : 32'hffff40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af3, value : 32'h20c28009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af4, value : 32'h1a060061},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af5, value : 32'hb5003003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af6, value : 32'hbced8fd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af7, value : 32'h20cafd6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af8, value : 32'hc6c600e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54af9, value : 32'h7fe0710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54afa, value : 32'hc420ab},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54afb, value : 32'h1e00710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54afc, value : 32'h900c7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54afd, value : 32'h7ee00088},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54afe, value : 32'h7014c2f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54aff, value : 32'h42c3c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b00, value : 32'h1238000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b01, value : 32'h901c43c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b02, value : 32'h404804b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b03, value : 32'hf8122ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b04, value : 32'h1248000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b05, value : 32'h8b2840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b06, value : 32'h23056ba4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b07, value : 32'hdf3f10c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b08, value : 32'h23058a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b09, value : 32'h91001343},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b0a, value : 32'hbf08e50c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b0b, value : 32'h12cd2505},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b0c, value : 32'h938078e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b0d, value : 32'h784595c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b0e, value : 32'h2404b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b0f, value : 32'h7ee413c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b10, value : 32'h7ac57845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b11, value : 32'hb540b300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b12, value : 32'h901c41d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b13, value : 32'h100004e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b14, value : 32'h21401080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b15, value : 32'h16002215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b16, value : 32'h80007081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b17, value : 32'h48350124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b18, value : 32'h14402305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b19, value : 32'h254090c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b1a, value : 32'h25ce2116},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b1b, value : 32'h26531021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b1c, value : 32'h23051181},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b1d, value : 32'h23051542},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b1e, value : 32'h25001583},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b1f, value : 32'h92209057},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b20, value : 32'h1131300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b21, value : 32'h1902153},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b22, value : 32'h1a4230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b23, value : 32'h23530024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b24, value : 32'h25002194},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b25, value : 32'he943e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b26, value : 32'h25000024},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b27, value : 32'h22953e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b28, value : 32'h752c0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b29, value : 32'h942700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b2a, value : 32'hb913f6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b2b, value : 32'h6832c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b2c, value : 32'h5832105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b2d, value : 32'h5422105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b2e, value : 32'h4402105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b2f, value : 32'h7ee44328},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b30, value : 32'h23d22204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b31, value : 32'h15c12605},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b32, value : 32'h23502000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b33, value : 32'h2305b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b34, value : 32'h901c1f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b35, value : 32'h270404e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b36, value : 32'h758214cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b37, value : 32'h2005b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b38, value : 32'h7de52480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b39, value : 32'hb3a0b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b3a, value : 32'h78e0c6d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b3b, value : 32'h4628c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b3c, value : 32'h16004508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b3d, value : 32'h90307100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b3e, value : 32'h1a2203bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b3f, value : 32'he909301c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b40, value : 32'h10710e3d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b41, value : 32'h724c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b42, value : 32'h30831a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b43, value : 32'h258cf020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b44, value : 32'h4e9804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b45, value : 32'h258c0029},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b46, value : 32'h629fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b47, value : 32'h258c002c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b48, value : 32'h258c9002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b49, value : 32'hf23d9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b4a, value : 32'h9404258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b4b, value : 32'h258cf23d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b4c, value : 32'hf44f9804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b4d, value : 32'h1a07754c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b4e, value : 32'hf00a3143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b4f, value : 32'h30341c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b50, value : 32'h8a60001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b51, value : 32'h42c1f6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b52, value : 32'h30821207},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b53, value : 32'h41c3d80a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b54, value : 32'h30304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b55, value : 32'h9b243a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b56, value : 32'h44c1f92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b57, value : 32'h258cc6c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b58, value : 32'hf6d597c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b59, value : 32'h9808258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b5a, value : 32'h258cf223},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b5b, value : 32'hf2259848},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b5c, value : 32'h9f800d97},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b5d, value : 32'he9010000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b5e, value : 32'hf223f02b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b5f, value : 32'h9402258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b60, value : 32'h714cf427},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b61, value : 32'h30431a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b62, value : 32'h258cf1e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b63, value : 32'hf21d9844},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b64, value : 32'h9408258c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b65, value : 32'hda07f41d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b66, value : 32'h31c31a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b67, value : 32'h734cf1d8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b68, value : 32'h30c31a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b69, value : 32'h744cf1d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b6a, value : 32'h31031a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b6b, value : 32'hda08f1d0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b6c, value : 32'h32031a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b6d, value : 32'hda09f1cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b6e, value : 32'h32431a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b6f, value : 32'h704cf1c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b70, value : 32'h30031a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b71, value : 32'h764cf1c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b72, value : 32'h31831a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b73, value : 32'hda0af1c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b74, value : 32'h32831a07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b75, value : 32'h78e0f1bc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b76, value : 32'h8fc3208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b77, value : 32'h821f209},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b78, value : 32'h41c301d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b79, value : 32'h470901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b7a, value : 32'h451900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b7b, value : 32'h41c3f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b7c, value : 32'h470901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b7d, value : 32'h1051900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b7e, value : 32'h51900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b7f, value : 32'h903041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b80, value : 32'hb10000c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b81, value : 32'h20001d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b82, value : 32'h51904},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b83, value : 32'h903041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b84, value : 32'hb10000c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b85, value : 32'hb104b830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b86, value : 32'h200009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b87, value : 32'h51904},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b88, value : 32'h903041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b89, value : 32'h91000010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b8a, value : 32'h801f08ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b8b, value : 32'hb822155},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b8c, value : 32'h80f9200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b8d, value : 32'h1a0408b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b8e, value : 32'h1ace0045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b8f, value : 32'h9100005d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b90, value : 32'h801e08ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b91, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b92, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b93, value : 32'h1078000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b94, value : 32'h1002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b95, value : 32'hb8227fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b96, value : 32'h343226f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b97, value : 32'h500120e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b98, value : 32'h70d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b99, value : 32'h700c0c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b9a, value : 32'h7c520e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b9b, value : 32'h50112e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b9c, value : 32'hf60be1ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b9d, value : 32'h2032142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b9e, value : 32'h940b23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54b9f, value : 32'h430092b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba0, value : 32'hf20fe1c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba1, value : 32'h218cf014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba2, value : 32'hf20b8002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba3, value : 32'h8010218c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba4, value : 32'h91df211},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba5, value : 32'hf81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba6, value : 32'h8a004000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba7, value : 32'h8a00f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba8, value : 32'h80206d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ba9, value : 32'h8a00f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54baa, value : 32'hb8c0781d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bab, value : 32'h20797fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bac, value : 32'h8a000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bad, value : 32'hc0206d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bae, value : 32'h78e0f1fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54baf, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb0, value : 32'h58000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb1, value : 32'h20797fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb2, value : 32'h78e00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb3, value : 32'hf8ec0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb4, value : 32'he809ffcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb5, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb6, value : 32'hf48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb7, value : 32'h710cb8e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb8, value : 32'h700cf402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bb9, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bba, value : 32'h5c3216f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bbb, value : 32'h895a8960},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bbc, value : 32'h12384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bbd, value : 32'h811135},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bbe, value : 32'h7945bb26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bbf, value : 32'hc02178},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc0, value : 32'h78647fe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc1, value : 32'hf43216f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc2, value : 32'hb8e18900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc3, value : 32'h7ce0700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc4, value : 32'h810011e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc5, value : 32'h7000263c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc6, value : 32'hc7f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc7, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc8, value : 32'h4300c0f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bc9, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bca, value : 32'h18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bcb, value : 32'h13f0825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bcc, value : 32'heaa4428},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bcd, value : 32'hd808ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bce, value : 32'hffef0ed6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bcf, value : 32'h232f4060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd0, value : 32'hf20880c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd1, value : 32'hffef0eca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd2, value : 32'h14001404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd3, value : 32'hf3f238c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd4, value : 32'h7ee0c0d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd5, value : 32'h44cbc5e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd6, value : 32'h28f00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd7, value : 32'h30d201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd8, value : 32'h786a789b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bd9, value : 32'h184229f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bda, value : 32'h2c4160bb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bdb, value : 32'h782a1080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bdc, value : 32'h605b6078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bdd, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bde, value : 32'h22561a46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bdf, value : 32'h63080800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be0, value : 32'h12315},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be1, value : 32'h60346a0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be2, value : 32'h9236151},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be3, value : 32'h700c0324},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be4, value : 32'hf822334},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be5, value : 32'h1b488000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be6, value : 32'h22cc7150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be7, value : 32'hf7878306},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be8, value : 32'h4a907942},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54be9, value : 32'h20ca7110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bea, value : 32'hc4c20045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54beb, value : 32'h1600c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bec, value : 32'h80007101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bed, value : 32'h47c3000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bee, value : 32'h18000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bef, value : 32'h21044010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf0, value : 32'h248a01c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf1, value : 32'h27507001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf2, value : 32'h700d0307},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf3, value : 32'h70cc702d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf4, value : 32'h70cd70ed},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf5, value : 32'h706d704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf6, value : 32'h20a8708d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf7, value : 32'h20150101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf8, value : 32'h906023c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bf9, value : 32'h87b9001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bfa, value : 32'h631d00e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bfb, value : 32'h6b014873},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bfc, value : 32'h7d0c73c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bfd, value : 32'h462340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bfe, value : 32'h21007034},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54bff, value : 32'h20da1349},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c00, value : 32'h20d503c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c01, value : 32'hf22d1001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c02, value : 32'h1e10915},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c03, value : 32'h8c07208b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c04, value : 32'h271a780c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c05, value : 32'h621a1003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c06, value : 32'hf0237e75},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c07, value : 32'h83bf20d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c08, value : 32'hdb08023f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c09, value : 32'h8003208b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c0a, value : 32'h262ff213},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c0b, value : 32'hdb07f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c0c, value : 32'h1a323ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c0d, value : 32'h204bf011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c0e, value : 32'hf2078300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c0f, value : 32'h736cb8e3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c10, value : 32'ha123ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c11, value : 32'h781df009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c12, value : 32'h432044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c13, value : 32'hb8e5f005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c14, value : 32'h23ca756c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c15, value : 32'h647c0121},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c16, value : 32'h23157bec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c17, value : 32'h71e510cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c18, value : 32'h300e4b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c19, value : 32'h2905d8c9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c1a, value : 32'h21781180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c1b, value : 32'h71f00003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c1c, value : 32'h767d729d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c1d, value : 32'h26ca7074},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c1e, value : 32'h20ca0081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c1f, value : 32'h71041381},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c20, value : 32'h118d2805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c21, value : 32'hffef0e4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c22, value : 32'he8897e1d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c23, value : 32'hbd2271a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c24, value : 32'h1fc0257c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c25, value : 32'h25ca7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c26, value : 32'h18821fe1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c27, value : 32'h2080239c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c28, value : 32'h18002084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c29, value : 32'h700c2342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c2a, value : 32'h41c3c6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c2b, value : 32'h20216},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c2c, value : 32'he564201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c2d, value : 32'h4321f8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c2e, value : 32'h21741c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c2f, value : 32'he4a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c30, value : 32'hd8c9f8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c31, value : 32'hc6c8730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c32, value : 32'h42c3c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c33, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c34, value : 32'h8a404300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c35, value : 32'h2c1239f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c36, value : 32'h582229f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c37, value : 32'h2232627a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c38, value : 32'h80010f8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c39, value : 32'h714c4e8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c3a, value : 32'he9047a18},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c3b, value : 32'h12012585},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c3c, value : 32'h9ae6a12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c3d, value : 32'h2005f72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c3e, value : 32'h252f008e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c3f, value : 32'h700c0387},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c40, value : 32'hda22762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c41, value : 32'h244a43a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c42, value : 32'h9da0480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c43, value : 32'h70ccf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c44, value : 32'hd907d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c45, value : 32'h706c724c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c46, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c47, value : 32'hf76f09c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c48, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c49, value : 32'hf76f096e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c4a, value : 32'hc6c4712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c4b, value : 32'hb80243e3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c4c, value : 32'hf822005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c4d, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c4e, value : 32'hfe6f0a4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c4f, value : 32'h7b204020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c50, value : 32'h78e0b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c51, value : 32'h4608c2e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c52, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c53, value : 32'h88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c54, value : 32'h72ad7214},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c55, value : 32'h94a4728},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c56, value : 32'h25caf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c57, value : 32'hc321161},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c58, value : 32'h926f74f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c59, value : 32'h819f70f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c5a, value : 32'h700c003f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c5b, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c5c, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c5d, value : 32'h96e70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c5e, value : 32'h70ccf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c5f, value : 32'h752cd809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c60, value : 32'h704cb813},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c61, value : 32'h8238a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c62, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c63, value : 32'hf76f0956},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c64, value : 32'hd80c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c65, value : 32'h42a1d92b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c66, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c67, value : 32'h94645c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c68, value : 32'h70ccf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c69, value : 32'hd92bd80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c6a, value : 32'h706c42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c6b, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c6c, value : 32'hf76f0932},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c6d, value : 32'hef0670cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c6e, value : 32'hd80c6d41},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c6f, value : 32'hf005d92b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c70, value : 32'hd92bd80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c71, value : 32'h706c42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c72, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c73, value : 32'hf76f0916},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c74, value : 32'h708c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c75, value : 32'h4788d92b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c76, value : 32'hbf9242a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c77, value : 32'h40e1726c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c78, value : 32'h90245c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c79, value : 32'h70ccf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c7a, value : 32'hd92bd80c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c7b, value : 32'h726c42a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c7c, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c7d, value : 32'hf76f08ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c7e, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c7f, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c80, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c81, value : 32'h8de70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c82, value : 32'h264af76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c83, value : 32'h7dfb0280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c84, value : 32'h40a1d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c85, value : 32'h706cda10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c86, value : 32'h45c1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c87, value : 32'hf76f08c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c88, value : 32'h2f4170cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c89, value : 32'hd90710c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c8a, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c8b, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c8c, value : 32'hf76f08b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c8d, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c8e, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c8f, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c90, value : 32'h8a270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c91, value : 32'h264af76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c92, value : 32'hb2e0bc0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c93, value : 32'h700cf74f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c94, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c95, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c96, value : 32'h88a70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c97, value : 32'h70ccf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c98, value : 32'h18002555},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c99, value : 32'h704cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c9a, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c9b, value : 32'h87645c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c9c, value : 32'h70ccf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c9d, value : 32'h78e0c6c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c9e, value : 32'hc1a6c3fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54c9f, value : 32'hc045d93b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca0, value : 32'hc86b911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca1, value : 32'h740cf8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca2, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca3, value : 32'h10020150},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca4, value : 32'h42830501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca5, value : 32'h1002b220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca6, value : 32'hb2210501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca7, value : 32'h5011002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca8, value : 32'h1002b222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ca9, value : 32'hb2230501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54caa, value : 32'h5011002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cab, value : 32'h9020b224},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cac, value : 32'h9021b225},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cad, value : 32'h9022b226},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cae, value : 32'h808010d7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54caf, value : 32'he805b227},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb0, value : 32'h30961210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb1, value : 32'h120ff003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb2, value : 32'h700e3096},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb3, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb4, value : 32'hc0441230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb5, value : 32'h1f07216},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb6, value : 32'h702c0026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb7, value : 32'h20510811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb8, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cb9, value : 32'h3f8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cba, value : 32'hf2e97014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cbb, value : 32'h2800710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cbc, value : 32'hd960400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cbd, value : 32'h780ff96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cbe, value : 32'h702ec005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cbf, value : 32'hf29c7014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc0, value : 32'h202fc704},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc1, value : 32'hc0803407},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc2, value : 32'h4402015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc3, value : 32'h40020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc4, value : 32'hf6ef0f8e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc5, value : 32'ha6e68b2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc6, value : 32'h78b0f76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc7, value : 32'h70ad45f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc8, value : 32'h10875d2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cc9, value : 32'h704e0026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cca, value : 32'h3540210a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ccb, value : 32'hbf7706e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ccc, value : 32'h11012095},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ccd, value : 32'h740c3494},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cce, value : 32'h1f8e2532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ccf, value : 32'h4788000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd0, value : 32'h41c34222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd1, value : 32'h50077},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd2, value : 32'h240a4362},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd3, value : 32'h45c10400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd4, value : 32'hf8ef0bb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd5, value : 32'h500260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd6, value : 32'h13310e1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd7, value : 32'h3083120e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd8, value : 32'h407202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cd9, value : 32'hfb6f0a86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cda, value : 32'h487212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cdb, value : 32'hda22e803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cdc, value : 32'h6b09f00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cdd, value : 32'h2538da22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cde, value : 32'h23781001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cdf, value : 32'h20052000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce0, value : 32'h7ac0807e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce1, value : 32'h4382710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce2, value : 32'h4c02800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce3, value : 32'h683244c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce4, value : 32'h782570cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce5, value : 32'h272f762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce6, value : 32'h700c2007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce7, value : 32'hf72f0f46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce8, value : 32'h5c0250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ce9, value : 32'h13310e79},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cea, value : 32'h1487262f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ceb, value : 32'ha3e4003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cec, value : 32'h41c1fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ced, value : 32'h244fe823},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cee, value : 32'h740c21d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cef, value : 32'h41c34222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf0, value : 32'h50078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf1, value : 32'h240a4362},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf2, value : 32'h254a0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf3, value : 32'hb3a0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf4, value : 32'h260af8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf5, value : 32'hb130500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf6, value : 32'h704c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf7, value : 32'h7704ca0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf8, value : 32'h10000d07},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cf9, value : 32'h700cda22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cfa, value : 32'h4382762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cfb, value : 32'h300244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cfc, value : 32'h5c0250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cfd, value : 32'hf72f0eee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cfe, value : 32'h400370cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54cff, value : 32'hfb6f09ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d00, value : 32'he88e41c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d01, value : 32'h742c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d02, value : 32'hf76f09ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d03, value : 32'hb11704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d04, value : 32'h700c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d05, value : 32'h9c2702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d06, value : 32'h704cf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d07, value : 32'h71667146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d08, value : 32'h74a6f187},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d09, value : 32'hf17e71a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d0a, value : 32'h74367126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d0b, value : 32'hffe506da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d0c, value : 32'hf045e72c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d0d, value : 32'h704e740f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d0e, value : 32'h72eec080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d0f, value : 32'h4802015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d10, value : 32'h70ad70ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d11, value : 32'h40020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d12, value : 32'h2005781b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d13, value : 32'h40f93},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d14, value : 32'he4d1000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d15, value : 32'h240a2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d16, value : 32'h25002580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d17, value : 32'h80002f95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d18, value : 32'h70ed1230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d19, value : 32'h2b00225a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d1a, value : 32'h1f822732},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d1b, value : 32'h4788000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d1c, value : 32'h7941c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d1d, value : 32'h78f50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d1e, value : 32'h4002014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d1f, value : 32'h200e2532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d20, value : 32'ha86740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d21, value : 32'h43c1f8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d22, value : 32'h71e578af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d23, value : 32'h71a57062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d24, value : 32'hb89cb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d25, value : 32'h248db89f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d26, value : 32'ha0c02a3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d27, value : 32'h26ff278d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d28, value : 32'hd1571ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d29, value : 32'h78af103e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d2a, value : 32'hb8027062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d2b, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d2c, value : 32'h4441800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d2d, value : 32'h30bf208d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d2e, value : 32'hc0047146},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d2f, value : 32'h72047106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d30, value : 32'hf10ac044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d31, value : 32'h901c40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d32, value : 32'hb02001f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d33, value : 32'h804418f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d34, value : 32'h78e0c7da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d35, value : 32'h716ec2f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d36, value : 32'h23064010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d37, value : 32'h16002013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d38, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d39, value : 32'h70140131},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d3a, value : 32'h2740224a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d3b, value : 32'h2100240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d3c, value : 32'h46504570},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d3d, value : 32'hdaa4628},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d3e, value : 32'h22caf6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d3f, value : 32'h70ad25a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d40, value : 32'h11c7552},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d41, value : 32'h40a20026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d42, value : 32'h1f912532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d43, value : 32'h6208000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d44, value : 32'hc8a4122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d45, value : 32'h2632faef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d46, value : 32'h8bd144f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d47, value : 32'hd1b0010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d48, value : 32'h700c1131},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d49, value : 32'h744cd910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d4a, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d4b, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d4c, value : 32'hf72f0db2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d4d, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d4e, value : 32'h704c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d4f, value : 32'h240a43e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d50, value : 32'h250a0440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d51, value : 32'hd9e0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d52, value : 32'h70ccf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d53, value : 32'hd922700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d54, value : 32'hf76f0886},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d55, value : 32'hd85704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d56, value : 32'he191755},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d57, value : 32'h1f08734e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d58, value : 32'h16000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d59, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d5a, value : 32'h85d00ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d5b, value : 32'hf034001f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d5c, value : 32'h734f0e55},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d5d, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d5e, value : 32'h14110d61},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d5f, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d60, value : 32'h8820122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d61, value : 32'h203c8803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d62, value : 32'h8620040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d63, value : 32'h4162fb6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d64, value : 32'ha32e81a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d65, value : 32'hd8fafbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d66, value : 32'h700c7910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d67, value : 32'hf76f083a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d68, value : 32'h274f704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d69, value : 32'h700c11c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d6a, value : 32'h704c762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d6b, value : 32'h440240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d6c, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d6d, value : 32'hf72f0d2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d6e, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d6f, value : 32'h81ad922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d70, value : 32'h704cf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d71, value : 32'h9fed8fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d72, value : 32'h7910fbcf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d73, value : 32'h80a700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d74, value : 32'h704cf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d75, value : 32'hf19671a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d76, value : 32'hc41edfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d77, value : 32'h8e012010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d78, value : 32'hdf080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d79, value : 32'h20538e14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d7a, value : 32'hf21880fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d7b, value : 32'hca6700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d7c, value : 32'h712cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d7d, value : 32'hf6cf0caa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d7e, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d7f, value : 32'h9963a98},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d80, value : 32'hd908fc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d81, value : 32'hfe6f0cda},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d82, value : 32'h40c340c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d83, value : 32'hd400003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d84, value : 32'hfc6f0982},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d85, value : 32'hf1e0d908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d86, value : 32'hf1d7d8c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d87, value : 32'hd941700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d88, value : 32'hf72f0fb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d89, value : 32'h700c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d8a, value : 32'hf72f0c6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d8b, value : 32'he41712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d8c, value : 32'h8e1c2010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d8d, value : 32'h15e0831},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d8e, value : 32'hf6cf0c66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d8f, value : 32'h20452053},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d90, value : 32'hd919d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d91, value : 32'hdb85744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d92, value : 32'hc9a708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d93, value : 32'h70ccf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d94, value : 32'hc42700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d95, value : 32'h712cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d96, value : 32'h5b40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d97, value : 32'h9368d80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d98, value : 32'h702cfc6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d99, value : 32'he56700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d9a, value : 32'h4102f8ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d9b, value : 32'h78e0c6d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d9c, value : 32'h716ec2f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d9d, value : 32'h23064010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d9e, value : 32'h16002013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54d9f, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da0, value : 32'h70140131},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da1, value : 32'h2740224a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da2, value : 32'h2140240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da3, value : 32'h2100250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da4, value : 32'h47504670},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da5, value : 32'h8664628},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da6, value : 32'h22caf9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da7, value : 32'hc0225a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da8, value : 32'haeef6cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54da9, value : 32'h70adfe4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54daa, value : 32'h12a7552},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dab, value : 32'h40c20026},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dac, value : 32'h1f912532},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dad, value : 32'h6208000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dae, value : 32'hae24122},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54daf, value : 32'h2632faef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db0, value : 32'h7014144f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db1, value : 32'hd11f285},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db2, value : 32'h700c2030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db3, value : 32'hf0ad91e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db4, value : 32'h714cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db5, value : 32'h11310d55},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db6, value : 32'h762c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db7, value : 32'hf72f0efa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db8, value : 32'h700c714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54db9, value : 32'h704cd92c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dba, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dbb, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dbc, value : 32'hf72f0bf2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dbd, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dbe, value : 32'h704cd92d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dbf, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc0, value : 32'h400250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc1, value : 32'hf72f0bde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc2, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc3, value : 32'heca762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc4, value : 32'h714cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc5, value : 32'h41e14022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc6, value : 32'hf72f0f9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc7, value : 32'h25424202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc8, value : 32'h8451600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dc9, value : 32'hf0500154},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dca, value : 32'h41e14022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dcb, value : 32'hf72f0f8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dcc, value : 32'hed234202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dcd, value : 32'h14d00d31},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dce, value : 32'h94110de7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dcf, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd0, value : 32'h8820122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd1, value : 32'h203c8803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd2, value : 32'hea20040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd3, value : 32'h4162fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd4, value : 32'h700ce867},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd5, value : 32'he82762c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd6, value : 32'h714cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd7, value : 32'h11c1274f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd8, value : 32'hf1dc4022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dd9, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dda, value : 32'hca8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ddb, value : 32'h3e0859},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ddc, value : 32'hd91e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ddd, value : 32'hc47f025},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dde, value : 32'h8e012010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ddf, value : 32'hdf080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de0, value : 32'h20538e14},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de1, value : 32'hf21b80fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de2, value : 32'hfe4f09e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de3, value : 32'hb06700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de4, value : 32'h712cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de5, value : 32'hf6cf0b0a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de6, value : 32'hfe4f09f6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de7, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de8, value : 32'hff23a98},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54de9, value : 32'hd908fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dea, value : 32'hfe6f0b36},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54deb, value : 32'h40c340c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dec, value : 32'hd400003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ded, value : 32'hfc2f0fde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dee, value : 32'h700cd908},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54def, value : 32'he1ad918},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df0, value : 32'h714cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df1, value : 32'h762c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df2, value : 32'hf72f0e0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df3, value : 32'h71a5714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df4, value : 32'h99af16c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df5, value : 32'h700cfe4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df6, value : 32'hf72f0aba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df7, value : 32'hf5b712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df8, value : 32'h8e1c2010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54df9, value : 32'h15e084b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dfa, value : 32'hf6cf0ab6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dfb, value : 32'hfe4f09a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dfc, value : 32'hd925700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dfd, value : 32'hdb85704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dfe, value : 32'h250a708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54dff, value : 32'hae60400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e00, value : 32'h70ccf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e01, value : 32'hd926700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e02, value : 32'hdb85704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e03, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e04, value : 32'hf72f0ad2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e05, value : 32'h95670cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e06, value : 32'h700cfe4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e07, value : 32'hf72f0a76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e08, value : 32'h40c3712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e09, value : 32'h8d80005b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e0a, value : 32'hfc2f0f6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e0b, value : 32'h710c702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e0c, value : 32'hf8ef0c8a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e0d, value : 32'he5e4102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e0e, value : 32'hc6d6f98f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e0f, value : 32'h2132c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e10, value : 32'h47680091},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e11, value : 32'h46284548},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e12, value : 32'hf6ef0a56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e13, value : 32'hf0f4010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e14, value : 32'heaa105f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e15, value : 32'h93af94f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e16, value : 32'h66a9fe4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e17, value : 32'he5a40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e18, value : 32'h4202f72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e19, value : 32'h13802542},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e1a, value : 32'hb50819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e1b, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e1c, value : 32'h706cda20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e1d, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e1e, value : 32'hf72f0a6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e1f, value : 32'hf01f70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e20, value : 32'h14310d3b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e21, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e22, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e23, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e24, value : 32'hf72f0a52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e25, value : 32'h93971cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e26, value : 32'h700c217e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e27, value : 32'hfacf082a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e28, value : 32'hfe4f08ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e29, value : 32'h9ee700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e2a, value : 32'h702cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e2b, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e2c, value : 32'hee21388},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e2d, value : 32'hd914fc2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e2e, value : 32'h700cf010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e2f, value : 32'h764cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e30, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e31, value : 32'ha1e70ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e32, value : 32'h70ccf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e33, value : 32'hfe4f089e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e34, value : 32'h9c2700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e35, value : 32'h712cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e36, value : 32'hdb8bfe0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e37, value : 32'hc6caf981},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e38, value : 32'h47cbc2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e39, value : 32'h2fe8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e3a, value : 32'h10911700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e3b, value : 32'hf92f0f9a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e3c, value : 32'h40c3730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e3d, value : 32'h11408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e3e, value : 32'he80b8800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e3f, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e40, value : 32'h18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e41, value : 32'h2002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e42, value : 32'h2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e43, value : 32'h700cf002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e44, value : 32'hcd6d987},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e45, value : 32'hb910f66f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e46, value : 32'h207e090b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e47, value : 32'hcbed820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e48, value : 32'hddaff8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e49, value : 32'h8fa1f94f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e4a, value : 32'h10901700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e4b, value : 32'hf6ef0972},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e4c, value : 32'h10022589},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e4d, value : 32'hfe4f085a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e4e, value : 32'h70cded1b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e4f, value : 32'h1f802600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e50, value : 32'h3808000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e51, value : 32'hda0f8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e52, value : 32'hf72f0d6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e53, value : 32'h80801080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e54, value : 32'h762c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e55, value : 32'hf72f0c82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e56, value : 32'h258d714c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e57, value : 32'h71c51cbf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e58, value : 32'hfe4f080a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e59, value : 32'h92e700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e5a, value : 32'h712cf72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e5b, value : 32'hffef003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e5c, value : 32'h80ffe0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e5d, value : 32'hd822207e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e5e, value : 32'hff8f0c62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e5f, value : 32'hd16f1d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e60, value : 32'h90df98f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e61, value : 32'hd821207e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e62, value : 32'hff8f0c52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e63, value : 32'h78e0c6ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e64, value : 32'h43c3c5e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e65, value : 32'h46a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e66, value : 32'h93034008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e67, value : 32'hf042242f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e68, value : 32'h7a1df215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e69, value : 32'h2200706d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e6a, value : 32'h40f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e6b, value : 32'h20a81000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e6c, value : 32'h201503c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e6d, value : 32'h716512c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e6e, value : 32'h924192a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e6f, value : 32'h7d45ba10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e70, value : 32'hba9c6c52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e71, value : 32'hba9f7185},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e72, value : 32'h6038a2a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e73, value : 32'h9300b303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e74, value : 32'hb3006038},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e75, value : 32'h78e0c4c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e76, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e77, value : 32'h4710b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e78, value : 32'hb89fd840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e79, value : 32'h2100240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e7a, value : 32'h45504378},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e7b, value : 32'h991000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e7c, value : 32'h10e54630},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e7d, value : 32'h700e8098},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e7e, value : 32'h716e724e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e7f, value : 32'h24002b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e80, value : 32'h2004722e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e81, value : 32'hb80206cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e82, value : 32'h40e200f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e83, value : 32'h70ad4003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e84, value : 32'hf23078eb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e85, value : 32'h23402b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e86, value : 32'hf92f0e6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e87, value : 32'h40c3780f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e88, value : 32'h11408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e89, value : 32'he8188800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e8a, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e8b, value : 32'h18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e8c, value : 32'hff0825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e8d, value : 32'h259f4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e8e, value : 32'h209f1582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e8f, value : 32'h42c202c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e90, value : 32'h708c43a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e91, value : 32'h500250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e92, value : 32'h651975e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e93, value : 32'hffef0c26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e94, value : 32'hf01078cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e95, value : 32'h259f4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e96, value : 32'h209f1582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e97, value : 32'h42c202c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e98, value : 32'h240a43a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e99, value : 32'h75e20500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e9a, value : 32'ha6e6519},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e9b, value : 32'h78cfffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e9c, value : 32'h218d4023},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e9d, value : 32'h71ad243f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e9e, value : 32'h20bf228d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54e9f, value : 32'he0a710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea0, value : 32'h730cf92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea1, value : 32'h341b1404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea2, value : 32'h78e0c6da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea3, value : 32'h4568c3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea4, value : 32'h47284648},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea5, value : 32'hb0091cf8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea6, value : 32'h30011c04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea7, value : 32'h30c21c01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea8, value : 32'hf72f0ae2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ea9, value : 32'h2578c360},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eaa, value : 32'h41c11000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eab, value : 32'h6841781b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eac, value : 32'hf72f0a86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ead, value : 32'hacec080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eae, value : 32'h40e1f72f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eaf, value : 32'hfd6700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb0, value : 32'h712cf6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb1, value : 32'h78e0c7c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb2, value : 32'h2945c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb3, value : 32'h4608018b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb4, value : 32'hd3d70ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb5, value : 32'h8e0112c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb6, value : 32'h8e228e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb7, value : 32'h7a05b808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb8, value : 32'hb8088e03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eb9, value : 32'hb8107825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eba, value : 32'h812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ebb, value : 32'h8e448e05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ebc, value : 32'hb8087734},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ebd, value : 32'hf2077845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ebe, value : 32'hb99cb902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ebf, value : 32'hb100b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec0, value : 32'hc06f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec1, value : 32'h76c5fc0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec2, value : 32'hf1e571a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec3, value : 32'h78e0c6c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec4, value : 32'h7034c2e4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec5, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec6, value : 32'hf22712e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec7, value : 32'hc1110a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec8, value : 32'h7180244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ec9, value : 32'h7b31c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eca, value : 32'h2144b923},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ecb, value : 32'h68520401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ecc, value : 32'h22057965},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ecd, value : 32'h90030f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ece, value : 32'h7b2fd580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ecf, value : 32'hf812205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed0, value : 32'hd5849003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed1, value : 32'h800042c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed2, value : 32'hb4600550},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed3, value : 32'h20a8b160},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed4, value : 32'h12100300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed5, value : 32'h79050401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed6, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed7, value : 32'h90030f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed8, value : 32'hb160c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ed9, value : 32'h2042f017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eda, value : 32'hf215803c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54edb, value : 32'h20a86944},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54edc, value : 32'h120604c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54edd, value : 32'hb8020400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ede, value : 32'hf832005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54edf, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee0, value : 32'h4c0120e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee1, value : 32'hb8237911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee2, value : 32'h4002044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee3, value : 32'h780f7825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee4, value : 32'h720cb300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee5, value : 32'h900345cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee6, value : 32'h46cbd478},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee7, value : 32'hf07c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee8, value : 32'h10c51d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ee9, value : 32'hfc2f0b62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eea, value : 32'h10c51e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eeb, value : 32'h900f41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eec, value : 32'h2150e008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eed, value : 32'h710c04c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eee, value : 32'h1451900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eef, value : 32'h1451a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef0, value : 32'hb200b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef1, value : 32'hb600b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef2, value : 32'h78e0c6c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef3, value : 32'h42c3c0e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef4, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef5, value : 32'h40288a81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef6, value : 32'hc518aa0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef7, value : 32'h43001364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef8, value : 32'h22479},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ef9, value : 32'he20970b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54efa, value : 32'h22cac809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54efb, value : 32'h20050062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54efc, value : 32'h221f00ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54efd, value : 32'h2d40034b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54efe, value : 32'h240a130f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54eff, value : 32'h7fc57080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f00, value : 32'h20a8706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f01, value : 32'h2b400440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f02, value : 32'h70b40200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f03, value : 32'h20f478c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f04, value : 32'h78e512c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f05, value : 32'hb8027164},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f06, value : 32'hb8927165},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f07, value : 32'hb89fb89c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f08, value : 32'h7591b020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f09, value : 32'hf7a971a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f0a, value : 32'h78e0c4c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f0b, value : 32'h4010c2e8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f0c, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f0d, value : 32'h47cb122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f0e, value : 32'h4db48001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f0f, value : 32'h2754e903},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f10, value : 32'h8ea01f0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f11, value : 32'h8578e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f12, value : 32'hd8c80364},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f13, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f14, value : 32'h880012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f15, value : 32'h36e0843},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f16, value : 32'heca79af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f17, value : 32'h4002fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f18, value : 32'hc8094408},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f19, value : 32'h13822d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f1a, value : 32'h7280244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f1b, value : 32'h700c6832},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f1c, value : 32'h20a87a25},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f1d, value : 32'hc2104c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f1e, value : 32'h255a100e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f1f, value : 32'h61f91501},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f20, value : 32'h321f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f21, value : 32'h2812840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f22, value : 32'h21057945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f23, value : 32'h90040f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f24, value : 32'hb1600320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f25, value : 32'h71a57104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f26, value : 32'had2f1d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f27, value : 32'hc6c8fc0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f28, value : 32'h718ec2f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f29, value : 32'h2c004610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f2a, value : 32'h16002040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f2b, value : 32'h80007093},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f2c, value : 32'hb8020004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f2d, value : 32'h200f4230},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f2e, value : 32'haaf0051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f2f, value : 32'h235302f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f30, value : 32'he28a20d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f31, value : 32'h700ef4b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f32, value : 32'h81372ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f33, value : 32'h16002010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f34, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f35, value : 32'h8890040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f36, value : 32'h272f0010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f37, value : 32'h40421400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f38, value : 32'hfaaf0c42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f39, value : 32'h260041e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f3a, value : 32'h42c323c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f3b, value : 32'hea48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f3c, value : 32'h89218960},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f3d, value : 32'h6149634d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f3e, value : 32'h6914e804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f3f, value : 32'hf0047d05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f40, value : 32'h7d25bd04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f41, value : 32'h2800710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f42, value : 32'hb7e0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f43, value : 32'h780ff92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f44, value : 32'h750c7eaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f45, value : 32'h41c34242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f46, value : 32'h301d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f47, value : 32'h9ea4302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f48, value : 32'h44c1f8af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f49, value : 32'h447212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f4a, value : 32'hfe2f0a2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f4b, value : 32'h235f40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f4c, value : 32'h60f82b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f4d, value : 32'h70c37042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f4e, value : 32'h12448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f4f, value : 32'h20300a15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f50, value : 32'hcc7a8a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f51, value : 32'h1e002010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f52, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f53, value : 32'hf008017e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f54, value : 32'h20100ccb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f55, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f56, value : 32'h17d8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f57, value : 32'h258d710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f58, value : 32'h708e2dfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f59, value : 32'h700ef064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f5a, value : 32'h81372ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f5b, value : 32'h16002010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f5c, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f5d, value : 32'h8890040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f5e, value : 32'h272f0010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f5f, value : 32'h40421400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f60, value : 32'hfaaf0ba2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f61, value : 32'h260041e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f62, value : 32'h42c323c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f63, value : 32'hea48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f64, value : 32'h89218960},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f65, value : 32'h6149634d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f66, value : 32'h6914e804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f67, value : 32'hf0047d05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f68, value : 32'h7d25bd04},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f69, value : 32'h2800710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f6a, value : 32'hade0400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f6b, value : 32'h780ff92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f6c, value : 32'h750c7eaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f6d, value : 32'h41c34242},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f6e, value : 32'h301d6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f6f, value : 32'h94a4302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f70, value : 32'h44c1f8af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f71, value : 32'h447212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f72, value : 32'hfe2f0822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f73, value : 32'h235f40c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f74, value : 32'h60f82b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f75, value : 32'h70c37042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f76, value : 32'h12408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f77, value : 32'h20300a15},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f78, value : 32'hc31a8a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f79, value : 32'h1e002010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f7a, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f7b, value : 32'hf00800f7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f7c, value : 32'h20100c35},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f7d, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f7e, value : 32'hf28000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f7f, value : 32'h258d710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f80, value : 32'h708e2dfe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f81, value : 32'h1e00f014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f82, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f83, value : 32'hf0100180},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f84, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f85, value : 32'h1018000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f86, value : 32'h1e00f00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f87, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f88, value : 32'hf006017f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f89, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f8a, value : 32'hfc8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f8b, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f8c, value : 32'h408000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f8d, value : 32'h730ce803},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f8e, value : 32'h710cf002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f8f, value : 32'hf90f0a4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f90, value : 32'h78e0c6d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f91, value : 32'hc1a8c3e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f92, value : 32'h1243276f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f93, value : 32'h800145cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f94, value : 32'h8fc04e7c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f95, value : 32'h1756712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f96, value : 32'h20441080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f97, value : 32'hbaa0202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f98, value : 32'h40a1fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f99, value : 32'hd91440a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f9a, value : 32'hf72f0cb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f9b, value : 32'h178a704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f9c, value : 32'h40a11082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f9d, value : 32'hb92bac3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f9e, value : 32'hd914fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54f9f, value : 32'hf92f09fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa0, value : 32'hab6c084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa1, value : 32'hc080fe2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa2, value : 32'hb0ac080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa3, value : 32'hd910f92f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa4, value : 32'h8358f17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa5, value : 32'h40c3001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa6, value : 32'h12e08000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa7, value : 32'he8148800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa8, value : 32'h41c3bec3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fa9, value : 32'h12308000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54faa, value : 32'h1b00265f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fab, value : 32'h6119602a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fac, value : 32'h1da28902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fad, value : 32'h89011002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fae, value : 32'h10021d57},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54faf, value : 32'had4c8903},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb0, value : 32'h10021ded},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb1, value : 32'hd91040a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb2, value : 32'hf72f0c52},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb3, value : 32'h40a1dafb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb4, value : 32'hb36d910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb5, value : 32'hda41fbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb6, value : 32'h702c40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb7, value : 32'hdbffc284},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb8, value : 32'hffef0afa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fb9, value : 32'h40a1708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fba, value : 32'hb1ed910},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fbb, value : 32'h744cfbaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fbc, value : 32'h702c40a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fbd, value : 32'h8c6c280},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fbe, value : 32'h716cf76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fbf, value : 32'h78e0c7c6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc0, value : 32'h78e07ee0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc1, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc2, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc3, value : 32'h46303604},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc4, value : 32'hc3a702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc5, value : 32'h4318f7ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc6, value : 32'h451071ad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc7, value : 32'h16c02d00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc8, value : 32'hfa2f0992},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fc9, value : 32'h99a68f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fca, value : 32'h4210fa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fcb, value : 32'h8e82208c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fcc, value : 32'h238a70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fcd, value : 32'hf7062f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fce, value : 32'hfa0f0986},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fcf, value : 32'h8932054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd0, value : 32'h70831600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd1, value : 32'h48000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd2, value : 32'h750cbbc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd3, value : 32'h41c34263},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd4, value : 32'h20409},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd5, value : 32'hf86f0fb2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd6, value : 32'h16d0270f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd7, value : 32'h41c3d82e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd8, value : 32'he010001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fd9, value : 32'hb70f478b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fda, value : 32'hb709d895},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fdb, value : 32'hb890d897},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fdc, value : 32'h41c3c155},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fdd, value : 32'h12a0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fde, value : 32'h2154c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fdf, value : 32'hb86c0942},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe0, value : 32'hc043c149},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe1, value : 32'hc809e115},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe2, value : 32'hc2466989},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe3, value : 32'h422005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe4, value : 32'h7224b755},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe5, value : 32'hba30c24f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe6, value : 32'hb7567905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe7, value : 32'hc14c6c49},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe8, value : 32'h812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fe9, value : 32'h3032005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fea, value : 32'h30441c42},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54feb, value : 32'h1c44b930},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fec, value : 32'h6a2e3044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fed, value : 32'h20057905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fee, value : 32'h10f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fef, value : 32'hb73b00fb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff0, value : 32'hb703b930},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff1, value : 32'hb73cb830},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff2, value : 32'hb704d90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff3, value : 32'h714cc080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff4, value : 32'h31c51c50},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff5, value : 32'h33441c4e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff6, value : 32'hb7aab7b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff7, value : 32'h1c58b7c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff8, value : 32'h1c523384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ff9, value : 32'h1c4c3384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ffa, value : 32'h1c463384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ffb, value : 32'h1c403384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ffc, value : 32'hb7dd3384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ffd, value : 32'hb7d7b7da},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54ffe, value : 32'hb7d1b7d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h54fff, value : 32'hb7cbb7ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55000, value : 32'hb7c5b7c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55001, value : 32'hfdef0af6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55002, value : 32'h1600c352},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55003, value : 32'h80007083},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55004, value : 32'h245512e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55005, value : 32'h244a3801},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55006, value : 32'h700c7200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55007, value : 32'h33801c8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55008, value : 32'h33801c88},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55009, value : 32'h33801c84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5500a, value : 32'h33801c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5500b, value : 32'h40020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5500c, value : 32'hb137a1d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5500d, value : 32'h2605008e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5500e, value : 32'h90381f82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5500f, value : 32'h9240012c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55010, value : 32'h7224b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55011, value : 32'h76c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55012, value : 32'h71044000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55013, value : 32'h1643276f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55014, value : 32'h20448f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55015, value : 32'hf2068202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55016, value : 32'h70851e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55017, value : 32'hc3789007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55018, value : 32'h41c3700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55019, value : 32'hc25c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5501a, value : 32'h800046cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5501b, value : 32'h1e00122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5501c, value : 32'h901c7004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5501d, value : 32'h1e000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5501e, value : 32'h90077004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5501f, value : 32'hb100f804},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55020, value : 32'h1964ea99},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55021, value : 32'hd9400205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55022, value : 32'h900740c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55023, value : 32'hb020c2c4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55024, value : 32'h8e41b0a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55025, value : 32'ha778e20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55026, value : 32'h7a5b0064},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55027, value : 32'h70402614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55028, value : 32'h48c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55029, value : 32'h412217},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5502a, value : 32'h8566942},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5502b, value : 32'h702cf62f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5502c, value : 32'h1600f02d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5502d, value : 32'h80007082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5502e, value : 32'h72540008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5502f, value : 32'h901c43c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55030, value : 32'h42c30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55031, value : 32'hf8009007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55032, value : 32'h1964f406},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55033, value : 32'hb3000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55034, value : 32'hf006b200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55035, value : 32'h1051964},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55036, value : 32'hb2a0b3a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55037, value : 32'h8e008e21},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55038, value : 32'h24092b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55039, value : 32'h71247902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5503a, value : 32'h7040240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5503b, value : 32'h3c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5503c, value : 32'h6812000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5503d, value : 32'h70022614},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5503e, value : 32'h48c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5503f, value : 32'h811120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55040, value : 32'h21787104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55041, value : 32'hb9080001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55042, value : 32'hd8aab220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55043, value : 32'h70041e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55044, value : 32'hc0b89007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55045, value : 32'hf68f098a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55046, value : 32'h407202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55047, value : 32'hc057d907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55048, value : 32'h145cd841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55049, value : 32'hb8133005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5504a, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5504b, value : 32'h9b6708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5504c, value : 32'h70ccf6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5504d, value : 32'hd907700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5504e, value : 32'h706cda08},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5504f, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55050, value : 32'hf6ef09a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55051, value : 32'h145c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55052, value : 32'hd8803005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55053, value : 32'hd907b893},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55054, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55055, value : 32'h98e708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55056, value : 32'h70ccf6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55057, value : 32'h936700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55058, value : 32'h712cf6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55059, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5505a, value : 32'he2a1388},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5505b, value : 32'h752cfbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5505c, value : 32'hd9ff710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5505d, value : 32'hfb6f0b7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5505e, value : 32'h216f704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5505f, value : 32'h40d32443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55060, value : 32'h48c8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55061, value : 32'h20801100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55062, value : 32'h1012078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55063, value : 32'h7424b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55064, value : 32'h180ab806},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55065, value : 32'h20892042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55066, value : 32'h41c30e43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55067, value : 32'h103df},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55068, value : 32'h740c6846},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55069, value : 32'hf86f0d62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5506a, value : 32'h20841808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5506b, value : 32'h6872c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5506c, value : 32'h901c40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5506d, value : 32'h23050504},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5506e, value : 32'hb1a00001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5506f, value : 32'hf812305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55070, value : 32'h4fc901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55071, value : 32'h834418a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55072, value : 32'hf802305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55073, value : 32'h4dc901c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55074, value : 32'h11009000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55075, value : 32'ha1b2082},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55076, value : 32'hb8c500b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55077, value : 32'h2c2204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55078, value : 32'h8f20b140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55079, value : 32'hfe0925},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5507a, value : 32'h301204f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5507b, value : 32'h204ff009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5507c, value : 32'hb1400302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5507d, value : 32'h9158f20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5507e, value : 32'h204f00fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5507f, value : 32'h23050341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55080, value : 32'h901c0f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55081, value : 32'hb02004f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55082, value : 32'hf802305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55083, value : 32'hc3ec9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55084, value : 32'h71051e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55085, value : 32'hc12c903b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55086, value : 32'hafeb0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55087, value : 32'h710cfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55088, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55089, value : 32'hf812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5508a, value : 32'h949004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5508b, value : 32'h1c909120},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5508c, value : 32'h8f203040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5508d, value : 32'hde091b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5508e, value : 32'hf812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5508f, value : 32'hc0949007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55090, value : 32'h30001490},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55091, value : 32'h80206c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55092, value : 32'hc02045},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55093, value : 32'h1600b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55094, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55095, value : 32'h22440126},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55096, value : 32'hb8e22051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55097, value : 32'hf9e20850},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55098, value : 32'h21004063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55099, value : 32'h42d32491},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5509a, value : 32'hfb88000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5509b, value : 32'h3a402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5509c, value : 32'h28012240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5509d, value : 32'he72da72},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5509e, value : 32'h2344f5ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5509f, value : 32'h40c32054},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a0, value : 32'hf0a70000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a1, value : 32'h30041c66},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a2, value : 32'h140c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a3, value : 32'hc058ff74},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a4, value : 32'h4208a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a5, value : 32'h30041c6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a6, value : 32'h100ad972},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a7, value : 32'h1c682080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a8, value : 32'hb8063344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a9, value : 32'h30041c64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550aa, value : 32'hffef0822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ab, value : 32'h3a402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ac, value : 32'h204b8f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ad, value : 32'hf4068e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ae, value : 32'h812c098},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550af, value : 32'hd90cffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b0, value : 32'hd90fd80f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b1, value : 32'h24cd2400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b2, value : 32'hf7af091e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b3, value : 32'h27912140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b4, value : 32'h204b8f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b5, value : 32'hf4088e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b6, value : 32'hf88f090a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b7, value : 32'hdee4063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b8, value : 32'h712cff6f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550b9, value : 32'h78afc217},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ba, value : 32'h447212f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550bb, value : 32'hfb2f0dd2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550bc, value : 32'h8f404118},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550bd, value : 32'h8e00224b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550be, value : 32'ha69f20b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550bf, value : 32'h700c00ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c0, value : 32'h41041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c1, value : 32'hae20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c2, value : 32'h271f60f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c3, value : 32'h41c30000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c4, value : 32'h40b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c5, value : 32'hf86f0bf2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c6, value : 32'hd861740c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c7, value : 32'h900745cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c8, value : 32'hb808c29c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550c9, value : 32'hb500712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ca, value : 32'hf6af0f6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550cb, value : 32'h208ad808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550cc, value : 32'h41c30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550cd, value : 32'h40c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ce, value : 32'hbceb500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550cf, value : 32'h740cf86f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d0, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d1, value : 32'h18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d2, value : 32'h1fcb8e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d3, value : 32'hdd0a0022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d4, value : 32'h21001008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d5, value : 32'hf6af0f3e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d6, value : 32'h258c712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d7, value : 32'hf0f91f3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d8, value : 32'h40d41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550d9, value : 32'hba20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550da, value : 32'h740cf86f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550db, value : 32'hf26710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550dc, value : 32'h712cf6af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550dd, value : 32'h3a402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550de, value : 32'hd6e4142},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550df, value : 32'hda10f5ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e0, value : 32'h39402455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e1, value : 32'h24012240},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e2, value : 32'hf5ef0d5e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e3, value : 32'h700cda10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e4, value : 32'hc05f8e20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e5, value : 32'hc05dc05e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e6, value : 32'h8e01c05c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e7, value : 32'h64082d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e8, value : 32'h68417822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550e9, value : 32'h240ac809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ea, value : 32'h68727080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550eb, value : 32'h38020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ec, value : 32'h3802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ed, value : 32'h7865c298},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ee, value : 32'h20057a35},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ef, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f0, value : 32'h900000a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f1, value : 32'ha2007124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f2, value : 32'heca700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f3, value : 32'h712cf6af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f4, value : 32'h258a8e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f5, value : 32'h8e202001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f6, value : 32'h64082d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f7, value : 32'h68617822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f8, value : 32'h240ac809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550f9, value : 32'h685270c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550fa, value : 32'h38020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550fb, value : 32'h3802940},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550fc, value : 32'h20057845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550fd, value : 32'h90040f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550fe, value : 32'h245500a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h550ff, value : 32'h48203a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55100, value : 32'hb3007124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55101, value : 32'hfd4f0fa2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55102, value : 32'he8a700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55103, value : 32'h712cf6af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55104, value : 32'h8e018ea0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55105, value : 32'h36408d7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55106, value : 32'h13912d40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55107, value : 32'h2105d889},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55108, value : 32'h90042f92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55109, value : 32'h1a0001c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5510a, value : 32'hade2004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5510b, value : 32'hd808fbef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5510c, value : 32'h234020f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5510d, value : 32'h3a532455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5510e, value : 32'h23532315},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5510f, value : 32'h39562455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55110, value : 32'h23562615},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55111, value : 32'h40e41c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55112, value : 32'h42a10005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55113, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55114, value : 32'h24540440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55115, value : 32'h20053e11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55116, value : 32'h90040f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55117, value : 32'h900001cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55118, value : 32'h23512115},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55119, value : 32'h20051a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5511a, value : 32'h582044},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5511b, value : 32'h740c4366},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5511c, value : 32'h20171600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5511d, value : 32'h600260a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5511e, value : 32'h20121100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5511f, value : 32'h5c0240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55120, value : 32'h480250a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55121, value : 32'hf86f0a82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55122, value : 32'h81d4470},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55123, value : 32'ha193011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55124, value : 32'h27402033},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55125, value : 32'h80d2040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55126, value : 32'h714e00f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55127, value : 32'hf00471ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55128, value : 32'h2fbf2f84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55129, value : 32'h3010081b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5512a, value : 32'h20720a17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5512b, value : 32'h20402740},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5512c, value : 32'hf5080b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5512d, value : 32'h77ee774e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5512e, value : 32'h2f84f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5512f, value : 32'ha1b2fbf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55130, value : 32'h20782031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55131, value : 32'h20793000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55132, value : 32'h791b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55133, value : 32'h2142b805},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55134, value : 32'h20420052},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55135, value : 32'h24000417},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55136, value : 32'h1e0025d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55137, value : 32'h190025c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55138, value : 32'h71a52480},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55139, value : 32'h25001b00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5513a, value : 32'h258cf195},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5513b, value : 32'h40632dfd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5513c, value : 32'hf7af0e5a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5513d, value : 32'h885702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5513e, value : 32'h8e210010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5513f, value : 32'h9438e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55140, value : 32'h204000a4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55141, value : 32'hc8090a83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55142, value : 32'h71247942},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55143, value : 32'h7040240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55144, value : 32'h5c020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55145, value : 32'h30c2a40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55146, value : 32'h24057c05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55147, value : 32'hb90210c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55148, value : 32'hf8d2105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55149, value : 32'h9004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5514a, value : 32'h21056c32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5514b, value : 32'h90040f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5514c, value : 32'h942000a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5514d, value : 32'hc198b520},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5514e, value : 32'h71444941},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5514f, value : 32'ha0eb420},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55150, value : 32'hf01cfd0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55151, value : 32'h21001008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55152, value : 32'hf6af0d4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55153, value : 32'h4063712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55154, value : 32'hff6f0b7a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55155, value : 32'h40c2702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55156, value : 32'hd9e702c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55157, value : 32'h724cfd2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55158, value : 32'h2a952540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55159, value : 32'h2005c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5515a, value : 32'h41c20540},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5515b, value : 32'h706c704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5515c, value : 32'he5e708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5515d, value : 32'h71acffaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5515e, value : 32'hfd4f0e2e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5515f, value : 32'h45cb70cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55160, value : 32'hc29c9007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55161, value : 32'h9d24063},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55162, value : 32'hb5c0faef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55163, value : 32'h41141c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55164, value : 32'h9760000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55165, value : 32'h740cf86f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55166, value : 32'h702c700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55167, value : 32'hfb2f0f56},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55168, value : 32'hb5d2704c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55169, value : 32'h8f00b5d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5516a, value : 32'hde081f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5516b, value : 32'hb802c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5516c, value : 32'hf812005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5516d, value : 32'hc0949007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5516e, value : 32'h30001490},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5516f, value : 32'h1e00b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55170, value : 32'h90077384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55171, value : 32'hcdac378},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55172, value : 32'h700cf64f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55173, value : 32'h80a752c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55174, value : 32'h714cf6ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55175, value : 32'hcbe700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55176, value : 32'h712cf6af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55177, value : 32'hfaef0f3a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55178, value : 32'hcbe700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55179, value : 32'h700cf64f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5517a, value : 32'h744cd907},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5517b, value : 32'h708c706c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5517c, value : 32'hcf270ac},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5517d, value : 32'h70ccf6af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5517e, value : 32'h145c708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5517f, value : 32'h40803005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55180, value : 32'hb890732c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55181, value : 32'h28414223},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55182, value : 32'hcda0103},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55183, value : 32'h70ccf6af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55184, value : 32'hd907d880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55185, value : 32'h706c744c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55186, value : 32'h70ac708c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55187, value : 32'hf6af0cc6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55188, value : 32'h700c70cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55189, value : 32'hf6af0c6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5518a, value : 32'h922712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5518b, value : 32'hd7afd0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5518c, value : 32'hc080fd4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5518d, value : 32'hcc6d90f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5518e, value : 32'h704cfdaf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5518f, value : 32'h708c1600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55190, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55191, value : 32'h38012455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55192, value : 32'h7200244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55193, value : 32'h20a8700c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55194, value : 32'h7a1d0440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55195, value : 32'h108e0c11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55196, value : 32'h26059140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55197, value : 32'h90381f83},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55198, value : 32'hb340012c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55199, value : 32'h76c37224},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5519a, value : 32'h40000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5519b, value : 32'h24807104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5519c, value : 32'h14043604},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5519d, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5519e, value : 32'h2482c3f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5519f, value : 32'h228a3102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a0, value : 32'h10822084},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a1, value : 32'h2033070f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a2, value : 32'h250a048e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a3, value : 32'h46702100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a4, value : 32'h43304450},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a5, value : 32'hff6f083a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a6, value : 32'he8084110},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a7, value : 32'h710478cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a8, value : 32'h2049b822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551a9, value : 32'hf0050fce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551aa, value : 32'h10320e45},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ab, value : 32'h2648700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ac, value : 32'h40d11000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ad, value : 32'h780f7104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ae, value : 32'h7000240a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551af, value : 32'h34020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b0, value : 32'h407202f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b1, value : 32'h20002115},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b2, value : 32'h9139020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b3, value : 32'h900103c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b4, value : 32'h10050f0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b5, value : 32'h700e7706},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b6, value : 32'hff6f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b7, value : 32'h7014ff0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b8, value : 32'h206220c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551b9, value : 32'hdd3fe6bf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ba, value : 32'hf01df6c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551bb, value : 32'hd940e6c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551bc, value : 32'h45c96e01},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551bd, value : 32'h4b20ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551be, value : 32'h240a78c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551bf, value : 32'h20a87000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c0, value : 32'h21150300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c1, value : 32'h90202340},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c2, value : 32'h3c50911},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c3, value : 32'hf0d9001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c4, value : 32'h71a51005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c5, value : 32'hf007dd3f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c6, value : 32'hff0f0fb6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c7, value : 32'h25c27014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c8, value : 32'hfae1062},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551c9, value : 32'he809ff0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ca, value : 32'h24802132},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551cb, value : 32'h79026d32},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551cc, value : 32'h4022018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551cd, value : 32'h4dd1f004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ce, value : 32'h14022602},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551cf, value : 32'h7e2f78cf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d0, value : 32'h200c2115},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d1, value : 32'h4f109400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d2, value : 32'h94017b10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d3, value : 32'h7f4f78e2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d4, value : 32'hf7e7810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d5, value : 32'h2009ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d6, value : 32'h701400cd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d7, value : 32'h138e2709},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d8, value : 32'hff2f0f6e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551d9, value : 32'h106225c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551da, value : 32'h40a17014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551db, value : 32'h138125ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551dc, value : 32'h710cf213},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551dd, value : 32'h20300b0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551de, value : 32'h30431c05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551df, value : 32'h704c712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e0, value : 32'h702cf003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e1, value : 32'h99642a2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e2, value : 32'hc380f9ef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e3, value : 32'h3100140c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e4, value : 32'h710478ca},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e5, value : 32'h7cb0b822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e6, value : 32'hc177b10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e7, value : 32'h24892030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e8, value : 32'he1b1fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551e9, value : 32'hb272051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ea, value : 32'hd9592071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551eb, value : 32'he17f016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ec, value : 32'hb232051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ed, value : 32'hd93e2071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ee, value : 32'hb17f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ef, value : 32'hd9552071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f0, value : 32'hb17f00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f1, value : 32'hd93a2071},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f2, value : 32'hd957f008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f3, value : 32'hd953f006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f4, value : 32'hd93cf004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f5, value : 32'hd938f002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f6, value : 32'h6909b99f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f7, value : 32'hc2608840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f8, value : 32'ha0dc220},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551f9, value : 32'h23890325},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551fa, value : 32'hc4200fc3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551fb, value : 32'h8900a880},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551fc, value : 32'hc020c060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551fd, value : 32'hc50807},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551fe, value : 32'ha960c320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h551ff, value : 32'h78e0c7d4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55200, value : 32'h1600c2ea},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55201, value : 32'h8000708e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55202, value : 32'h7114122a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55203, value : 32'hdd75d870},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55204, value : 32'h25ca4130},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55205, value : 32'h16001001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55206, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55207, value : 32'h877122b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55208, value : 32'h16000384},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55209, value : 32'h80007080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5520a, value : 32'h86712e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5520b, value : 32'h79cf03ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5520c, value : 32'hfdef0af2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5520d, value : 32'h46004022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5520e, value : 32'h742d70ec},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5520f, value : 32'h702c720d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55210, value : 32'h3822114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55211, value : 32'hba0cc809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55212, value : 32'h27157845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55213, value : 32'h702c0042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55214, value : 32'h2450937},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55215, value : 32'hae0e2d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55216, value : 32'h7b0561bb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55217, value : 32'h2305bb02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55218, value : 32'h90380f8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55219, value : 32'h265a0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5521a, value : 32'h7b541503},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5521b, value : 32'hf8b2334},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5521c, value : 32'h4db48001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5521d, value : 32'h800043c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5521e, value : 32'h23f40f68},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5521f, value : 32'hb46002c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55220, value : 32'h71447124},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55221, value : 32'h712cf1e6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55222, value : 32'h173f208d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55223, value : 32'h71c5752d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55224, value : 32'hc6caf1c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55225, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55226, value : 32'h44d3b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55227, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55228, value : 32'h14014018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55229, value : 32'h14002080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5522a, value : 32'h200c2090},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5522b, value : 32'h11aa000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5522c, value : 32'h4748002d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5522d, value : 32'hc172140},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5522e, value : 32'he45d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5522f, value : 32'h21400000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55230, value : 32'h21400816},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55231, value : 32'h21540402},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55232, value : 32'h21050819},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55233, value : 32'h2705055b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55234, value : 32'h26052557},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55235, value : 32'h25052556},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55236, value : 32'h46cb2095},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55237, value : 32'h9000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55238, value : 32'h800041c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55239, value : 32'h892012e1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5523a, value : 32'h40e09d5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5523b, value : 32'h2513205a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5523c, value : 32'h800145cb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5523d, value : 32'h7f604db4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5523e, value : 32'h23402334},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5523f, value : 32'h23512840},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55240, value : 32'h21055021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55241, value : 32'h75622612},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55242, value : 32'h26c22205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55243, value : 32'hb9027945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55244, value : 32'hb10079c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55245, value : 32'h95017f60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55246, value : 32'h25422205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55247, value : 32'h79455021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55248, value : 32'h79c5b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55249, value : 32'h7f60b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5524a, value : 32'h22059502},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5524b, value : 32'h50212582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5524c, value : 32'hb9027945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5524d, value : 32'hb10079c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5524e, value : 32'h95037f60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5524f, value : 32'h25d22205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55250, value : 32'h21055021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55251, value : 32'hb9020481},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55252, value : 32'hb10079c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55253, value : 32'h95047f60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55254, value : 32'h26112100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55255, value : 32'h21964100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55256, value : 32'hc8092008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55257, value : 32'h26c22105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55258, value : 32'hb8027845},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55259, value : 32'hb02078c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5525a, value : 32'h95057f60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5525b, value : 32'h25422105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5525c, value : 32'h79455021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5525d, value : 32'h79c5b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5525e, value : 32'h7f60b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5525f, value : 32'h21059506},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55260, value : 32'h50212582},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55261, value : 32'hb9027945},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55262, value : 32'hb10079c5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55263, value : 32'h95077f60},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55264, value : 32'h25c22105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55265, value : 32'h79455021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55266, value : 32'h79c5b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55267, value : 32'h7f60b100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55268, value : 32'h21059508},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55269, value : 32'h50212651},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5526a, value : 32'h4412105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5526b, value : 32'h2105b902},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5526c, value : 32'h90380f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5526d, value : 32'hb1000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5526e, value : 32'h20801401},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5526f, value : 32'ha000200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55270, value : 32'hffe50720},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55271, value : 32'h14047106},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55272, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55273, value : 32'h1cfcc2fa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55274, value : 32'h2482b6c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55275, value : 32'h45683802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55276, value : 32'hc0414630},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55277, value : 32'h700c702e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55278, value : 32'h31001c90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55279, value : 32'h30801c8c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5527a, value : 32'heb05c040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5527b, value : 32'hf84f0ab6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5527c, value : 32'h40dbc040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5527d, value : 32'hc0c49007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5527e, value : 32'hff2f0cd6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5527f, value : 32'h30451800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55280, value : 32'h30021c0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55281, value : 32'h702c710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55282, value : 32'hf1242a1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55283, value : 32'hc382f9af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55284, value : 32'h47d3722f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55285, value : 32'h122a8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55286, value : 32'hb89fd825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55287, value : 32'h881b8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55288, value : 32'h710c7905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55289, value : 32'h4402800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5528a, value : 32'h200fb802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5528b, value : 32'h782b0440},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5528c, value : 32'h1023c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5528d, value : 32'h208e1700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5528e, value : 32'h20801701},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5528f, value : 32'h2307610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55290, value : 32'h40c3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55291, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55292, value : 32'h20118800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55293, value : 32'h21a8380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55294, value : 32'h79cf0021},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55295, value : 32'hfdef08ce},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55296, value : 32'h3000148c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55297, value : 32'h131b2e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55298, value : 32'h1c94700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55299, value : 32'h14943000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5529a, value : 32'h20113000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5529b, value : 32'hf2f18400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5529c, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5529d, value : 32'h7a1b28f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5529e, value : 32'h211fc101},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5529f, value : 32'hb822200c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a0, value : 32'h230a794a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a1, value : 32'h261a1400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a2, value : 32'h42c31003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a3, value : 32'h1b448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a4, value : 32'h1184239a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a5, value : 32'h3088140d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a6, value : 32'h61796199},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a7, value : 32'h62387161},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a8, value : 32'h88a26157},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552a9, value : 32'h10300817},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552aa, value : 32'h14149022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ab, value : 32'h78aa3100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ac, value : 32'h71044528},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ad, value : 32'h671fb822},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ae, value : 32'h65fdf003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552af, value : 32'h28404728},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b0, value : 32'hc8092201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b1, value : 32'h6c12105},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b2, value : 32'hc0017905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b3, value : 32'h412214f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b4, value : 32'he80a4330},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b5, value : 32'h875639b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b6, value : 32'h23001030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b7, value : 32'h605802c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b8, value : 32'hf0399002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552b9, value : 32'h20110e23},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ba, value : 32'h1a00265a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552bb, value : 32'h4002015},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552bc, value : 32'h4402014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552bd, value : 32'hf812000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552be, value : 32'hbecc8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552bf, value : 32'h800070c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c0, value : 32'hb1e0c00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c1, value : 32'h2455b0a0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c2, value : 32'hd6239c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c3, value : 32'h78b0f96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c4, value : 32'he807ca05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c5, value : 32'h39c02455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c6, value : 32'hfb2f0c76},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c7, value : 32'h98e41c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c8, value : 32'he80afc8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552c9, value : 32'h16802600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ca, value : 32'h81101c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552cb, value : 32'hfb2f0c62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552cc, value : 32'h39c02455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552cd, value : 32'h24402205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ce, value : 32'h2005b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552cf, value : 32'h90000f8d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d0, value : 32'h24550048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d1, value : 32'hf07839c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d2, value : 32'h60506219},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d3, value : 32'h60388922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d4, value : 32'hd1a7810},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d5, value : 32'h2455f96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d6, value : 32'h240039c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d7, value : 32'h3f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d8, value : 32'hd0a009a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552d9, value : 32'h78b0f96f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552da, value : 32'he806c000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552db, value : 32'h3100149a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552dc, value : 32'h30041c9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552dd, value : 32'he80eca05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552de, value : 32'h39c02455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552df, value : 32'hfb2f0c12},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e0, value : 32'h240041c2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e1, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e2, value : 32'hc06009a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e3, value : 32'h41c2fb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e4, value : 32'hfc8f091a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e5, value : 32'h2600e811},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e6, value : 32'h24551694},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e7, value : 32'hbf239c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e8, value : 32'h141cfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552e9, value : 32'h24002081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ea, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552eb, value : 32'hbe2009a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ec, value : 32'h141cfb2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ed, value : 32'hca052081},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ee, value : 32'h8f2e887},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ef, value : 32'h89ffc8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f0, value : 32'h24550030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f1, value : 32'h245539c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f2, value : 32'h240039c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f3, value : 32'h3f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f4, value : 32'h724c009a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f5, value : 32'hfd0f08ae},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f6, value : 32'h20310e35},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f7, value : 32'h39c02455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f8, value : 32'h1a15265a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552f9, value : 32'h800044d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552fa, value : 32'h2515c00c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552fb, value : 32'h25142415},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552fc, value : 32'hbd62455},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552fd, value : 32'h2400f82f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552fe, value : 32'h1c002554},
                          '{ step_type : REG_WRITE, reg_addr : 32'h552ff, value : 32'h25002004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55300, value : 32'h80002f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55301, value : 32'h1ca0becc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55302, value : 32'hb0e02344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55303, value : 32'h244d2205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55304, value : 32'h2505bd02},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55305, value : 32'h90001f92},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55306, value : 32'hba20048},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55307, value : 32'h2455f82f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55308, value : 32'hbd8639c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55309, value : 32'h20041a00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5530a, value : 32'h2400bd9c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5530b, value : 32'h3f80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5530c, value : 32'hbd9f009a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5530d, value : 32'hf80f0b86},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5530e, value : 32'h1490b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5530f, value : 32'he8093000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55310, value : 32'h20802b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55311, value : 32'hf802005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55312, value : 32'h3209004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55313, value : 32'h7106b0e0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55314, value : 32'ha240204c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55315, value : 32'hffc50612},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55316, value : 32'h2400f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55317, value : 32'h3f81},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55318, value : 32'h714c009a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55319, value : 32'h5d5f1b8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5531a, value : 32'h71c5ffef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5531b, value : 32'h35bb218d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5531c, value : 32'h1800712e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5531d, value : 32'h24803005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5531e, value : 32'h14043802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5531f, value : 32'hc6da341b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55320, value : 32'h1600c3f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55321, value : 32'h80007091},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55322, value : 32'ha460004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55323, value : 32'h2482ff2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55324, value : 32'h1c053102},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55325, value : 32'h710c3002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55326, value : 32'h704c712c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55327, value : 32'hf9af0c7e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55328, value : 32'h2153c380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55329, value : 32'h718e20d1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5532a, value : 32'h726e700e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5532b, value : 32'h47cb714e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5532c, value : 32'h12288000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5532d, value : 32'hb89fd825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5532e, value : 32'h881b8820},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5532f, value : 32'h2c007905},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55330, value : 32'hb8022400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55331, value : 32'h400200f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55332, value : 32'hf2c1782b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55333, value : 32'h8f038fc2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55334, value : 32'h17a7610},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55335, value : 32'h40c3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55336, value : 32'h12e18000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55337, value : 32'h20118800},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55338, value : 32'hf2b38380},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55339, value : 32'h13002e40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5533a, value : 32'h30881405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5533b, value : 32'h4012005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5533c, value : 32'h7825c809},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5533d, value : 32'h7280244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5533e, value : 32'h706d6892},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5533f, value : 32'h1f892405},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55340, value : 32'ha09004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55341, value : 32'ha0020a8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55342, value : 32'h40c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55343, value : 32'h68320a3c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55344, value : 32'h201f78cc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55345, value : 32'h41c32042},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55346, value : 32'h1b448000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55347, value : 32'h4061621a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55348, value : 32'h184209a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55349, value : 32'h1030080d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5534a, value : 32'h60386058},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5534b, value : 32'hf0069002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5534c, value : 32'h6030611b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5534d, value : 32'h60788b62},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5534e, value : 32'h12710b0f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5534f, value : 32'h12832b40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55350, value : 32'h10041900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55351, value : 32'h7b85f007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55352, value : 32'hf832305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55353, value : 32'h1e89004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55354, value : 32'h7165b300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55355, value : 32'h70801600},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55356, value : 32'hee8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55357, value : 32'hf4757014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55358, value : 32'h10100821},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55359, value : 32'h6159622d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5535a, value : 32'h140c8922},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5535b, value : 32'h782a3100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5535c, value : 32'h20047104},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5535d, value : 32'hf80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5535e, value : 32'hb822fffc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5535f, value : 32'hf004651d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55360, value : 32'h89a46159},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55361, value : 32'h8118f05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55362, value : 32'h720c03a5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55363, value : 32'hf88f0afa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55364, value : 32'hf006710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55365, value : 32'hf8af0af2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55366, value : 32'h700c710c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55367, value : 32'h4002af00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55368, value : 32'hfa2f0b82},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55369, value : 32'h451041c1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5536a, value : 32'hb7a4002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5536b, value : 32'h41c1fa2f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5536c, value : 32'h2b01215f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5536d, value : 32'h2078},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5536e, value : 32'h7404b802},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5536f, value : 32'h8f006119},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55370, value : 32'h2114},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55371, value : 32'h700279af},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55372, value : 32'ha8a860f8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55373, value : 32'h20002578},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55374, value : 32'hb526841},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55375, value : 32'h4002f62f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55376, value : 32'h20300d17},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55377, value : 32'he8118f00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55378, value : 32'h20100a3b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55379, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5537a, value : 32'h508000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5537b, value : 32'he810f02a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5537c, value : 32'h20100a35},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5537d, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5537e, value : 32'hfa8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5537f, value : 32'ha33f022},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55380, value : 32'h1e002010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55381, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55382, value : 32'hf01c0035},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55383, value : 32'h20100a2d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55384, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55385, value : 32'hf08000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55386, value : 32'h1e00f014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55387, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55388, value : 32'hf0100051},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55389, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5538a, value : 32'hff8000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5538b, value : 32'h1e00f00a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5538c, value : 32'h80007342},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5538d, value : 32'hf0060036},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5538e, value : 32'h73421e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5538f, value : 32'hf58000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55390, value : 32'hf8af0a46},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55391, value : 32'h71c5730c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55392, value : 32'h704ef143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55393, value : 32'h2d3c238d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55394, value : 32'hc7d2710e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55395, value : 32'h7a00244a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55396, value : 32'h800040c3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55397, value : 32'h20a8c44c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55398, value : 32'h180001c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h55399, value : 32'h20800003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5539a, value : 32'h7ee0000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5539b, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5539c, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5539d, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5539e, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5539f, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h553a0, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h553a1, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h553a2, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h553a3, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0080, value : 32'h7}, // [dwc_ddrphy_phyinit_D_loadIMEM] WriteImem: COMPLETED
//phyinit_io_write: 0xc0080, 0x7
// [dwc_ddrphy_phyinit_D_loadIMEM] End of dwc_ddrphy_phyinit_D_loadIMEM
// [dwc_ddrphy_phyinit_getPsExecOrder] pRuntimeConfig->psExecOrder[3] = 0x0
//Start of dwc_ddrphy_phyinit_C_initPhyConfigPsLoop(), PState=1, tck_ps=1666ps
                          '{ step_type : REG_WRITE, reg_addr : 32'h2008b, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, programming PState = 1
                          '{ step_type : REG_WRITE, reg_addr : 32'h190801, value : 32'hc0a2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming Seq0BGPR1 to 0xc0a2
                          '{ step_type : REG_WRITE, reg_addr : 32'h190802, value : 32'h0}, //phyinit_io_write: 0x190801, 0xc0a2
                          '{ step_type : REG_WRITE, reg_addr : 32'h190806, value : 32'h1}, //phyinit_io_write: 0x190802, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1a03ff, value : 32'h4101}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming OdtSeg120 to 0x4101
                          '{ step_type : REG_WRITE, reg_addr : 32'h1a030b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming ZCalCompCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h160008, value : 32'ha9a}, //[dwc_ddrphy_phyinit_programPLL] [phyinit_C_initPhyConfigPsLoop] Pstate=1,  Memclk=600MHz, Programming CpllCtrl5 to 0xa9a.
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e0, value : 32'h4b}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY0 to 0x4b (0.5us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e1, value : 32'he1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY1 to 0xe1 (tZQCal PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e2, value : 32'h5dc}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY2 to 0x5dc (10.us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e3, value : 32'h58}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY3 to 0x58 (dllLock PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e4, value : 32'hf}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY4 to 0xf (0.1us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e5, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY5 to 0x0 (RxReplicaCalWait delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e6, value : 32'h43}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY6 to 0x43 (Oscillator PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e7, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY7 to 0x0 (tXDSM_XP PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908ea, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY10 to 0x3 (tPDXCSODTON 20ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908eb, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY11 to 0x3 (20ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908ec, value : 32'h8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY12 to 0x8 (50ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908ed, value : 32'h3b}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming Seq0BDLY13 to 0x3b (tXSR PIE delay, tRFCab delay is 380ns)
                          '{ step_type : REG_WRITE, reg_addr : 32'h120002, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming PclkPtrInitVal to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h160040, value : 32'h3}, //phyinit_io_write: 0x120002, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h120000, value : 32'h2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DfiFreqRatio to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h1100fb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming RxDigStrbEn to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1110fb, value : 32'h0}, //phyinit_io_write: 0x1100fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1120fb, value : 32'h0}, //phyinit_io_write: 0x1110fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1130fb, value : 32'h0}, //phyinit_io_write: 0x1120fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e000b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DxDigStrobeMode HMDBYTE to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e100b, value : 32'h0}, //phyinit_io_write: 0x1e000b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e200b, value : 32'h0}, //phyinit_io_write: 0x1e100b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e300b, value : 32'h0}, //phyinit_io_write: 0x1e200b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e400b, value : 32'h0}, //phyinit_io_write: 0x1e300b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e500b, value : 32'h0}, //phyinit_io_write: 0x1e400b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e600b, value : 32'h0}, //phyinit_io_write: 0x1e500b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e700b, value : 32'h0}, //phyinit_io_write: 0x1e600b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h110024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE0.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h111024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE1.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h112024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE2.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h113024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE3.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h110025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE0.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h111025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE1.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h112025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE2.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h113025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE3.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h110004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE0.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h110003, value : 32'h0}, //phyinit_io_write: 0x110004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h111004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE1.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h111003, value : 32'h0}, //phyinit_io_write: 0x111004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h112004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE2.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h112003, value : 32'h0}, //phyinit_io_write: 0x112004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h113004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE3.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h113003, value : 32'h0}, //phyinit_io_write: 0x113004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1b0004, value : 32'h258}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ZCalClkInfo::ZCalDfiClkTicksPer1uS to 0x258
                          '{ step_type : REG_WRITE, reg_addr : 32'h1a030c, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h11003e, value : 32'h5}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE RxGainCurrAdjRxReplica to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h11103e, value : 32'h5}, //phyinit_io_write: 0x11003e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h11203e, value : 32'h5}, //phyinit_io_write: 0x11103e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h11303e, value : 32'h5}, //phyinit_io_write: 0x11203e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h120003, value : 32'h1}, //phyinit_io_write: 0x11303e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h12000b, value : 32'h1111}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming CPclkDivRatio to 0x1111
                          '{ step_type : REG_WRITE, reg_addr : 32'h110108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE0.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h111108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE1.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h112108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE2.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h113108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming DBYTE3.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70005, value : 32'h0}, //[phyinit_C_initPhyConfig] Programming EnPhyUpdZQCalUpdate to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h7000f, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming DisableZQupdateOnSnoop to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11000e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h11100e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h11200e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h11300e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h120019, value : 32'h4}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming EnRxDqsTracking::DqsSampNegRxEnSense to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e002c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 0 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e102c, value : 32'h33}, //phyinit_io_write: 0x1e002c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e002d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 0 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e102d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 0 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e202c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 1 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e302c, value : 32'h33}, //phyinit_io_write: 0x1e202c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e202d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 1 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e302d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 1 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e402c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 2 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e502c, value : 32'h33}, //phyinit_io_write: 0x1e402c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e402d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 2 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e502d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 2 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e602c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 3 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e702c, value : 32'h33}, //phyinit_io_write: 0x1e602c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e602d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 3 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e702d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 3 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h100070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC0 Instance0 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h101070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC1 Instance1 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h102070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC2 Instance2 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h103070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC3 Instance3 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h104070, value : 32'hff}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming AC0 HMAC4 Instance4 CS TxImpedanceAC::TxStrenCodePDAC to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h105070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC5 Instance5 TxImpedanceAC::TxStrenCodePD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h107070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC0 Instance7 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h108070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC1 Instance8 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h109070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC2 Instance9 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC3 Instance10 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b070, value : 32'hff}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming AC1 HMAC4 Instance11 CS TxImpedanceAC::TxStrenCodePDAC to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC5 Instance12 TxImpedanceAC::TxStrenCodePD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e002e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 0 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e102e, value : 32'h30}, //phyinit_io_write: 0x1e002e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e002f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 0 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e102f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 0 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e202e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 1 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e302e, value : 32'h30}, //phyinit_io_write: 0x1e202e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e202f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 1 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e302f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 1 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e402e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 2 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e502e, value : 32'h30}, //phyinit_io_write: 0x1e402e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e402f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 2 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e502f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 2 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e602e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 3 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e702e, value : 32'h30}, //phyinit_io_write: 0x1e602e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e602f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 3 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e702f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 3 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h100079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC0 Instance0 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h101079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC1 Instance1 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h102079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC2 Instance2 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h103079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC3 Instance3 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h104079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC4 Instance4 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h105079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC5 DIFF5 OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h107079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC0 Instance7 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h108079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC1 Instance8 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h109079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC2 Instance9 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC3 Instance10 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC4 Instance11 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC5 DIFF12 OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e001c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 0 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e101c, value : 32'h3}, //phyinit_io_write: 0x1e001c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e201c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 1 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e301c, value : 32'h3}, //phyinit_io_write: 0x1e201c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e401c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 2 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e501c, value : 32'h3}, //phyinit_io_write: 0x1e401c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e601c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming HMDBYTE 3 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e701c, value : 32'h3}, //phyinit_io_write: 0x1e601c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h10006d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC0 Instance0 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10106d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC1 Instance1 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10206d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC2 Instance2 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10306d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC3 Instance3 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10406d, value : 32'hf8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC4 Instance4 CS TxSlewAC::TxSlewPDAC to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h10506d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX0 HMAC5 Instance5 TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10706d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC0 Instance7 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10806d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC1 Instance8 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10906d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC2 Instance9 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a06d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC3 Instance10 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b06d, value : 32'hf8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC4 Instance11 CS TxSlewAC::TxSlewPDAC to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c06d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACX1 HMAC5 Instance12 TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e003e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Programming HMDBYTE RxDQSCtrl::RxDQSDiffSeVrefDACEn to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e103e, value : 32'h0}, //phyinit_io_write: 0x1e003e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e203e, value : 32'h0}, //phyinit_io_write: 0x1e103e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e303e, value : 32'h0}, //phyinit_io_write: 0x1e203e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e403e, value : 32'h0}, //phyinit_io_write: 0x1e303e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e503e, value : 32'h0}, //phyinit_io_write: 0x1e403e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e603e, value : 32'h0}, //phyinit_io_write: 0x1e503e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e703e, value : 32'h0}, //phyinit_io_write: 0x1e603e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h110001, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming WriteLinkEcc to 0
                          '{ step_type : REG_WRITE, reg_addr : 32'h111001, value : 32'h0}, //phyinit_io_write: 0x110001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h112001, value : 32'h0}, //phyinit_io_write: 0x111001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h113001, value : 32'h0}, //phyinit_io_write: 0x112001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h170040, value : 32'h5a}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming PPTTrainSetup::PhyMstrMaxReqToAck to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h170041, value : 32'hf}, //phyinit_io_write: 0x170040, 0x5a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1100a5, value : 32'h1}, //phyinit_io_write: 0x170041, 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h1110a5, value : 32'h1}, //phyinit_io_write: 0x1100a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1120a5, value : 32'h1}, //phyinit_io_write: 0x1110a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1130a5, value : 32'h1}, //phyinit_io_write: 0x1120a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h110209, value : 32'h3232}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Programming RxReplicaRangeVal 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h111209, value : 32'h3232}, //phyinit_io_write: 0x110209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h112209, value : 32'h3232}, //phyinit_io_write: 0x111209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h113209, value : 32'h3232}, //phyinit_io_write: 0x112209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h11020f, value : 32'h6}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Programming RxReplicaCtl04 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h11120f, value : 32'h6}, //phyinit_io_write: 0x11020f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h11220f, value : 32'h6}, //phyinit_io_write: 0x11120f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h11320f, value : 32'h6}, //phyinit_io_write: 0x11220f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h120005, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, DfiFreq=600MHz, Programming PipeCtl[AcInPipeEn]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h110008, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, DfiFreq=600MHz, Programming DBYTE0.LP5DfiDataEnLatency[LP5RLm13]=0x1 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h111008, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, DfiFreq=600MHz, Programming DBYTE1.LP5DfiDataEnLatency[LP5RLm13]=0x1 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h112008, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, DfiFreq=600MHz, Programming DBYTE2.LP5DfiDataEnLatency[LP5RLm13]=0x1 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h113008, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, DfiFreq=600MHz, Programming DBYTE3.LP5DfiDataEnLatency[LP5RLm13]=0x1 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h17006b, value : 32'h222}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, DfiFreq=600MHz, Programming DfiHandshakeDelays[PhyUpdReqDelay]=0x2 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h170066, value : 32'h20}, //phyinit_io_write: 0x17006b, 0x222
                          '{ step_type : REG_WRITE, reg_addr : 32'h1700eb, value : 32'h222}, //phyinit_io_write: 0x170066, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h1700e6, value : 32'h20}, //phyinit_io_write: 0x1700eb, 0x222
                          '{ step_type : REG_WRITE, reg_addr : 32'h170135, value : 32'hc08}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACSMWckWriteFastTogglePulse::ACSMWckWriteFastToggleWidth to 0x19, ACSMWckWriteFastTogglePulse::ACSMWckWriteFastToggleDelay to 0x18
                          '{ step_type : REG_WRITE, reg_addr : 32'h170136, value : 32'hc08}, //phyinit_io_write: 0x170135, 0xc08
                          '{ step_type : REG_WRITE, reg_addr : 32'h170137, value : 32'h414}, //phyinit_io_write: 0x170136, 0xc08
                          '{ step_type : REG_WRITE, reg_addr : 32'h170138, value : 32'h1918}, //phyinit_io_write: 0x170137, 0x414
                          '{ step_type : REG_WRITE, reg_addr : 32'h170139, value : 32'hc10}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACSMWckReadFastTogglePulse::ACSMWckReadFastToggleWidth to 0x29, ACSMWckReadFastTogglePulse::ACSMWckReadFastToggleDelay to 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h17013a, value : 32'hc10}, //phyinit_io_write: 0x170139, 0xc10
                          '{ step_type : REG_WRITE, reg_addr : 32'h17013b, value : 32'h41c}, //phyinit_io_write: 0x17013a, 0xc10
                          '{ step_type : REG_WRITE, reg_addr : 32'h17013c, value : 32'h2920}, //phyinit_io_write: 0x17013b, 0x41c
                          '{ step_type : REG_WRITE, reg_addr : 32'h17013d, value : 32'hc04}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACSMWckFreqFastTogglePulse::ACSMWckFreqFastToggleWidth to 0x11, ACSMWckFreqFastTogglePulse::ACSMWckFreqFastToggleDelay to 0x14
                          '{ step_type : REG_WRITE, reg_addr : 32'h17013e, value : 32'hc04}, //phyinit_io_write: 0x17013d, 0xc04
                          '{ step_type : REG_WRITE, reg_addr : 32'h17013f, value : 32'h410}, //phyinit_io_write: 0x17013e, 0xc04
                          '{ step_type : REG_WRITE, reg_addr : 32'h170140, value : 32'h1114}, //phyinit_io_write: 0x17013f, 0x410
                          '{ step_type : REG_WRITE, reg_addr : 32'h17012c, value : 32'h827}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACSMRxValPulse::ACSMRxValDelay to 0x27, ACSMRxValPulse::ACSMRxValWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h17012d, value : 32'h827}, //phyinit_io_write: 0x17012c, 0x827
                          '{ step_type : REG_WRITE, reg_addr : 32'h170130, value : 32'h827}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACSMRdcsPulse::ACSMRdcsDelay to 0x27, ACSMRdcsPulse::ACSMRdcsWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h17012e, value : 32'h817}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACSMTxEnPulse::ACSMTxEnDelay to 0x17, ACSMTxEnPulse::ACSMTxEnWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h17012f, value : 32'h817}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming ACSMWrcsPulse::ACSMWrcsDelay to 0x17, ACSMWrcsPulse::ACSMWrcsWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h130008, value : 32'h0}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming AcPipeEn AC0 to 0. DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h131008, value : 32'h0}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, Programming AcPipeEn AC1 to 0. DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1013, value : 32'h0}, //phyinit_io_write: 0x1e0013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3013, value : 32'h0}, //phyinit_io_write: 0x1e2013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5013, value : 32'h0}, //phyinit_io_write: 0x1e4013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7013, value : 32'h0}, //phyinit_io_write: 0x1e6013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1005e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC0 Instance0 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1015e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC1 Instance1 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1025e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC2 Instance2 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1035e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC3 Instance3 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1045e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC4 Instance4 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1055e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC5 Instance5 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1075e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC0 Instance7 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1085e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC1 Instance8 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1095e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC2 Instance9 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a5e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC3 Instance10 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b5e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC4 Instance11 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c5e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC5 Instance12 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e05e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming HMDBYTE0 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e15e3, value : 32'h4}, //phyinit_io_write: 0x1e05e3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e25e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming HMDBYTE1 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e35e3, value : 32'h4}, //phyinit_io_write: 0x1e25e3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e45e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming HMDBYTE2 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e55e3, value : 32'h4}, //phyinit_io_write: 0x1e45e3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e65e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming HMDBYTE3 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e75e3, value : 32'h4}, //phyinit_io_write: 0x1e65e3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h10050a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC0 Instance0 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10150a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC1 Instance1 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10250a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC2 Instance2 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10350a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC3 Instance3 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10450a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC4 Instance4 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10550a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC5 Instance5 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10750a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC0 Instance7 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10850a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC1 Instance8 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10950a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC2 Instance9 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a50a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC3 Instance10 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b50a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC4 Instance11 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c50a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC5 Instance12 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11080b, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming DBYTE0 PclkDCASampDelayLCDLDB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11180b, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming DBYTE1 PclkDCASampDelayLCDLDB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11280b, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming DBYTE2 PclkDCASampDelayLCDLDB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11380b, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming DBYTE3 PclkDCASampDelayLCDLDB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h130803, value : 32'h105a}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming PclkDCAStaticCtr0AC to 0x105a
                          '{ step_type : REG_WRITE, reg_addr : 32'h131803, value : 32'h105a}, //phyinit_io_write: 0x130803, 0x105a
                          '{ step_type : REG_WRITE, reg_addr : 32'h110803, value : 32'h105a}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming PclkDCAStaticCtr0DB to 0x105a
                          '{ step_type : REG_WRITE, reg_addr : 32'h111803, value : 32'h105a}, //phyinit_io_write: 0x110803, 0x105a
                          '{ step_type : REG_WRITE, reg_addr : 32'h112803, value : 32'h105a}, //phyinit_io_write: 0x111803, 0x105a
                          '{ step_type : REG_WRITE, reg_addr : 32'h113803, value : 32'h105a}, //phyinit_io_write: 0x112803, 0x105a
                          '{ step_type : REG_WRITE, reg_addr : 32'h100503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC0 Instance0 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h101503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC1 Instance1 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h102503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC2 Instance2 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h103503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC3 Instance3 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h104503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC4 Instance4 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h105503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC5 Instance5 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h107503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC0 Instance7 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h108503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC1 Instance8 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h109503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC2 Instance9 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC3 Instance10 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC4 Instance11 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c503, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC5 Instance12 PclkDCAStaticCtrl1AC to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h110c03, value : 32'h1b}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming PclkDCAStaticCtrl1DB to 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h111c03, value : 32'h1b}, //phyinit_io_write: 0x110c03, 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h112c03, value : 32'h1b}, //phyinit_io_write: 0x111c03, 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h113c03, value : 32'h1b}, //phyinit_io_write: 0x112c03, 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h100110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC0 Instance0 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h101110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC1 Instance1 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h102110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC2 Instance2 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h103110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC3 Instance3 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h104110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC4 Instance4 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h105110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX0 HMAC5 Instance5 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h107110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC0 Instance7 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h108110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC1 Instance8 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h109110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC2 Instance9 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC3 Instance10 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC4 Instance11 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming ACX1 HMAC5 Instance12 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming HMDBYTE0 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1110, value : 32'h1f}, //phyinit_io_write: 0x1e0110, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming HMDBYTE1 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3110, value : 32'h1f}, //phyinit_io_write: 0x1e2110, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming HMDBYTE2 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5110, value : 32'h1f}, //phyinit_io_write: 0x1e4110, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming HMDBYTE3 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7110, value : 32'h1f}, //phyinit_io_write: 0x1e6110, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e8, value : 32'h11}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=1, Programming Seq0BDLY9 to 57
                          '{ step_type : REG_WRITE, reg_addr : 32'h1908e9, value : 32'h39}, //phyinit_io_write: 0x1908e8, 0x11
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0002, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Programming HMDBYTE RxDFECtrlDq to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1002, value : 32'h0}, //phyinit_io_write: 0x1e0002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2002, value : 32'h0}, //phyinit_io_write: 0x1e1002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3002, value : 32'h0}, //phyinit_io_write: 0x1e2002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4002, value : 32'h0}, //phyinit_io_write: 0x1e3002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5002, value : 32'h0}, //phyinit_io_write: 0x1e4002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6002, value : 32'h0}, //phyinit_io_write: 0x1e5002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7002, value : 32'h0}, //phyinit_io_write: 0x1e6002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11010b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=1, Memclk=600MHz, freqThreshold=200MHz, NoRDQS=0 Programming InhibitTxRdPtrInit::DisableRxEnDlyLoad to 0x0, InhibitTxRdPtrInit::DisableTxDqDly to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11110b, value : 32'h0}, //phyinit_io_write: 0x11010b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11210b, value : 32'h0}, //phyinit_io_write: 0x11110b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11310b, value : 32'h0}, //phyinit_io_write: 0x11210b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h100063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC0 Instance0 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h101063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC1 Instance1 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h102063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC2 Instance2 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h103063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC3 Instance3 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h104063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC4 Instance4 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h105063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC5 Instance5 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h107063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC0 Instance7 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h108063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC1 Instance8 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h109063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC2 Instance9 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC3 Instance10 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC4 Instance11 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c063, value : 32'h8a}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC5 Instance12 HMTxLcdlSeed HMTxSeed to 0x8a HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h19080a, value : 32'h28a}, //[dwc_ddrphy_phyinit_programLCDLSeed] Programming Seq0BGPR10 to HMTxLcdlSeed Full search value = 0x28a
                          '{ step_type : REG_WRITE, reg_addr : 32'h19080b, value : 32'h8a}, //phyinit_io_write: 0x19080a, 0x28a
                          '{ step_type : REG_WRITE, reg_addr : 32'h190815, value : 32'h28a}, //[dwc_ddrphy_phyinit_programLCDLSeed] Programming Seq0BGPR21 to ACHMTxLcdlSeed Full search value = 0x28a
                          '{ step_type : REG_WRITE, reg_addr : 32'h190816, value : 32'h8a}, //phyinit_io_write: 0x190815, 0x28a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0063, value : 32'h8a}, //phyinit_io_write: 0x190816, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0064, value : 32'h8a}, //phyinit_io_write: 0x1e0063, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0087, value : 32'h8a}, //phyinit_io_write: 0x1e0064, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1063, value : 32'h8a}, //phyinit_io_write: 0x1e0087, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1064, value : 32'h8a}, //phyinit_io_write: 0x1e1063, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1087, value : 32'h8a}, //phyinit_io_write: 0x1e1064, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2063, value : 32'h8a}, //phyinit_io_write: 0x1e1087, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2064, value : 32'h8a}, //phyinit_io_write: 0x1e2063, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2087, value : 32'h8a}, //phyinit_io_write: 0x1e2064, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3063, value : 32'h8a}, //phyinit_io_write: 0x1e2087, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3064, value : 32'h8a}, //phyinit_io_write: 0x1e3063, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3087, value : 32'h8a}, //phyinit_io_write: 0x1e3064, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4063, value : 32'h8a}, //phyinit_io_write: 0x1e3087, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4064, value : 32'h8a}, //phyinit_io_write: 0x1e4063, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4087, value : 32'h8a}, //phyinit_io_write: 0x1e4064, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5063, value : 32'h8a}, //phyinit_io_write: 0x1e4087, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5064, value : 32'h8a}, //phyinit_io_write: 0x1e5063, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5087, value : 32'h8a}, //phyinit_io_write: 0x1e5064, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6063, value : 32'h8a}, //phyinit_io_write: 0x1e5087, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6064, value : 32'h8a}, //phyinit_io_write: 0x1e6063, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6087, value : 32'h8a}, //phyinit_io_write: 0x1e6064, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7063, value : 32'h8a}, //phyinit_io_write: 0x1e6087, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7064, value : 32'h8a}, //phyinit_io_write: 0x1e7063, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7087, value : 32'h8a}, //phyinit_io_write: 0x1e7064, 0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0080, value : 32'h7}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming UcclkHclkEnables to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e003c, value : 32'h80}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming RxDQSSeVrefDAC0 to 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e103c, value : 32'h80}, //phyinit_io_write: 0x1e003c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e203c, value : 32'h80}, //phyinit_io_write: 0x1e103c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e303c, value : 32'h80}, //phyinit_io_write: 0x1e203c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e403c, value : 32'h80}, //phyinit_io_write: 0x1e303c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e503c, value : 32'h80}, //phyinit_io_write: 0x1e403c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e603c, value : 32'h80}, //phyinit_io_write: 0x1e503c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e703c, value : 32'h80}, //phyinit_io_write: 0x1e603c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h190817, value : 32'h3e}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 1 Seq0BGPR23 to 0x3e, NumMemClk_tRFCab=246.0, NumMemClk_7p5ns=4.5, NumMemClk_tXSR=250.5
                          '{ step_type : REG_WRITE, reg_addr : 32'h190818, value : 32'h0}, //phyinit_io_write: 0x190817, 0x3e
                          '{ step_type : REG_WRITE, reg_addr : 32'h190819, value : 32'h0}, //phyinit_io_write: 0x190818, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1300eb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 1 AC0 AcLcdlUpdInterval to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1310eb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 1 AC1 AcLcdlUpdInterval to 0x0
//[dwc_ddrphy_phyinit_programDfiMode] Skip DfiMode Programming: Keeping the reset value of 0x3
//End of dwc_ddrphy_phyinit_C_initPhyConfigPsLoop(), Pstate=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h60006, value : 32'h1f0}, //[dwc_ddrphy_phyinit_progCsrSkipTrain] Programming CPllCtrl3 to 0x1f0
                          '{ step_type : REG_WRITE, reg_addr : 32'h100d9, value : 32'h9c}, //[dwc_ddrphy_phyinit_progCsrSkipTrain] RxReplica Programming RxReplicaUICalWait to 0x9c
                          '{ step_type : REG_WRITE, reg_addr : 32'h110d9, value : 32'h9c}, //phyinit_io_write: 0x100d9, 0x9c
                          '{ step_type : REG_WRITE, reg_addr : 32'h120d9, value : 32'h9c}, //phyinit_io_write: 0x110d9, 0x9c
                          '{ step_type : REG_WRITE, reg_addr : 32'h130d9, value : 32'h9c}, //phyinit_io_write: 0x120d9, 0x9c
                          '{ step_type : REG_WRITE, reg_addr : 32'h10027, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrain] Programming RxClkCntl1 to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h11027, value : 32'h1}, //phyinit_io_write: 0x10027, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h12027, value : 32'h1}, //phyinit_io_write: 0x11027, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h13027, value : 32'h1}, //phyinit_io_write: 0x12027, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h30022, value : 32'h3}, // [dwc_ddrphy_phyinit_programMemResetL] Programming MemResetL AC 0to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h31022, value : 32'h3}, // [dwc_ddrphy_phyinit_programMemResetL] Programming MemResetL AC 1to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1300d9, value : 32'h40}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming CKXTxDly to 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1300d8, value : 32'h40}, //phyinit_io_write: 0x1300d9, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1301d8, value : 32'h40}, //phyinit_io_write: 0x1300d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1302d8, value : 32'h40}, //phyinit_io_write: 0x1301d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303d8, value : 32'h40}, //phyinit_io_write: 0x1302d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1304d8, value : 32'h40}, //phyinit_io_write: 0x1303d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1305d8, value : 32'h40}, //phyinit_io_write: 0x1304d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1306d8, value : 32'h40}, //phyinit_io_write: 0x1305d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1308d8, value : 32'h40}, //phyinit_io_write: 0x1306d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1309d8, value : 32'h40}, //phyinit_io_write: 0x1308d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1310d9, value : 32'h40}, //phyinit_io_write: 0x1309d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1310d8, value : 32'h40}, //phyinit_io_write: 0x1310d9, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1311d8, value : 32'h40}, //phyinit_io_write: 0x1310d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1312d8, value : 32'h40}, //phyinit_io_write: 0x1311d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1313d8, value : 32'h40}, //phyinit_io_write: 0x1312d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1314d8, value : 32'h40}, //phyinit_io_write: 0x1313d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1315d8, value : 32'h40}, //phyinit_io_write: 0x1314d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1316d8, value : 32'h40}, //phyinit_io_write: 0x1315d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1318d8, value : 32'h40}, //phyinit_io_write: 0x1316d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h1319d8, value : 32'h40}, //phyinit_io_write: 0x1318d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h110000, value : 32'h7}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming HwtMRL to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h111000, value : 32'h7}, //phyinit_io_write: 0x110000, 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h112000, value : 32'h7}, //phyinit_io_write: 0x111000, 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h113000, value : 32'h7}, //phyinit_io_write: 0x112000, 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h17000d, value : 32'h7}, //phyinit_io_write: 0x113000, 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h11002a, value : 32'h200}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming TxWckDlyTg0/Tg1 to 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h11002b, value : 32'h200}, //phyinit_io_write: 0x11002a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h11102a, value : 32'h200}, //phyinit_io_write: 0x11002b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h11102b, value : 32'h200}, //phyinit_io_write: 0x11102a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h11202a, value : 32'h200}, //phyinit_io_write: 0x11102b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h11202b, value : 32'h200}, //phyinit_io_write: 0x11202a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h11302a, value : 32'h200}, //phyinit_io_write: 0x11202b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h11302b, value : 32'h200}, //phyinit_io_write: 0x11302a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h110028, value : 32'hba}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming TxDqsDlyTg0/Tg1 to 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h110029, value : 32'hba}, //phyinit_io_write: 0x110028, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h111028, value : 32'hba}, //phyinit_io_write: 0x110029, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h111029, value : 32'hba}, //phyinit_io_write: 0x111028, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h112028, value : 32'hba}, //phyinit_io_write: 0x111029, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h112029, value : 32'hba}, //phyinit_io_write: 0x112028, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h113028, value : 32'hba}, //phyinit_io_write: 0x112029, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h113029, value : 32'hba}, //phyinit_io_write: 0x113028, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11007a, value : 32'hba}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming TxDqDlyTg0/Tg1 to 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11007b, value : 32'hba}, //phyinit_io_write: 0x11007a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11017a, value : 32'hba}, //phyinit_io_write: 0x11007b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11017b, value : 32'hba}, //phyinit_io_write: 0x11017a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11027a, value : 32'hba}, //phyinit_io_write: 0x11017b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11027b, value : 32'hba}, //phyinit_io_write: 0x11027a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11037a, value : 32'hba}, //phyinit_io_write: 0x11027b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11037b, value : 32'hba}, //phyinit_io_write: 0x11037a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11047a, value : 32'hba}, //phyinit_io_write: 0x11037b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11047b, value : 32'hba}, //phyinit_io_write: 0x11047a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11057a, value : 32'hba}, //phyinit_io_write: 0x11047b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11057b, value : 32'hba}, //phyinit_io_write: 0x11057a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11067a, value : 32'hba}, //phyinit_io_write: 0x11057b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11067b, value : 32'hba}, //phyinit_io_write: 0x11067a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11077a, value : 32'hba}, //phyinit_io_write: 0x11067b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11077b, value : 32'hba}, //phyinit_io_write: 0x11077a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11087a, value : 32'hba}, //phyinit_io_write: 0x11077b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11087b, value : 32'hba}, //phyinit_io_write: 0x11087a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11107a, value : 32'hba}, //phyinit_io_write: 0x11087b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11107b, value : 32'hba}, //phyinit_io_write: 0x11107a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11117a, value : 32'hba}, //phyinit_io_write: 0x11107b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11117b, value : 32'hba}, //phyinit_io_write: 0x11117a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11127a, value : 32'hba}, //phyinit_io_write: 0x11117b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11127b, value : 32'hba}, //phyinit_io_write: 0x11127a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11137a, value : 32'hba}, //phyinit_io_write: 0x11127b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11137b, value : 32'hba}, //phyinit_io_write: 0x11137a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11147a, value : 32'hba}, //phyinit_io_write: 0x11137b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11147b, value : 32'hba}, //phyinit_io_write: 0x11147a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11157a, value : 32'hba}, //phyinit_io_write: 0x11147b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11157b, value : 32'hba}, //phyinit_io_write: 0x11157a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11167a, value : 32'hba}, //phyinit_io_write: 0x11157b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11167b, value : 32'hba}, //phyinit_io_write: 0x11167a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11177a, value : 32'hba}, //phyinit_io_write: 0x11167b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11177b, value : 32'hba}, //phyinit_io_write: 0x11177a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11187a, value : 32'hba}, //phyinit_io_write: 0x11177b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11187b, value : 32'hba}, //phyinit_io_write: 0x11187a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11207a, value : 32'hba}, //phyinit_io_write: 0x11187b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11207b, value : 32'hba}, //phyinit_io_write: 0x11207a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11217a, value : 32'hba}, //phyinit_io_write: 0x11207b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11217b, value : 32'hba}, //phyinit_io_write: 0x11217a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11227a, value : 32'hba}, //phyinit_io_write: 0x11217b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11227b, value : 32'hba}, //phyinit_io_write: 0x11227a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11237a, value : 32'hba}, //phyinit_io_write: 0x11227b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11237b, value : 32'hba}, //phyinit_io_write: 0x11237a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11247a, value : 32'hba}, //phyinit_io_write: 0x11237b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11247b, value : 32'hba}, //phyinit_io_write: 0x11247a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11257a, value : 32'hba}, //phyinit_io_write: 0x11247b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11257b, value : 32'hba}, //phyinit_io_write: 0x11257a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11267a, value : 32'hba}, //phyinit_io_write: 0x11257b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11267b, value : 32'hba}, //phyinit_io_write: 0x11267a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11277a, value : 32'hba}, //phyinit_io_write: 0x11267b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11277b, value : 32'hba}, //phyinit_io_write: 0x11277a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11287a, value : 32'hba}, //phyinit_io_write: 0x11277b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11287b, value : 32'hba}, //phyinit_io_write: 0x11287a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11307a, value : 32'hba}, //phyinit_io_write: 0x11287b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11307b, value : 32'hba}, //phyinit_io_write: 0x11307a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11317a, value : 32'hba}, //phyinit_io_write: 0x11307b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11317b, value : 32'hba}, //phyinit_io_write: 0x11317a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11327a, value : 32'hba}, //phyinit_io_write: 0x11317b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11327b, value : 32'hba}, //phyinit_io_write: 0x11327a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11337a, value : 32'hba}, //phyinit_io_write: 0x11327b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11337b, value : 32'hba}, //phyinit_io_write: 0x11337a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11347a, value : 32'hba}, //phyinit_io_write: 0x11337b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11347b, value : 32'hba}, //phyinit_io_write: 0x11347a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11357a, value : 32'hba}, //phyinit_io_write: 0x11347b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11357b, value : 32'hba}, //phyinit_io_write: 0x11357a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11367a, value : 32'hba}, //phyinit_io_write: 0x11357b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11367b, value : 32'hba}, //phyinit_io_write: 0x11367a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11377a, value : 32'hba}, //phyinit_io_write: 0x11367b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11377b, value : 32'hba}, //phyinit_io_write: 0x11377a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11387a, value : 32'hba}, //phyinit_io_write: 0x11377b, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h11387b, value : 32'hba}, //phyinit_io_write: 0x11387a, 0xba
                          '{ step_type : REG_WRITE, reg_addr : 32'h110078, value : 32'h352}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming RxDigStrbDlyTg0/Tg1 to 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110079, value : 32'h352}, //phyinit_io_write: 0x110078, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110178, value : 32'h352}, //phyinit_io_write: 0x110079, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110179, value : 32'h352}, //phyinit_io_write: 0x110178, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110278, value : 32'h352}, //phyinit_io_write: 0x110179, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110279, value : 32'h352}, //phyinit_io_write: 0x110278, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110378, value : 32'h352}, //phyinit_io_write: 0x110279, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110379, value : 32'h352}, //phyinit_io_write: 0x110378, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110478, value : 32'h352}, //phyinit_io_write: 0x110379, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110479, value : 32'h352}, //phyinit_io_write: 0x110478, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110578, value : 32'h352}, //phyinit_io_write: 0x110479, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110579, value : 32'h352}, //phyinit_io_write: 0x110578, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110678, value : 32'h352}, //phyinit_io_write: 0x110579, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110679, value : 32'h352}, //phyinit_io_write: 0x110678, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110778, value : 32'h352}, //phyinit_io_write: 0x110679, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110779, value : 32'h352}, //phyinit_io_write: 0x110778, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110878, value : 32'h352}, //phyinit_io_write: 0x110779, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110879, value : 32'h352}, //phyinit_io_write: 0x110878, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111078, value : 32'h352}, //phyinit_io_write: 0x110879, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111079, value : 32'h352}, //phyinit_io_write: 0x111078, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111178, value : 32'h352}, //phyinit_io_write: 0x111079, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111179, value : 32'h352}, //phyinit_io_write: 0x111178, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111278, value : 32'h352}, //phyinit_io_write: 0x111179, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111279, value : 32'h352}, //phyinit_io_write: 0x111278, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111378, value : 32'h352}, //phyinit_io_write: 0x111279, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111379, value : 32'h352}, //phyinit_io_write: 0x111378, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111478, value : 32'h352}, //phyinit_io_write: 0x111379, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111479, value : 32'h352}, //phyinit_io_write: 0x111478, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111578, value : 32'h352}, //phyinit_io_write: 0x111479, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111579, value : 32'h352}, //phyinit_io_write: 0x111578, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111678, value : 32'h352}, //phyinit_io_write: 0x111579, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111679, value : 32'h352}, //phyinit_io_write: 0x111678, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111778, value : 32'h352}, //phyinit_io_write: 0x111679, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111779, value : 32'h352}, //phyinit_io_write: 0x111778, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111878, value : 32'h352}, //phyinit_io_write: 0x111779, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h111879, value : 32'h352}, //phyinit_io_write: 0x111878, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112078, value : 32'h352}, //phyinit_io_write: 0x111879, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112079, value : 32'h352}, //phyinit_io_write: 0x112078, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112178, value : 32'h352}, //phyinit_io_write: 0x112079, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112179, value : 32'h352}, //phyinit_io_write: 0x112178, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112278, value : 32'h352}, //phyinit_io_write: 0x112179, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112279, value : 32'h352}, //phyinit_io_write: 0x112278, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112378, value : 32'h352}, //phyinit_io_write: 0x112279, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112379, value : 32'h352}, //phyinit_io_write: 0x112378, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112478, value : 32'h352}, //phyinit_io_write: 0x112379, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112479, value : 32'h352}, //phyinit_io_write: 0x112478, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112578, value : 32'h352}, //phyinit_io_write: 0x112479, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112579, value : 32'h352}, //phyinit_io_write: 0x112578, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112678, value : 32'h352}, //phyinit_io_write: 0x112579, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112679, value : 32'h352}, //phyinit_io_write: 0x112678, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112778, value : 32'h352}, //phyinit_io_write: 0x112679, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112779, value : 32'h352}, //phyinit_io_write: 0x112778, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112878, value : 32'h352}, //phyinit_io_write: 0x112779, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h112879, value : 32'h352}, //phyinit_io_write: 0x112878, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113078, value : 32'h352}, //phyinit_io_write: 0x112879, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113079, value : 32'h352}, //phyinit_io_write: 0x113078, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113178, value : 32'h352}, //phyinit_io_write: 0x113079, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113179, value : 32'h352}, //phyinit_io_write: 0x113178, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113278, value : 32'h352}, //phyinit_io_write: 0x113179, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113279, value : 32'h352}, //phyinit_io_write: 0x113278, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113378, value : 32'h352}, //phyinit_io_write: 0x113279, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113379, value : 32'h352}, //phyinit_io_write: 0x113378, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113478, value : 32'h352}, //phyinit_io_write: 0x113379, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113479, value : 32'h352}, //phyinit_io_write: 0x113478, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113578, value : 32'h352}, //phyinit_io_write: 0x113479, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113579, value : 32'h352}, //phyinit_io_write: 0x113578, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113678, value : 32'h352}, //phyinit_io_write: 0x113579, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113679, value : 32'h352}, //phyinit_io_write: 0x113678, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113778, value : 32'h352}, //phyinit_io_write: 0x113679, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113779, value : 32'h352}, //phyinit_io_write: 0x113778, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113878, value : 32'h352}, //phyinit_io_write: 0x113779, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h113879, value : 32'h352}, //phyinit_io_write: 0x113878, 0x352
                          '{ step_type : REG_WRITE, reg_addr : 32'h110020, value : 32'h2b3}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming RxEnDlyTg0/Tg1 to 0x2b3
                          '{ step_type : REG_WRITE, reg_addr : 32'h110021, value : 32'h2b3}, //phyinit_io_write: 0x110020, 0x2b3
                          '{ step_type : REG_WRITE, reg_addr : 32'h111020, value : 32'h2b3}, //phyinit_io_write: 0x110021, 0x2b3
                          '{ step_type : REG_WRITE, reg_addr : 32'h111021, value : 32'h2b3}, //phyinit_io_write: 0x111020, 0x2b3
                          '{ step_type : REG_WRITE, reg_addr : 32'h112020, value : 32'h2b3}, //phyinit_io_write: 0x111021, 0x2b3
                          '{ step_type : REG_WRITE, reg_addr : 32'h112021, value : 32'h2b3}, //phyinit_io_write: 0x112020, 0x2b3
                          '{ step_type : REG_WRITE, reg_addr : 32'h113020, value : 32'h2b3}, //phyinit_io_write: 0x112021, 0x2b3
                          '{ step_type : REG_WRITE, reg_addr : 32'h113021, value : 32'h2b3}, //phyinit_io_write: 0x113020, 0x2b3
                          '{ step_type : REG_WRITE, reg_addr : 32'h110010, value : 32'h188}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming RxClkT2UIDlyTg0/Tg1 and RxClkC2UIDlyTg0/Tg1 to 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110011, value : 32'h188}, //phyinit_io_write: 0x110010, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110012, value : 32'h188}, //phyinit_io_write: 0x110011, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110013, value : 32'h188}, //phyinit_io_write: 0x110012, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110110, value : 32'h188}, //phyinit_io_write: 0x110013, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110111, value : 32'h188}, //phyinit_io_write: 0x110110, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110112, value : 32'h188}, //phyinit_io_write: 0x110111, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110113, value : 32'h188}, //phyinit_io_write: 0x110112, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110210, value : 32'h188}, //phyinit_io_write: 0x110113, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110211, value : 32'h188}, //phyinit_io_write: 0x110210, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110212, value : 32'h188}, //phyinit_io_write: 0x110211, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110213, value : 32'h188}, //phyinit_io_write: 0x110212, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110310, value : 32'h188}, //phyinit_io_write: 0x110213, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110311, value : 32'h188}, //phyinit_io_write: 0x110310, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110312, value : 32'h188}, //phyinit_io_write: 0x110311, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110313, value : 32'h188}, //phyinit_io_write: 0x110312, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110410, value : 32'h188}, //phyinit_io_write: 0x110313, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110411, value : 32'h188}, //phyinit_io_write: 0x110410, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110412, value : 32'h188}, //phyinit_io_write: 0x110411, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110413, value : 32'h188}, //phyinit_io_write: 0x110412, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110510, value : 32'h188}, //phyinit_io_write: 0x110413, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110511, value : 32'h188}, //phyinit_io_write: 0x110510, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110512, value : 32'h188}, //phyinit_io_write: 0x110511, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110513, value : 32'h188}, //phyinit_io_write: 0x110512, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110610, value : 32'h188}, //phyinit_io_write: 0x110513, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110611, value : 32'h188}, //phyinit_io_write: 0x110610, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110612, value : 32'h188}, //phyinit_io_write: 0x110611, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110613, value : 32'h188}, //phyinit_io_write: 0x110612, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110710, value : 32'h188}, //phyinit_io_write: 0x110613, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110711, value : 32'h188}, //phyinit_io_write: 0x110710, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110712, value : 32'h188}, //phyinit_io_write: 0x110711, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110713, value : 32'h188}, //phyinit_io_write: 0x110712, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110810, value : 32'h188}, //phyinit_io_write: 0x110713, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110811, value : 32'h188}, //phyinit_io_write: 0x110810, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110812, value : 32'h188}, //phyinit_io_write: 0x110811, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h110813, value : 32'h188}, //phyinit_io_write: 0x110812, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111010, value : 32'h188}, //phyinit_io_write: 0x110813, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111011, value : 32'h188}, //phyinit_io_write: 0x111010, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111012, value : 32'h188}, //phyinit_io_write: 0x111011, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111013, value : 32'h188}, //phyinit_io_write: 0x111012, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111110, value : 32'h188}, //phyinit_io_write: 0x111013, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111111, value : 32'h188}, //phyinit_io_write: 0x111110, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111112, value : 32'h188}, //phyinit_io_write: 0x111111, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111113, value : 32'h188}, //phyinit_io_write: 0x111112, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111210, value : 32'h188}, //phyinit_io_write: 0x111113, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111211, value : 32'h188}, //phyinit_io_write: 0x111210, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111212, value : 32'h188}, //phyinit_io_write: 0x111211, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111213, value : 32'h188}, //phyinit_io_write: 0x111212, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111310, value : 32'h188}, //phyinit_io_write: 0x111213, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111311, value : 32'h188}, //phyinit_io_write: 0x111310, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111312, value : 32'h188}, //phyinit_io_write: 0x111311, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111313, value : 32'h188}, //phyinit_io_write: 0x111312, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111410, value : 32'h188}, //phyinit_io_write: 0x111313, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111411, value : 32'h188}, //phyinit_io_write: 0x111410, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111412, value : 32'h188}, //phyinit_io_write: 0x111411, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111413, value : 32'h188}, //phyinit_io_write: 0x111412, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111510, value : 32'h188}, //phyinit_io_write: 0x111413, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111511, value : 32'h188}, //phyinit_io_write: 0x111510, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111512, value : 32'h188}, //phyinit_io_write: 0x111511, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111513, value : 32'h188}, //phyinit_io_write: 0x111512, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111610, value : 32'h188}, //phyinit_io_write: 0x111513, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111611, value : 32'h188}, //phyinit_io_write: 0x111610, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111612, value : 32'h188}, //phyinit_io_write: 0x111611, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111613, value : 32'h188}, //phyinit_io_write: 0x111612, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111710, value : 32'h188}, //phyinit_io_write: 0x111613, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111711, value : 32'h188}, //phyinit_io_write: 0x111710, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111712, value : 32'h188}, //phyinit_io_write: 0x111711, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111713, value : 32'h188}, //phyinit_io_write: 0x111712, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111810, value : 32'h188}, //phyinit_io_write: 0x111713, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111811, value : 32'h188}, //phyinit_io_write: 0x111810, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111812, value : 32'h188}, //phyinit_io_write: 0x111811, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h111813, value : 32'h188}, //phyinit_io_write: 0x111812, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112010, value : 32'h188}, //phyinit_io_write: 0x111813, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112011, value : 32'h188}, //phyinit_io_write: 0x112010, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112012, value : 32'h188}, //phyinit_io_write: 0x112011, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112013, value : 32'h188}, //phyinit_io_write: 0x112012, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112110, value : 32'h188}, //phyinit_io_write: 0x112013, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112111, value : 32'h188}, //phyinit_io_write: 0x112110, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112112, value : 32'h188}, //phyinit_io_write: 0x112111, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112113, value : 32'h188}, //phyinit_io_write: 0x112112, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112210, value : 32'h188}, //phyinit_io_write: 0x112113, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112211, value : 32'h188}, //phyinit_io_write: 0x112210, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112212, value : 32'h188}, //phyinit_io_write: 0x112211, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112213, value : 32'h188}, //phyinit_io_write: 0x112212, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112310, value : 32'h188}, //phyinit_io_write: 0x112213, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112311, value : 32'h188}, //phyinit_io_write: 0x112310, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112312, value : 32'h188}, //phyinit_io_write: 0x112311, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112313, value : 32'h188}, //phyinit_io_write: 0x112312, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112410, value : 32'h188}, //phyinit_io_write: 0x112313, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112411, value : 32'h188}, //phyinit_io_write: 0x112410, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112412, value : 32'h188}, //phyinit_io_write: 0x112411, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112413, value : 32'h188}, //phyinit_io_write: 0x112412, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112510, value : 32'h188}, //phyinit_io_write: 0x112413, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112511, value : 32'h188}, //phyinit_io_write: 0x112510, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112512, value : 32'h188}, //phyinit_io_write: 0x112511, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112513, value : 32'h188}, //phyinit_io_write: 0x112512, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112610, value : 32'h188}, //phyinit_io_write: 0x112513, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112611, value : 32'h188}, //phyinit_io_write: 0x112610, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112612, value : 32'h188}, //phyinit_io_write: 0x112611, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112613, value : 32'h188}, //phyinit_io_write: 0x112612, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112710, value : 32'h188}, //phyinit_io_write: 0x112613, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112711, value : 32'h188}, //phyinit_io_write: 0x112710, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112712, value : 32'h188}, //phyinit_io_write: 0x112711, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112713, value : 32'h188}, //phyinit_io_write: 0x112712, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112810, value : 32'h188}, //phyinit_io_write: 0x112713, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112811, value : 32'h188}, //phyinit_io_write: 0x112810, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112812, value : 32'h188}, //phyinit_io_write: 0x112811, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h112813, value : 32'h188}, //phyinit_io_write: 0x112812, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113010, value : 32'h188}, //phyinit_io_write: 0x112813, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113011, value : 32'h188}, //phyinit_io_write: 0x113010, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113012, value : 32'h188}, //phyinit_io_write: 0x113011, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113013, value : 32'h188}, //phyinit_io_write: 0x113012, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113110, value : 32'h188}, //phyinit_io_write: 0x113013, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113111, value : 32'h188}, //phyinit_io_write: 0x113110, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113112, value : 32'h188}, //phyinit_io_write: 0x113111, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113113, value : 32'h188}, //phyinit_io_write: 0x113112, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113210, value : 32'h188}, //phyinit_io_write: 0x113113, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113211, value : 32'h188}, //phyinit_io_write: 0x113210, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113212, value : 32'h188}, //phyinit_io_write: 0x113211, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113213, value : 32'h188}, //phyinit_io_write: 0x113212, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113310, value : 32'h188}, //phyinit_io_write: 0x113213, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113311, value : 32'h188}, //phyinit_io_write: 0x113310, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113312, value : 32'h188}, //phyinit_io_write: 0x113311, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113313, value : 32'h188}, //phyinit_io_write: 0x113312, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113410, value : 32'h188}, //phyinit_io_write: 0x113313, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113411, value : 32'h188}, //phyinit_io_write: 0x113410, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113412, value : 32'h188}, //phyinit_io_write: 0x113411, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113413, value : 32'h188}, //phyinit_io_write: 0x113412, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113510, value : 32'h188}, //phyinit_io_write: 0x113413, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113511, value : 32'h188}, //phyinit_io_write: 0x113510, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113512, value : 32'h188}, //phyinit_io_write: 0x113511, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113513, value : 32'h188}, //phyinit_io_write: 0x113512, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113610, value : 32'h188}, //phyinit_io_write: 0x113513, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113611, value : 32'h188}, //phyinit_io_write: 0x113610, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113612, value : 32'h188}, //phyinit_io_write: 0x113611, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113613, value : 32'h188}, //phyinit_io_write: 0x113612, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113710, value : 32'h188}, //phyinit_io_write: 0x113613, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113711, value : 32'h188}, //phyinit_io_write: 0x113710, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113712, value : 32'h188}, //phyinit_io_write: 0x113711, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113713, value : 32'h188}, //phyinit_io_write: 0x113712, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113810, value : 32'h188}, //phyinit_io_write: 0x113713, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113811, value : 32'h188}, //phyinit_io_write: 0x113810, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113812, value : 32'h188}, //phyinit_io_write: 0x113811, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h113813, value : 32'h188}, //phyinit_io_write: 0x113812, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h11000c, value : 32'h9a}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming PptWck2DqoCntInvTrn1 to 0x133
                          '{ step_type : REG_WRITE, reg_addr : 32'h11000d, value : 32'h9a}, //phyinit_io_write: 0x11000c, 0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h110014, value : 32'h133}, //phyinit_io_write: 0x11000d, 0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h110015, value : 32'h133}, //phyinit_io_write: 0x110014, 0x133
                          '{ step_type : REG_WRITE, reg_addr : 32'h11100c, value : 32'h9a}, //phyinit_io_write: 0x110015, 0x133
                          '{ step_type : REG_WRITE, reg_addr : 32'h11100d, value : 32'h9a}, //phyinit_io_write: 0x11100c, 0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h111014, value : 32'h133}, //phyinit_io_write: 0x11100d, 0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h111015, value : 32'h133}, //phyinit_io_write: 0x111014, 0x133
                          '{ step_type : REG_WRITE, reg_addr : 32'h11200c, value : 32'h9a}, //phyinit_io_write: 0x111015, 0x133
                          '{ step_type : REG_WRITE, reg_addr : 32'h11200d, value : 32'h9a}, //phyinit_io_write: 0x11200c, 0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h112014, value : 32'h133}, //phyinit_io_write: 0x11200d, 0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h112015, value : 32'h133}, //phyinit_io_write: 0x112014, 0x133
                          '{ step_type : REG_WRITE, reg_addr : 32'h11300c, value : 32'h9a}, //phyinit_io_write: 0x112015, 0x133
                          '{ step_type : REG_WRITE, reg_addr : 32'h11300d, value : 32'h9a}, //phyinit_io_write: 0x11300c, 0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h113014, value : 32'h133}, //phyinit_io_write: 0x11300d, 0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h113015, value : 32'h133}, //phyinit_io_write: 0x113014, 0x133
                          '{ step_type : REG_WRITE, reg_addr : 32'h70077, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming HwtCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h120071, value : 32'h55}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming HMRxReplicaLcdlSeed HMRxSeed to 0x83 HMRxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h100063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC0 Instance0 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h101063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC1 Instance1 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h102063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC2 Instance2 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h103063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC3 Instance3 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h104063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC4 Instance4 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h105063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX0 HMAC5 Instance5 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h107063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC0 Instance7 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h108063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC1 Instance8 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h109063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC2 Instance9 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h10a063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC3 Instance10 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h10b063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC4 Instance11 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c063, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=1, Memclk=600MHz, Programming ACX1 HMAC5 Instance12 HMTxLcdlSeed HMTxSeed to 0x83 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0063, value : 32'h83}, //phyinit_io_write: 0x10c063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0064, value : 32'h83}, //phyinit_io_write: 0x1e0063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e0087, value : 32'h83}, //phyinit_io_write: 0x1e0064, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1063, value : 32'h83}, //phyinit_io_write: 0x1e0087, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1064, value : 32'h83}, //phyinit_io_write: 0x1e1063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e1087, value : 32'h83}, //phyinit_io_write: 0x1e1064, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2063, value : 32'h83}, //phyinit_io_write: 0x1e1087, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2064, value : 32'h83}, //phyinit_io_write: 0x1e2063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e2087, value : 32'h83}, //phyinit_io_write: 0x1e2064, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3063, value : 32'h83}, //phyinit_io_write: 0x1e2087, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3064, value : 32'h83}, //phyinit_io_write: 0x1e3063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e3087, value : 32'h83}, //phyinit_io_write: 0x1e3064, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4063, value : 32'h83}, //phyinit_io_write: 0x1e3087, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4064, value : 32'h83}, //phyinit_io_write: 0x1e4063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e4087, value : 32'h83}, //phyinit_io_write: 0x1e4064, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5063, value : 32'h83}, //phyinit_io_write: 0x1e4087, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5064, value : 32'h83}, //phyinit_io_write: 0x1e5063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e5087, value : 32'h83}, //phyinit_io_write: 0x1e5064, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6063, value : 32'h83}, //phyinit_io_write: 0x1e5087, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6064, value : 32'h83}, //phyinit_io_write: 0x1e6063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e6087, value : 32'h83}, //phyinit_io_write: 0x1e6064, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7063, value : 32'h83}, //phyinit_io_write: 0x1e6087, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7064, value : 32'h83}, //phyinit_io_write: 0x1e7063, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e7087, value : 32'h83}, //phyinit_io_write: 0x1e7064, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h19080a, value : 32'h283}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=1 Programming Seq0bGPR10 to mission mode HMTxLcdlSeed value 0x283
                          '{ step_type : REG_WRITE, reg_addr : 32'h19080b, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=1 Programming Seq0bGPR11 to mission mode HMTxLcdlSeed value 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h190815, value : 32'h283}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=1 Programming Seq0bGPR21 to mission mode HMTxLcdlSeed value 0x283
                          '{ step_type : REG_WRITE, reg_addr : 32'h190816, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=1 Programming Seq0bGPR22 to mission mode HMTxLcdlSeed value 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h11015f, value : 32'h83}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=1, Memclk=600MHz, Programming RDqRDqsCntrl to 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h11115f, value : 32'h83}, //phyinit_io_write: 0x11015f, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h11215f, value : 32'h83}, //phyinit_io_write: 0x11115f, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h11315f, value : 32'h83}, //phyinit_io_write: 0x11215f, 0x83
                          '{ step_type : REG_WRITE, reg_addr : 32'h160009, value : 32'h10}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Memclk=600MHz, Programming CPllDacValIn to 0x10
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE0.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102a1, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE0.RxReplicaPathPhase1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102a2, value : 32'h2c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE0.RxReplicaPathPhase2 to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102a3, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE0.RxReplicaPathPhase3 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102a4, value : 32'hb7}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE0.RxReplicaPathPhase4 to 0xb7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1112a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE1.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1112a1, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE1.RxReplicaPathPhase1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1112a2, value : 32'h2c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE1.RxReplicaPathPhase2 to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h1112a3, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE1.RxReplicaPathPhase3 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h1112a4, value : 32'hb7}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE1.RxReplicaPathPhase4 to 0xb7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1122a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE2.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1122a1, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE2.RxReplicaPathPhase1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1122a2, value : 32'h2c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE2.RxReplicaPathPhase2 to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h1122a3, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE2.RxReplicaPathPhase3 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h1122a4, value : 32'hb7}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE2.RxReplicaPathPhase4 to 0xb7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1132a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE3.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1132a1, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE3.RxReplicaPathPhase1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1132a2, value : 32'h2c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE3.RxReplicaPathPhase2 to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h1132a3, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE3.RxReplicaPathPhase3 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h1132a4, value : 32'hb7}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE3.RxReplicaPathPhase4 to 0xb7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102ad, value : 32'h2}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE0.RxReplicaCtl01::RxReplicaSelPathPhase to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h1112ad, value : 32'h2}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE1.RxReplicaCtl01::RxReplicaSelPathPhase to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h1122ad, value : 32'h2}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE2.RxReplicaCtl01::RxReplicaSelPathPhase to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h1132ad, value : 32'h2}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE3.RxReplicaCtl01::RxReplicaSelPathPhase to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102af, value : 32'h28}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE0.RxReplicaCtl03 to 0x28
                          '{ step_type : REG_WRITE, reg_addr : 32'h1112af, value : 32'h28}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE1.RxReplicaCtl03 to 0x28
                          '{ step_type : REG_WRITE, reg_addr : 32'h1122af, value : 32'h28}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE2.RxReplicaCtl03 to 0x28
                          '{ step_type : REG_WRITE, reg_addr : 32'h1132af, value : 32'h28}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming DBYTE3.RxReplicaCtl03 to 0x28
                          '{ step_type : REG_WRITE, reg_addr : 32'h190807, value : 32'h9701}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming Seq0BGPR7 to save ZQCalCodeOvrValPU=0x12e and ZQCalCodeOvrEnPU=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h190808, value : 32'hb681}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=1, Programming Seq0BGPR8 to save ZQCalCodeOvrValPD=0x16d and ZQCalCodeOvrEnPD=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h0} //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
//[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] End of dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop(), PState=1
   },
                  
// [dwc_ddrphy_phyinit_userCustom_E_setDfiClk] Start of dwc_ddrphy_phyinit_userCustom_E_setDfiClk()
// [dwc_ddrphy_phyinit_userCustom_E_setDfiClk] End of dwc_ddrphy_phyinit_userCustom_E_setDfiClk()
 
   "F" : '{                 
// [dwc_ddrphy_phyinit_F_loadDMEM1D] Start of dwc_ddrphy_phyinit_F_loadDMEM (pstate=1, Train2D=0)
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0088, value : 32'h1}, //[dwc_ddrphy_phyinit_F_loadDMEM] Program csr StartDccmClear to 1 to clear DCCM.
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 8300},
//Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 8300 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0088, value : 32'h0}, //[dwc_ddrphy_phyinit_F_loadDMEM] Program csr StartDccmClear to 0 after DCCM clear is done.
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}, //Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 40 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'h58000, value : 32'h600}, // [dwc_ddrphy_phyinit_WriteOutMem] STARTING. offset 0x58000 size 0x6000, sparse_write=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h58001, value : 32'h12c00011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58002, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58004, value : 32'hff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58005, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58009, value : 32'h310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5800f, value : 32'h10000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58010, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58016, value : 32'h80800000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58017, value : 32'h88888080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58018, value : 32'he0e8888},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58019, value : 32'h54540e0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801a, value : 32'h44445454},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801b, value : 32'h50504444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801c, value : 32'h5050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801d, value : 32'h50500000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801e, value : 32'h50505050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801f, value : 32'h5050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58020, value : 32'hac840000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58021, value : 32'hac84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58023, value : 32'h2020000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58024, value : 32'h202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5802a, value : 32'h4040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5802b, value : 32'h404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58032, value : 32'h60600000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58033, value : 32'h6060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58048, value : 32'h2b000001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58049, value : 32'h27},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58054, value : 32'h5c0032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58055, value : 32'he000b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58056, value : 32'h164013a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58057, value : 32'h1e801be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58062, value : 32'h6400c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58103, value : 32'h50b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58104, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58108, value : 32'h8080808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58110, value : 32'hef0f4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811b, value : 32'h4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811d, value : 32'h40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811e, value : 32'h180f0e0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811f, value : 32'h4746451e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58120, value : 32'h4a4948},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58121, value : 32'h1000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58125, value : 32'h40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58126, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58129, value : 32'hffffffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5812e, value : 32'h2f059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5812f, value : 32'hffb50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58130, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58131, value : 32'h1f0b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58132, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58133, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58134, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58135, value : 32'hf0b00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58136, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58137, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58138, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58139, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813a, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813b, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813c, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813d, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813e, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813f, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58140, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58141, value : 32'hff740182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58142, value : 32'h800001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58143, value : 32'h1ffbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58144, value : 32'hf0be0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58145, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58146, value : 32'h1f0a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58147, value : 32'hf0a20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58148, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58149, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814a, value : 32'h40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814b, value : 32'h308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814c, value : 32'h560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814e, value : 32'h80000dbc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814f, value : 32'h309},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58150, value : 32'h561},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58151, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58152, value : 32'h80000dcd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58153, value : 32'he0305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58154, value : 32'he0205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58155, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58156, value : 32'h80000dde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58157, value : 32'he0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58158, value : 32'he0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58159, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815a, value : 32'h80000e44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815b, value : 32'he0301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815c, value : 32'he0201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815d, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815e, value : 32'h80000e57},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815f, value : 32'he0302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58160, value : 32'he0202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58161, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58162, value : 32'h80000e6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58163, value : 32'he0303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58164, value : 32'he0203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58165, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58166, value : 32'h80000e7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58167, value : 32'he0304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58168, value : 32'he0204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58169, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816a, value : 32'h80000e90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816b, value : 32'h1ff01ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816c, value : 32'he0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816e, value : 32'h63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816f, value : 32'h64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58170, value : 32'h660},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58172, value : 32'h80000d8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58173, value : 32'h661},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58174, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58175, value : 32'h80000dad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58176, value : 32'he00f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58177, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58178, value : 32'h80000def},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58179, value : 32'he00f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817a, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817b, value : 32'h80000e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817c, value : 32'he00f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817d, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817e, value : 32'h80000e11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817f, value : 32'he00f3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58180, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58181, value : 32'h80000e22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58182, value : 32'he00f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58183, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58184, value : 32'h80000e33},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58185, value : 32'he00f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58186, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58187, value : 32'h80000d9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58188, value : 32'h2011210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58189, value : 32'h1c0a1403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818a, value : 32'hb112e29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818b, value : 32'h1916150d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818c, value : 32'h180f0e0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818d, value : 32'h453a131e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818e, value : 32'h49484746},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818f, value : 32'h2006e4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58190, value : 32'h100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58191, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58192, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58194, value : 32'h2150001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58195, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58196, value : 32'h1010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58197, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58198, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58199, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819a, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819b, value : 32'h6400002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819c, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819d, value : 32'h30215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819e, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819f, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a0, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a1, value : 32'h10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a2, value : 32'habe0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a3, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a4, value : 32'h50320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a5, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c5, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c6, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c7, value : 32'h43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c8, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c9, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ca, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cb, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cc, value : 32'h42b0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cd, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ce, value : 32'h200c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cf, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d0, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d1, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d2, value : 32'h10003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d3, value : 32'h8550002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d4, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d5, value : 32'h40158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d6, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d7, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d8, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d9, value : 32'h10005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581da, value : 32'hc800002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581db, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581dc, value : 32'h601d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581dd, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581de, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581df, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e0, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e1, value : 32'h10ab0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e2, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e3, value : 32'h80258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e4, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e5, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e6, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e7, value : 32'h20009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e8, value : 32'h157c0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e9, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ea, value : 32'ha02ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581eb, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ec, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ed, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ee, value : 32'h2000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ef, value : 32'h19000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f0, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f1, value : 32'hc03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f2, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f3, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f4, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f5, value : 32'h3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f6, value : 32'h21550006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f7, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f8, value : 32'he04b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f9, value : 32'h70003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fa, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fb, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fc, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fd, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fe, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ff, value : 32'h2150004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58200, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58201, value : 32'h4010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58202, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58203, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58204, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58205, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58206, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58207, value : 32'h80006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58208, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58209, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820a, value : 32'h6400006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820b, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820c, value : 32'h80215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820d, value : 32'h2000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820e, value : 32'h30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820f, value : 32'h70004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58210, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58211, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58212, value : 32'he0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58213, value : 32'h70001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58214, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58215, value : 32'habe0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58216, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58217, value : 32'ha0320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58218, value : 32'h30010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58219, value : 32'h40009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5821a, value : 32'h80004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824c, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824d, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824e, value : 32'h20043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824f, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58250, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58251, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58252, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58253, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58254, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58255, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58256, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58257, value : 32'h42b0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58258, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58259, value : 32'h300c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825a, value : 32'h10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825b, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825c, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825d, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825e, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825f, value : 32'h50004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58260, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58261, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58262, value : 32'h8550004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58263, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58264, value : 32'h40158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58265, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58266, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58267, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58268, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58269, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826a, value : 32'h80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826b, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826c, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826d, value : 32'hc800004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826e, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826f, value : 32'h601d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58270, value : 32'h20009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58271, value : 32'h30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58272, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58273, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58274, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58275, value : 32'hb0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58276, value : 32'h70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58277, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58278, value : 32'h10ab0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58279, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827a, value : 32'h70258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827b, value : 32'h3000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827c, value : 32'h30008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827d, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827e, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827f, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58280, value : 32'he0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58281, value : 32'h90003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58282, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58283, value : 32'h157c0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58284, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58285, value : 32'h902ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58286, value : 32'h4000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58287, value : 32'h4000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58288, value : 32'h60002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58289, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828a, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828b, value : 32'h100009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828c, value : 32'hb0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828d, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828e, value : 32'h19000006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828f, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58290, value : 32'hb03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58291, value : 32'h50013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58292, value : 32'h5000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58293, value : 32'h70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58294, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58295, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58296, value : 32'h16000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58297, value : 32'hf0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58298, value : 32'h20006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58299, value : 32'h21550008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829a, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829b, value : 32'he04b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829c, value : 32'h60018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829d, value : 32'h70010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829e, value : 32'h90002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829f, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a0, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a1, value : 32'h60006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a2, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a4, value : 32'h60001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a5, value : 32'h2150007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a6, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a7, value : 32'h8010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a8, value : 32'h80008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582aa, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ab, value : 32'h90007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ac, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ad, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ae, value : 32'ha000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582af, value : 32'h1000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b0, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b1, value : 32'h80002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b2, value : 32'h640000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b3, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b4, value : 32'hc0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b5, value : 32'he000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b6, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b7, value : 32'h30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b8, value : 32'hb0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b9, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ba, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bb, value : 32'h100010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bc, value : 32'h30012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bd, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582be, value : 32'ha0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bf, value : 32'habe000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c0, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c1, value : 32'h120320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c2, value : 32'h140014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c3, value : 32'h70005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c4, value : 32'h40007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c5, value : 32'he000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58300, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58301, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58302, value : 32'h30043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58303, value : 32'h30003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58305, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58306, value : 32'h40003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58307, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58308, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58309, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830a, value : 32'h4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830c, value : 32'h40001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830d, value : 32'h42b0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830e, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830f, value : 32'h500c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58310, value : 32'h50005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58311, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58312, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58313, value : 32'h50004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58314, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58315, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58316, value : 32'h70006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58317, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58318, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58319, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831a, value : 32'h8550006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831b, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831c, value : 32'h80158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831d, value : 32'h90008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831e, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831f, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58320, value : 32'h70005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58321, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58322, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58323, value : 32'ha0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58324, value : 32'h3000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58325, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58326, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58327, value : 32'hc800007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58328, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58329, value : 32'ha01d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832a, value : 32'hc000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832b, value : 32'h40003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832c, value : 32'h30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832d, value : 32'h80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832e, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832f, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58330, value : 32'hd000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58331, value : 32'h4000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58332, value : 32'h60005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58333, value : 32'h60003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58334, value : 32'h10ab0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58335, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58336, value : 32'hd0258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58337, value : 32'hf000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58338, value : 32'h60005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58339, value : 32'h30007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833a, value : 32'h90006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833b, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833c, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833d, value : 32'h10000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833e, value : 32'h60011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833f, value : 32'h80007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58340, value : 32'h60004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58341, value : 32'h157c000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58342, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58343, value : 32'h1002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58344, value : 32'h130011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58345, value : 32'h70006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58346, value : 32'h40009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58347, value : 32'hb0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58348, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58349, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834a, value : 32'h120011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834b, value : 32'h70014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834c, value : 32'ha0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834d, value : 32'h70004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834e, value : 32'h1900000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834f, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58350, value : 32'h1403aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58351, value : 32'h180016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58352, value : 32'h90007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58353, value : 32'h5000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58354, value : 32'he0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58355, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58356, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58357, value : 32'h190017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58358, value : 32'h8001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58359, value : 32'hb000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835a, value : 32'ha0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835b, value : 32'h21550010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835c, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835d, value : 32'h1904b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835e, value : 32'h1d001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835f, value : 32'hb0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58360, value : 32'h7000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58361, value : 32'h12000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58362, value : 32'ha05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58363, value : 32'h50000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58364, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58365, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58366, value : 32'h43416564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58367, value : 32'h63500030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58368, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58369, value : 32'h646f4341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836a, value : 32'h53514465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836b, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836c, value : 32'h4143446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836d, value : 32'h65646f43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836e, value : 32'h314341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836f, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58370, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58371, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58372, value : 32'h30434174},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58373, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58374, value : 32'h4443446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58375, value : 32'h7366664f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58376, value : 32'h43417465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58377, value : 32'h63500031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58378, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58379, value : 32'h66664f44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837a, value : 32'h44746573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837b, value : 32'h50005351},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837c, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837d, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837e, value : 32'h71446564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837f, value : 32'h306e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58380, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58381, value : 32'h43414344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58382, value : 32'h4465646f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58383, value : 32'h316e4c71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58384, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58385, value : 32'h4143446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58386, value : 32'h65646f43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58387, value : 32'h6e4c7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58388, value : 32'h63500032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58389, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838a, value : 32'h646f4341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838b, value : 32'h4c714465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838c, value : 32'h5000336e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838d, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838e, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838f, value : 32'h71446564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58390, value : 32'h346e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58391, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58392, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58393, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58394, value : 32'h4c714474},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58395, value : 32'h5000306e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58396, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58397, value : 32'h664f4443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58398, value : 32'h74657366},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58399, value : 32'h6e4c7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839a, value : 32'h63500031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839b, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839c, value : 32'h66664f44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839d, value : 32'h44746573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839e, value : 32'h326e4c71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839f, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a0, value : 32'h4443446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a1, value : 32'h7366664f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a2, value : 32'h71447465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a3, value : 32'h336e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a4, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a5, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a6, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a7, value : 32'h4c714474},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a8, value : 32'h346e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a9, value : 32'h4050607},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583aa, value : 32'h10203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ab, value : 32'hc0b0a09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ac, value : 32'hb50f0e0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ad, value : 32'h1ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ae, value : 32'h1f0b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583af, value : 32'hb3000100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b0, value : 32'h1f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b1, value : 32'h1f0b400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b2, value : 32'hb0000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b3, value : 32'h300001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b4, value : 32'h7f00300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b5, value : 32'h4000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b6, value : 32'h7f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b7, value : 32'h1fe0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b8, value : 32'h4000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b9, value : 32'h1fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ba, value : 32'h7f01100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bb, value : 32'h21000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bc, value : 32'h1fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bd, value : 32'h1ffbe00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583be, value : 32'hbe000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bf, value : 32'h10001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c0, value : 32'h1f0a700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c1, value : 32'ha2000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c2, value : 32'h20001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c3, value : 32'h2007900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c4, value : 32'h4000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c5, value : 32'h1008b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c6, value : 32'hf05f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c7, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c8, value : 32'h1ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c9, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ca, value : 32'h1ff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cb, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cc, value : 32'hf0b001ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cd, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ce, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cf, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d0, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d1, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d2, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d3, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d4, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d5, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d6, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d7, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d8, value : 32'hf0a70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d9, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583da, value : 32'he000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583db, value : 32'hc000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583dc, value : 32'ha000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583dd, value : 32'h80009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583de, value : 32'h60007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583df, value : 32'h40005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e0, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e1, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e2, value : 32'h110010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e3, value : 32'h130012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e4, value : 32'h150014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e5, value : 32'h170016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e6, value : 32'h190018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e7, value : 32'h1b001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e8, value : 32'h1d001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e9, value : 32'h1f001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ea, value : 32'hef77dbb7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583eb, value : 32'hfbdff7bd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ec, value : 32'hbddfb76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ed, value : 32'hbdffbdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ee, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ef, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f0, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f1, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f2, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f3, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f4, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f5, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f6, value : 32'h1ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f7, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f8, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f9, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fa, value : 32'hf0b90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fb, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fc, value : 32'h1f0ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fd, value : 32'hf0b10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fe, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ff, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58400, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58401, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58402, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58403, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58404, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58405, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58406, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58407, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58408, value : 32'h7f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58409, value : 32'hfe200002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840a, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840b, value : 32'h7f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840c, value : 32'hf01cffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840d, value : 32'hffff0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840e, value : 32'h1fe2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840f, value : 32'hfe2bffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58410, value : 32'hffff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58411, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58412, value : 32'hffb50040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58413, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58414, value : 32'h1f0b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58415, value : 32'hf0b40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58416, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58417, value : 32'h1f0b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58418, value : 32'hf0ba0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58419, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841a, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841b, value : 32'hf0b00002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841c, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841d, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841e, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841f, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58420, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58421, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58422, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58423, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58424, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58425, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58426, value : 32'h7f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58427, value : 32'hfe200002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58428, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58429, value : 32'h7f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842a, value : 32'hf01cffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842b, value : 32'hffff0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842c, value : 32'h1fe2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842d, value : 32'hfe2bffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842e, value : 32'hffff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842f, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58430, value : 32'h40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58431, value : 32'h8840884},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58432, value : 32'h20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58433, value : 32'h10010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58434, value : 32'h10012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58435, value : 32'h1007a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58436, value : 32'h10028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58437, value : 32'h60000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58438, value : 32'h50005000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58439, value : 32'h2008050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843b, value : 32'h60080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843c, value : 32'h3c5a5555},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843d, value : 32'h600000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58440, value : 32'h70},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58441, value : 32'h75},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58442, value : 32'h26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58443, value : 32'ha0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58444, value : 32'ha1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58445, value : 32'ha4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58446, value : 32'ha5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58447, value : 32'ha030201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58448, value : 32'he0d0c0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58449, value : 32'h1413120f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844a, value : 32'h18171615},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844b, value : 32'h1e1c1a19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844c, value : 32'h2221201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844d, value : 32'h2e292825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844e, value : 32'h4746453a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844f, value : 32'h4a4948},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1} //This allows the firmware unrestricted access to the configuration CSRs.
//[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
// [dwc_ddrphy_phyinit_F_loadDMEM1D] End of dwc_ddrphy_phyinit_F_loadDMEM, Pstate=1
   },
   "G" : '{                 
// [dwc_ddrphy_phyinit_G_execFW] Start of dwc_ddrphy_phyinit_G_execFW
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1}, ////     Then rewrite the CSR so that only the StallToMicro remains set (all other fields should be zero).
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h9}, //[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h0}, // [dwc_ddrphy_phyinit_userCustom_G_waitFwDone] Start of dwc_ddrphy_phyinit_userCustom_G_waitFwDone()
// [dwc_ddrphy_phyinit_userCustom_G_waitFwDone] End of dwc_ddrphy_phyinit_userCustom_G_waitFwDone()
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h1}, //// 4.   Halt the microcontroller."
// [dwc_ddrphy_phyinit_G_execFW] End of dwc_ddrphy_phyinit_G_execFW
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}    },
                  
// [dwc_ddrphy_phyinit_userCustom_H_readMsgBlock] Start of dwc_ddrphy_phyinit_userCustom_H_readMsgBlock()
// [dwc_ddrphy_phyinit_userCustom_H_readMsgBlock] End of dwc_ddrphy_phyinit_userCustom_H_readMsgBlock ()
// 3. If training is required at another frequency, repeat the operations starting at step (E).
// [dwc_ddrphy_phyinit_H_readMsgBlock] End of dwc_ddrphy_phyinit_H_readMsgBlock
 
   "I" : '{                 
//[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Start of dwc_ddrphy_phyinit_I_loadPIEImagePsLoop(), PState=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h160008, value : 32'h956}, //[dwc_ddrphy_phyinit_programPLL] [phyinit_I_loadPIEImagePsLoop] Pstate=1,  Memclk=600MHz, Programming CpllCtrl5 to 0x956.
                          '{ step_type : REG_WRITE, reg_addr : 32'h60006, value : 32'h3f0}, //End of dwc_ddrphy_phyinit_programPLL(), PState=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h130015, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h131015, value : 32'h0}, //phyinit_io_write: 0x130015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11007c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11107c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11207c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11307c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11007c, value : 32'h0}, //phyinit_io_write: 0x11307c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11107c, value : 32'h0}, //phyinit_io_write: 0x11007c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11207c, value : 32'h0}, //phyinit_io_write: 0x11107c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11307c, value : 32'h0}, //phyinit_io_write: 0x11207c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h130015, value : 32'h0}, //phyinit_io_write: 0x11307c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h131015, value : 32'h0}, //phyinit_io_write: 0x130015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h170141, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming ACSMWckFreeRunMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h19080c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming GPR12 with Zcalkclkdiv to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h110027, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming RxClkCntl1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h111027, value : 32'h0}, //phyinit_io_write: 0x110027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h112027, value : 32'h0}, //phyinit_io_write: 0x111027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h113027, value : 32'h0}, //phyinit_io_write: 0x112027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11020f, value : 32'h8}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=1, Programming RxReplicaCtl04 to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h11120f, value : 32'h8}, //phyinit_io_write: 0x11020f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h11220f, value : 32'h8}, //phyinit_io_write: 0x11120f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h11320f, value : 32'h8}, //phyinit_io_write: 0x11220f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e003f, value : 32'h0}, //phyinit_io_write: 0x11320f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e008d, value : 32'h0}, //phyinit_io_write: 0x1e003f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e103f, value : 32'h0}, //phyinit_io_write: 0x1e008d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e108d, value : 32'h0}, //phyinit_io_write: 0x1e103f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e203f, value : 32'h0}, //phyinit_io_write: 0x1e108d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e208d, value : 32'h0}, //phyinit_io_write: 0x1e203f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e303f, value : 32'h0}, //phyinit_io_write: 0x1e208d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e308d, value : 32'h0}, //phyinit_io_write: 0x1e303f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e403f, value : 32'h0}, //phyinit_io_write: 0x1e308d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e408d, value : 32'h0}, //phyinit_io_write: 0x1e403f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e503f, value : 32'h0}, //phyinit_io_write: 0x1e408d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e508d, value : 32'h0}, //phyinit_io_write: 0x1e503f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e603f, value : 32'h0}, //phyinit_io_write: 0x1e508d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e608d, value : 32'h0}, //phyinit_io_write: 0x1e603f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e703f, value : 32'h0}, //phyinit_io_write: 0x1e608d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1e708d, value : 32'h0}, //phyinit_io_write: 0x1e703f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h190903, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] PState=1, Programming RtrnMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70072, value : 32'h3}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming HwtLpCsEnA to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h19080e, value : 32'h3}, //phyinit_io_write: 0x70072, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h70073, value : 32'h3}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming HwtLpCsEnB to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h19080f, value : 32'h3}, //phyinit_io_write: 0x70073, 0x3
//phyinit_io_write: 0x19080f, 0x3
//[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] End of dwc_ddrphy_phyinit_I_loadPIEImagePsLoop(), PState=1
//[dwc_ddrphy_phyinit_userCustom_customPostTrainPsLoop] End of dwc_ddrphy_phyinit_userCustom_customPostTrainPsLoop(), PState=1
//Start of dwc_ddrphy_phyinit_C_initPhyConfigPsLoop(), PState=2, tck_ps=2500ps
                          '{ step_type : REG_WRITE, reg_addr : 32'h2008b, value : 32'h2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, programming PState = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h290801, value : 32'ha692}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming Seq0BGPR1 to 0xa692
                          '{ step_type : REG_WRITE, reg_addr : 32'h290802, value : 32'h0}, //phyinit_io_write: 0x290801, 0xa692
                          '{ step_type : REG_WRITE, reg_addr : 32'h290806, value : 32'h1}, //phyinit_io_write: 0x290802, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2a03ff, value : 32'h4101}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming OdtSeg120 to 0x4101
                          '{ step_type : REG_WRITE, reg_addr : 32'h2a030b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming ZCalCompCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h260008, value : 32'h4a96}, //[dwc_ddrphy_phyinit_programPLL] [phyinit_C_initPhyConfigPsLoop] Pstate=2,  Memclk=400MHz, Programming CpllCtrl5 to 0x4a96.
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908e0, value : 32'h32}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY0 to 0x32 (0.5us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908e1, value : 32'h96}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY1 to 0x96 (tZQCal PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908e2, value : 32'h3e8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY2 to 0x3e8 (10.us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908e3, value : 32'h58}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY3 to 0x58 (dllLock PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908e4, value : 32'ha}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY4 to 0xa (0.1us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908e5, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY5 to 0x0 (RxReplicaCalWait delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908e6, value : 32'h43}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY6 to 0x43 (Oscillator PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908e7, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY7 to 0x0 (tXDSM_XP PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908ea, value : 32'h2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY10 to 0x2 (tPDXCSODTON 20ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908eb, value : 32'h2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY11 to 0x2 (20ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908ec, value : 32'h5}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY12 to 0x5 (50ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h2908ed, value : 32'h27}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming Seq0BDLY13 to 0x27 (tXSR PIE delay, tRFCab delay is 380ns)
                          '{ step_type : REG_WRITE, reg_addr : 32'h220002, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming PclkPtrInitVal to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h260040, value : 32'h3}, //phyinit_io_write: 0x220002, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h220000, value : 32'h2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DfiFreqRatio to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h2100fb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming RxDigStrbEn to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2110fb, value : 32'h0}, //phyinit_io_write: 0x2100fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2120fb, value : 32'h0}, //phyinit_io_write: 0x2110fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2130fb, value : 32'h0}, //phyinit_io_write: 0x2120fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e000b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DxDigStrobeMode HMDBYTE to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e100b, value : 32'h0}, //phyinit_io_write: 0x2e000b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e200b, value : 32'h0}, //phyinit_io_write: 0x2e100b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e300b, value : 32'h0}, //phyinit_io_write: 0x2e200b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e400b, value : 32'h0}, //phyinit_io_write: 0x2e300b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e500b, value : 32'h0}, //phyinit_io_write: 0x2e400b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e600b, value : 32'h0}, //phyinit_io_write: 0x2e500b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e700b, value : 32'h0}, //phyinit_io_write: 0x2e600b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h210024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE0.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h211024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE1.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h212024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE2.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h213024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE3.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h210025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE0.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h211025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE1.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h212025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE2.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h213025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE3.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h210004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE0.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h210003, value : 32'h0}, //phyinit_io_write: 0x210004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h211004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE1.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h211003, value : 32'h0}, //phyinit_io_write: 0x211004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h212004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE2.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h212003, value : 32'h0}, //phyinit_io_write: 0x212004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h213004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE3.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h213003, value : 32'h0}, //phyinit_io_write: 0x213004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2b0004, value : 32'h190}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ZCalClkInfo::ZCalDfiClkTicksPer1uS to 0x190
                          '{ step_type : REG_WRITE, reg_addr : 32'h2a030c, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h21003e, value : 32'h5}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE RxGainCurrAdjRxReplica to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h21103e, value : 32'h5}, //phyinit_io_write: 0x21003e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h21203e, value : 32'h5}, //phyinit_io_write: 0x21103e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h21303e, value : 32'h5}, //phyinit_io_write: 0x21203e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h220003, value : 32'h1}, //phyinit_io_write: 0x21303e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h22000b, value : 32'h1111}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming CPclkDivRatio to 0x1111
                          '{ step_type : REG_WRITE, reg_addr : 32'h210108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE0.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h211108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE1.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h212108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE2.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h213108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming DBYTE3.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70005, value : 32'h0}, //[phyinit_C_initPhyConfig] Programming EnPhyUpdZQCalUpdate to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h7000f, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming DisableZQupdateOnSnoop to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21000e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h21100e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h21200e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h21300e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h220019, value : 32'h4}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming EnRxDqsTracking::DqsSampNegRxEnSense to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e002c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 0 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e102c, value : 32'h33}, //phyinit_io_write: 0x2e002c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e002d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 0 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e102d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 0 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e202c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 1 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e302c, value : 32'h33}, //phyinit_io_write: 0x2e202c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e202d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 1 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e302d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 1 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e402c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 2 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e502c, value : 32'h33}, //phyinit_io_write: 0x2e402c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e402d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 2 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e502d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 2 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e602c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 3 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e702c, value : 32'h33}, //phyinit_io_write: 0x2e602c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e602d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 3 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e702d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 3 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h200070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC0 Instance0 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h201070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC1 Instance1 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h202070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC2 Instance2 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h203070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC3 Instance3 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h204070, value : 32'hff}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming AC0 HMAC4 Instance4 CS TxImpedanceAC::TxStrenCodePDAC to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h205070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC5 Instance5 TxImpedanceAC::TxStrenCodePD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h207070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC0 Instance7 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h208070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC1 Instance8 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h209070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC2 Instance9 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h20a070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC3 Instance10 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h20b070, value : 32'hff}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming AC1 HMAC4 Instance11 CS TxImpedanceAC::TxStrenCodePDAC to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h20c070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC5 Instance12 TxImpedanceAC::TxStrenCodePD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e002e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 0 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e102e, value : 32'h30}, //phyinit_io_write: 0x2e002e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e002f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 0 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e102f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 0 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e202e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 1 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e302e, value : 32'h30}, //phyinit_io_write: 0x2e202e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e202f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 1 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e302f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 1 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e402e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 2 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e502e, value : 32'h30}, //phyinit_io_write: 0x2e402e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e402f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 2 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e502f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 2 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e602e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 3 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e702e, value : 32'h30}, //phyinit_io_write: 0x2e602e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e602f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 3 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e702f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 3 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h200079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC0 Instance0 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h201079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC1 Instance1 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h202079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC2 Instance2 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h203079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC3 Instance3 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h204079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC4 Instance4 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h205079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC5 DIFF5 OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h207079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC0 Instance7 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h208079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC1 Instance8 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h209079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC2 Instance9 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h20a079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC3 Instance10 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h20b079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC4 Instance11 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h20c079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC5 DIFF12 OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e001c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 0 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e101c, value : 32'h3}, //phyinit_io_write: 0x2e001c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e201c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 1 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e301c, value : 32'h3}, //phyinit_io_write: 0x2e201c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e401c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 2 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e501c, value : 32'h3}, //phyinit_io_write: 0x2e401c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e601c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming HMDBYTE 3 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e701c, value : 32'h3}, //phyinit_io_write: 0x2e601c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h20006d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC0 Instance0 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20106d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC1 Instance1 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20206d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC2 Instance2 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20306d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC3 Instance3 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20406d, value : 32'hf8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC4 Instance4 CS TxSlewAC::TxSlewPDAC to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h20506d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX0 HMAC5 Instance5 TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20706d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC0 Instance7 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20806d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC1 Instance8 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20906d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC2 Instance9 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20a06d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC3 Instance10 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20b06d, value : 32'hf8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC4 Instance11 CS TxSlewAC::TxSlewPDAC to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h20c06d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACX1 HMAC5 Instance12 TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e003e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Programming HMDBYTE RxDQSCtrl::RxDQSDiffSeVrefDACEn to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e103e, value : 32'h0}, //phyinit_io_write: 0x2e003e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e203e, value : 32'h0}, //phyinit_io_write: 0x2e103e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e303e, value : 32'h0}, //phyinit_io_write: 0x2e203e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e403e, value : 32'h0}, //phyinit_io_write: 0x2e303e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e503e, value : 32'h0}, //phyinit_io_write: 0x2e403e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e603e, value : 32'h0}, //phyinit_io_write: 0x2e503e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e703e, value : 32'h0}, //phyinit_io_write: 0x2e603e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h210001, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming WriteLinkEcc to 0
                          '{ step_type : REG_WRITE, reg_addr : 32'h211001, value : 32'h0}, //phyinit_io_write: 0x210001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h212001, value : 32'h0}, //phyinit_io_write: 0x211001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h213001, value : 32'h0}, //phyinit_io_write: 0x212001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h270040, value : 32'h5a}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming PPTTrainSetup::PhyMstrMaxReqToAck to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h270041, value : 32'hf}, //phyinit_io_write: 0x270040, 0x5a
                          '{ step_type : REG_WRITE, reg_addr : 32'h2100a5, value : 32'h1}, //phyinit_io_write: 0x270041, 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h2110a5, value : 32'h1}, //phyinit_io_write: 0x2100a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h2120a5, value : 32'h1}, //phyinit_io_write: 0x2110a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h2130a5, value : 32'h1}, //phyinit_io_write: 0x2120a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h210209, value : 32'h3232}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Programming RxReplicaRangeVal 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h211209, value : 32'h3232}, //phyinit_io_write: 0x210209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h212209, value : 32'h3232}, //phyinit_io_write: 0x211209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h213209, value : 32'h3232}, //phyinit_io_write: 0x212209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h21020f, value : 32'h6}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Programming RxReplicaCtl04 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h21120f, value : 32'h6}, //phyinit_io_write: 0x21020f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h21220f, value : 32'h6}, //phyinit_io_write: 0x21120f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h21320f, value : 32'h6}, //phyinit_io_write: 0x21220f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h220005, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, DfiFreq=400MHz, Programming PipeCtl[AcInPipeEn]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h210008, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, DfiFreq=400MHz, Programming DBYTE0.LP5DfiDataEnLatency[LP5RLm13]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h211008, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, DfiFreq=400MHz, Programming DBYTE1.LP5DfiDataEnLatency[LP5RLm13]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h212008, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, DfiFreq=400MHz, Programming DBYTE2.LP5DfiDataEnLatency[LP5RLm13]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h213008, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, DfiFreq=400MHz, Programming DBYTE3.LP5DfiDataEnLatency[LP5RLm13]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h27006b, value : 32'h222}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, DfiFreq=400MHz, Programming DfiHandshakeDelays[PhyUpdReqDelay]=0x2 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h270066, value : 32'h20}, //phyinit_io_write: 0x27006b, 0x222
                          '{ step_type : REG_WRITE, reg_addr : 32'h2700eb, value : 32'h222}, //phyinit_io_write: 0x270066, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h2700e6, value : 32'h20}, //phyinit_io_write: 0x2700eb, 0x222
                          '{ step_type : REG_WRITE, reg_addr : 32'h270135, value : 32'h804}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACSMWckWriteFastTogglePulse::ACSMWckWriteFastToggleWidth to 0x19, ACSMWckWriteFastTogglePulse::ACSMWckWriteFastToggleDelay to 0x10
                          '{ step_type : REG_WRITE, reg_addr : 32'h270136, value : 32'h804}, //phyinit_io_write: 0x270135, 0x804
                          '{ step_type : REG_WRITE, reg_addr : 32'h270137, value : 32'h40c}, //phyinit_io_write: 0x270136, 0x804
                          '{ step_type : REG_WRITE, reg_addr : 32'h270138, value : 32'h1910}, //phyinit_io_write: 0x270137, 0x40c
                          '{ step_type : REG_WRITE, reg_addr : 32'h270139, value : 32'h808}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACSMWckReadFastTogglePulse::ACSMWckReadFastToggleWidth to 0x25, ACSMWckReadFastTogglePulse::ACSMWckReadFastToggleDelay to 0x14
                          '{ step_type : REG_WRITE, reg_addr : 32'h27013a, value : 32'h808}, //phyinit_io_write: 0x270139, 0x808
                          '{ step_type : REG_WRITE, reg_addr : 32'h27013b, value : 32'h410}, //phyinit_io_write: 0x27013a, 0x808
                          '{ step_type : REG_WRITE, reg_addr : 32'h27013c, value : 32'h2514}, //phyinit_io_write: 0x27013b, 0x410
                          '{ step_type : REG_WRITE, reg_addr : 32'h27013d, value : 32'h800}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACSMWckFreqFastTogglePulse::ACSMWckFreqFastToggleWidth to 0x11, ACSMWckFreqFastTogglePulse::ACSMWckFreqFastToggleDelay to 0xc
                          '{ step_type : REG_WRITE, reg_addr : 32'h27013e, value : 32'h800}, //phyinit_io_write: 0x27013d, 0x800
                          '{ step_type : REG_WRITE, reg_addr : 32'h27013f, value : 32'h408}, //phyinit_io_write: 0x27013e, 0x800
                          '{ step_type : REG_WRITE, reg_addr : 32'h270140, value : 32'h110c}, //phyinit_io_write: 0x27013f, 0x408
                          '{ step_type : REG_WRITE, reg_addr : 32'h27012c, value : 32'h81f}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACSMRxValPulse::ACSMRxValDelay to 0x1f, ACSMRxValPulse::ACSMRxValWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h27012d, value : 32'h81f}, //phyinit_io_write: 0x27012c, 0x81f
                          '{ step_type : REG_WRITE, reg_addr : 32'h270130, value : 32'h81f}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACSMRdcsPulse::ACSMRdcsDelay to 0x1f, ACSMRdcsPulse::ACSMRdcsWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h27012e, value : 32'h80f}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACSMTxEnPulse::ACSMTxEnDelay to 0xf, ACSMTxEnPulse::ACSMTxEnWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h27012f, value : 32'h80f}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming ACSMWrcsPulse::ACSMWrcsDelay to 0xf, ACSMWrcsPulse::ACSMWrcsWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h230008, value : 32'h0}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming AcPipeEn AC0 to 0. DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h231008, value : 32'h0}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, Programming AcPipeEn AC1 to 0. DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e0013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e1013, value : 32'h0}, //phyinit_io_write: 0x2e0013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e2013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e3013, value : 32'h0}, //phyinit_io_write: 0x2e2013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e4013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e5013, value : 32'h0}, //phyinit_io_write: 0x2e4013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e6013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e7013, value : 32'h0}, //phyinit_io_write: 0x2e6013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e0002, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Programming HMDBYTE RxDFECtrlDq to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e1002, value : 32'h0}, //phyinit_io_write: 0x2e0002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e2002, value : 32'h0}, //phyinit_io_write: 0x2e1002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e3002, value : 32'h0}, //phyinit_io_write: 0x2e2002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e4002, value : 32'h0}, //phyinit_io_write: 0x2e3002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e5002, value : 32'h0}, //phyinit_io_write: 0x2e4002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e6002, value : 32'h0}, //phyinit_io_write: 0x2e5002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e7002, value : 32'h0}, //phyinit_io_write: 0x2e6002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21010b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=2, Memclk=400MHz, freqThreshold=200MHz, NoRDQS=0 Programming InhibitTxRdPtrInit::DisableRxEnDlyLoad to 0x0, InhibitTxRdPtrInit::DisableTxDqDly to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21110b, value : 32'h0}, //phyinit_io_write: 0x21010b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21210b, value : 32'h0}, //phyinit_io_write: 0x21110b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21310b, value : 32'h0}, //phyinit_io_write: 0x21210b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h200063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC0 Instance0 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h201063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC1 Instance1 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h202063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC2 Instance2 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h203063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC3 Instance3 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h204063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC4 Instance4 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h205063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC5 Instance5 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h207063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC0 Instance7 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h208063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC1 Instance8 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h209063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC2 Instance9 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h20a063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC3 Instance10 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h20b063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC4 Instance11 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h20c063, value : 32'hd0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC5 Instance12 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h29080a, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Programming Seq0BGPR10 to HMTxLcdlSeed Full search value = 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h29080b, value : 32'hd0}, //phyinit_io_write: 0x29080a, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h290815, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Programming Seq0BGPR21 to ACHMTxLcdlSeed Full search value = 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h290816, value : 32'hd0}, //phyinit_io_write: 0x290815, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e0063, value : 32'hd0}, //phyinit_io_write: 0x290816, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e0064, value : 32'hd0}, //phyinit_io_write: 0x2e0063, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e0087, value : 32'hd0}, //phyinit_io_write: 0x2e0064, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e1063, value : 32'hd0}, //phyinit_io_write: 0x2e0087, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e1064, value : 32'hd0}, //phyinit_io_write: 0x2e1063, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e1087, value : 32'hd0}, //phyinit_io_write: 0x2e1064, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e2063, value : 32'hd0}, //phyinit_io_write: 0x2e1087, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e2064, value : 32'hd0}, //phyinit_io_write: 0x2e2063, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e2087, value : 32'hd0}, //phyinit_io_write: 0x2e2064, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e3063, value : 32'hd0}, //phyinit_io_write: 0x2e2087, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e3064, value : 32'hd0}, //phyinit_io_write: 0x2e3063, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e3087, value : 32'hd0}, //phyinit_io_write: 0x2e3064, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e4063, value : 32'hd0}, //phyinit_io_write: 0x2e3087, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e4064, value : 32'hd0}, //phyinit_io_write: 0x2e4063, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e4087, value : 32'hd0}, //phyinit_io_write: 0x2e4064, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e5063, value : 32'hd0}, //phyinit_io_write: 0x2e4087, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e5064, value : 32'hd0}, //phyinit_io_write: 0x2e5063, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e5087, value : 32'hd0}, //phyinit_io_write: 0x2e5064, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e6063, value : 32'hd0}, //phyinit_io_write: 0x2e5087, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e6064, value : 32'hd0}, //phyinit_io_write: 0x2e6063, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e6087, value : 32'hd0}, //phyinit_io_write: 0x2e6064, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e7063, value : 32'hd0}, //phyinit_io_write: 0x2e6087, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e7064, value : 32'hd0}, //phyinit_io_write: 0x2e7063, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e7087, value : 32'hd0}, //phyinit_io_write: 0x2e7064, 0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0080, value : 32'h7}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming UcclkHclkEnables to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e003c, value : 32'h80}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming RxDQSSeVrefDAC0 to 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e103c, value : 32'h80}, //phyinit_io_write: 0x2e003c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e203c, value : 32'h80}, //phyinit_io_write: 0x2e103c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e303c, value : 32'h80}, //phyinit_io_write: 0x2e203c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e403c, value : 32'h80}, //phyinit_io_write: 0x2e303c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e503c, value : 32'h80}, //phyinit_io_write: 0x2e403c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e603c, value : 32'h80}, //phyinit_io_write: 0x2e503c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e703c, value : 32'h80}, //phyinit_io_write: 0x2e603c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h290817, value : 32'h29}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 2 Seq0BGPR23 to 0x29, NumMemClk_tRFCab=164.0, NumMemClk_7p5ns=3.0, NumMemClk_tXSR=167.0
                          '{ step_type : REG_WRITE, reg_addr : 32'h290818, value : 32'h0}, //phyinit_io_write: 0x290817, 0x29
                          '{ step_type : REG_WRITE, reg_addr : 32'h290819, value : 32'h0}, //phyinit_io_write: 0x290818, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2300eb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 2 AC0 AcLcdlUpdInterval to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2310eb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 2 AC1 AcLcdlUpdInterval to 0x0
//[dwc_ddrphy_phyinit_programDfiMode] Skip DfiMode Programming: Keeping the reset value of 0x3
//End of dwc_ddrphy_phyinit_C_initPhyConfigPsLoop(), Pstate=2
                          '{ step_type : REG_WRITE, reg_addr : 32'h2300d9, value : 32'h40}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming CKXTxDly to 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2300d8, value : 32'h40}, //phyinit_io_write: 0x2300d9, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2301d8, value : 32'h40}, //phyinit_io_write: 0x2300d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2302d8, value : 32'h40}, //phyinit_io_write: 0x2301d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2303d8, value : 32'h40}, //phyinit_io_write: 0x2302d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2304d8, value : 32'h40}, //phyinit_io_write: 0x2303d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2305d8, value : 32'h40}, //phyinit_io_write: 0x2304d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2306d8, value : 32'h40}, //phyinit_io_write: 0x2305d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2308d8, value : 32'h40}, //phyinit_io_write: 0x2306d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2309d8, value : 32'h40}, //phyinit_io_write: 0x2308d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2310d9, value : 32'h40}, //phyinit_io_write: 0x2309d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2310d8, value : 32'h40}, //phyinit_io_write: 0x2310d9, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2311d8, value : 32'h40}, //phyinit_io_write: 0x2310d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2312d8, value : 32'h40}, //phyinit_io_write: 0x2311d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2313d8, value : 32'h40}, //phyinit_io_write: 0x2312d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2314d8, value : 32'h40}, //phyinit_io_write: 0x2313d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2315d8, value : 32'h40}, //phyinit_io_write: 0x2314d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2316d8, value : 32'h40}, //phyinit_io_write: 0x2315d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2318d8, value : 32'h40}, //phyinit_io_write: 0x2316d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h2319d8, value : 32'h40}, //phyinit_io_write: 0x2318d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h210000, value : 32'h6}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming HwtMRL to 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h211000, value : 32'h6}, //phyinit_io_write: 0x210000, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h212000, value : 32'h6}, //phyinit_io_write: 0x211000, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h213000, value : 32'h6}, //phyinit_io_write: 0x212000, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h27000d, value : 32'h6}, //phyinit_io_write: 0x213000, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h21002a, value : 32'h200}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming TxWckDlyTg0/Tg1 to 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h21002b, value : 32'h200}, //phyinit_io_write: 0x21002a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h21102a, value : 32'h200}, //phyinit_io_write: 0x21002b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h21102b, value : 32'h200}, //phyinit_io_write: 0x21102a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h21202a, value : 32'h200}, //phyinit_io_write: 0x21102b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h21202b, value : 32'h200}, //phyinit_io_write: 0x21202a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h21302a, value : 32'h200}, //phyinit_io_write: 0x21202b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h21302b, value : 32'h200}, //phyinit_io_write: 0x21302a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h210028, value : 32'h87}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming TxDqsDlyTg0/Tg1 to 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h210029, value : 32'h87}, //phyinit_io_write: 0x210028, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h211028, value : 32'h87}, //phyinit_io_write: 0x210029, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h211029, value : 32'h87}, //phyinit_io_write: 0x211028, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h212028, value : 32'h87}, //phyinit_io_write: 0x211029, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h212029, value : 32'h87}, //phyinit_io_write: 0x212028, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h213028, value : 32'h87}, //phyinit_io_write: 0x212029, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h213029, value : 32'h87}, //phyinit_io_write: 0x213028, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21007a, value : 32'h87}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming TxDqDlyTg0/Tg1 to 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21007b, value : 32'h87}, //phyinit_io_write: 0x21007a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21017a, value : 32'h87}, //phyinit_io_write: 0x21007b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21017b, value : 32'h87}, //phyinit_io_write: 0x21017a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21027a, value : 32'h87}, //phyinit_io_write: 0x21017b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21027b, value : 32'h87}, //phyinit_io_write: 0x21027a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21037a, value : 32'h87}, //phyinit_io_write: 0x21027b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21037b, value : 32'h87}, //phyinit_io_write: 0x21037a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21047a, value : 32'h87}, //phyinit_io_write: 0x21037b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21047b, value : 32'h87}, //phyinit_io_write: 0x21047a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21057a, value : 32'h87}, //phyinit_io_write: 0x21047b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21057b, value : 32'h87}, //phyinit_io_write: 0x21057a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21067a, value : 32'h87}, //phyinit_io_write: 0x21057b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21067b, value : 32'h87}, //phyinit_io_write: 0x21067a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21077a, value : 32'h87}, //phyinit_io_write: 0x21067b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21077b, value : 32'h87}, //phyinit_io_write: 0x21077a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21087a, value : 32'h87}, //phyinit_io_write: 0x21077b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21087b, value : 32'h87}, //phyinit_io_write: 0x21087a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21107a, value : 32'h87}, //phyinit_io_write: 0x21087b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21107b, value : 32'h87}, //phyinit_io_write: 0x21107a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21117a, value : 32'h87}, //phyinit_io_write: 0x21107b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21117b, value : 32'h87}, //phyinit_io_write: 0x21117a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21127a, value : 32'h87}, //phyinit_io_write: 0x21117b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21127b, value : 32'h87}, //phyinit_io_write: 0x21127a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21137a, value : 32'h87}, //phyinit_io_write: 0x21127b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21137b, value : 32'h87}, //phyinit_io_write: 0x21137a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21147a, value : 32'h87}, //phyinit_io_write: 0x21137b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21147b, value : 32'h87}, //phyinit_io_write: 0x21147a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21157a, value : 32'h87}, //phyinit_io_write: 0x21147b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21157b, value : 32'h87}, //phyinit_io_write: 0x21157a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21167a, value : 32'h87}, //phyinit_io_write: 0x21157b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21167b, value : 32'h87}, //phyinit_io_write: 0x21167a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21177a, value : 32'h87}, //phyinit_io_write: 0x21167b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21177b, value : 32'h87}, //phyinit_io_write: 0x21177a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21187a, value : 32'h87}, //phyinit_io_write: 0x21177b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21187b, value : 32'h87}, //phyinit_io_write: 0x21187a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21207a, value : 32'h87}, //phyinit_io_write: 0x21187b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21207b, value : 32'h87}, //phyinit_io_write: 0x21207a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21217a, value : 32'h87}, //phyinit_io_write: 0x21207b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21217b, value : 32'h87}, //phyinit_io_write: 0x21217a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21227a, value : 32'h87}, //phyinit_io_write: 0x21217b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21227b, value : 32'h87}, //phyinit_io_write: 0x21227a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21237a, value : 32'h87}, //phyinit_io_write: 0x21227b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21237b, value : 32'h87}, //phyinit_io_write: 0x21237a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21247a, value : 32'h87}, //phyinit_io_write: 0x21237b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21247b, value : 32'h87}, //phyinit_io_write: 0x21247a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21257a, value : 32'h87}, //phyinit_io_write: 0x21247b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21257b, value : 32'h87}, //phyinit_io_write: 0x21257a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21267a, value : 32'h87}, //phyinit_io_write: 0x21257b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21267b, value : 32'h87}, //phyinit_io_write: 0x21267a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21277a, value : 32'h87}, //phyinit_io_write: 0x21267b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21277b, value : 32'h87}, //phyinit_io_write: 0x21277a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21287a, value : 32'h87}, //phyinit_io_write: 0x21277b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21287b, value : 32'h87}, //phyinit_io_write: 0x21287a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21307a, value : 32'h87}, //phyinit_io_write: 0x21287b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21307b, value : 32'h87}, //phyinit_io_write: 0x21307a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21317a, value : 32'h87}, //phyinit_io_write: 0x21307b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21317b, value : 32'h87}, //phyinit_io_write: 0x21317a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21327a, value : 32'h87}, //phyinit_io_write: 0x21317b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21327b, value : 32'h87}, //phyinit_io_write: 0x21327a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21337a, value : 32'h87}, //phyinit_io_write: 0x21327b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21337b, value : 32'h87}, //phyinit_io_write: 0x21337a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21347a, value : 32'h87}, //phyinit_io_write: 0x21337b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21347b, value : 32'h87}, //phyinit_io_write: 0x21347a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21357a, value : 32'h87}, //phyinit_io_write: 0x21347b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21357b, value : 32'h87}, //phyinit_io_write: 0x21357a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21367a, value : 32'h87}, //phyinit_io_write: 0x21357b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21367b, value : 32'h87}, //phyinit_io_write: 0x21367a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21377a, value : 32'h87}, //phyinit_io_write: 0x21367b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21377b, value : 32'h87}, //phyinit_io_write: 0x21377a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21387a, value : 32'h87}, //phyinit_io_write: 0x21377b, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h21387b, value : 32'h87}, //phyinit_io_write: 0x21387a, 0x87
                          '{ step_type : REG_WRITE, reg_addr : 32'h210078, value : 32'h2ec}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming RxDigStrbDlyTg0/Tg1 to 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210079, value : 32'h2ec}, //phyinit_io_write: 0x210078, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210178, value : 32'h2ec}, //phyinit_io_write: 0x210079, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210179, value : 32'h2ec}, //phyinit_io_write: 0x210178, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210278, value : 32'h2ec}, //phyinit_io_write: 0x210179, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210279, value : 32'h2ec}, //phyinit_io_write: 0x210278, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210378, value : 32'h2ec}, //phyinit_io_write: 0x210279, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210379, value : 32'h2ec}, //phyinit_io_write: 0x210378, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210478, value : 32'h2ec}, //phyinit_io_write: 0x210379, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210479, value : 32'h2ec}, //phyinit_io_write: 0x210478, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210578, value : 32'h2ec}, //phyinit_io_write: 0x210479, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210579, value : 32'h2ec}, //phyinit_io_write: 0x210578, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210678, value : 32'h2ec}, //phyinit_io_write: 0x210579, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210679, value : 32'h2ec}, //phyinit_io_write: 0x210678, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210778, value : 32'h2ec}, //phyinit_io_write: 0x210679, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210779, value : 32'h2ec}, //phyinit_io_write: 0x210778, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210878, value : 32'h2ec}, //phyinit_io_write: 0x210779, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210879, value : 32'h2ec}, //phyinit_io_write: 0x210878, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211078, value : 32'h2ec}, //phyinit_io_write: 0x210879, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211079, value : 32'h2ec}, //phyinit_io_write: 0x211078, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211178, value : 32'h2ec}, //phyinit_io_write: 0x211079, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211179, value : 32'h2ec}, //phyinit_io_write: 0x211178, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211278, value : 32'h2ec}, //phyinit_io_write: 0x211179, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211279, value : 32'h2ec}, //phyinit_io_write: 0x211278, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211378, value : 32'h2ec}, //phyinit_io_write: 0x211279, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211379, value : 32'h2ec}, //phyinit_io_write: 0x211378, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211478, value : 32'h2ec}, //phyinit_io_write: 0x211379, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211479, value : 32'h2ec}, //phyinit_io_write: 0x211478, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211578, value : 32'h2ec}, //phyinit_io_write: 0x211479, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211579, value : 32'h2ec}, //phyinit_io_write: 0x211578, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211678, value : 32'h2ec}, //phyinit_io_write: 0x211579, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211679, value : 32'h2ec}, //phyinit_io_write: 0x211678, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211778, value : 32'h2ec}, //phyinit_io_write: 0x211679, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211779, value : 32'h2ec}, //phyinit_io_write: 0x211778, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211878, value : 32'h2ec}, //phyinit_io_write: 0x211779, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h211879, value : 32'h2ec}, //phyinit_io_write: 0x211878, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212078, value : 32'h2ec}, //phyinit_io_write: 0x211879, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212079, value : 32'h2ec}, //phyinit_io_write: 0x212078, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212178, value : 32'h2ec}, //phyinit_io_write: 0x212079, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212179, value : 32'h2ec}, //phyinit_io_write: 0x212178, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212278, value : 32'h2ec}, //phyinit_io_write: 0x212179, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212279, value : 32'h2ec}, //phyinit_io_write: 0x212278, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212378, value : 32'h2ec}, //phyinit_io_write: 0x212279, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212379, value : 32'h2ec}, //phyinit_io_write: 0x212378, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212478, value : 32'h2ec}, //phyinit_io_write: 0x212379, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212479, value : 32'h2ec}, //phyinit_io_write: 0x212478, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212578, value : 32'h2ec}, //phyinit_io_write: 0x212479, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212579, value : 32'h2ec}, //phyinit_io_write: 0x212578, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212678, value : 32'h2ec}, //phyinit_io_write: 0x212579, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212679, value : 32'h2ec}, //phyinit_io_write: 0x212678, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212778, value : 32'h2ec}, //phyinit_io_write: 0x212679, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212779, value : 32'h2ec}, //phyinit_io_write: 0x212778, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212878, value : 32'h2ec}, //phyinit_io_write: 0x212779, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h212879, value : 32'h2ec}, //phyinit_io_write: 0x212878, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213078, value : 32'h2ec}, //phyinit_io_write: 0x212879, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213079, value : 32'h2ec}, //phyinit_io_write: 0x213078, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213178, value : 32'h2ec}, //phyinit_io_write: 0x213079, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213179, value : 32'h2ec}, //phyinit_io_write: 0x213178, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213278, value : 32'h2ec}, //phyinit_io_write: 0x213179, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213279, value : 32'h2ec}, //phyinit_io_write: 0x213278, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213378, value : 32'h2ec}, //phyinit_io_write: 0x213279, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213379, value : 32'h2ec}, //phyinit_io_write: 0x213378, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213478, value : 32'h2ec}, //phyinit_io_write: 0x213379, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213479, value : 32'h2ec}, //phyinit_io_write: 0x213478, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213578, value : 32'h2ec}, //phyinit_io_write: 0x213479, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213579, value : 32'h2ec}, //phyinit_io_write: 0x213578, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213678, value : 32'h2ec}, //phyinit_io_write: 0x213579, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213679, value : 32'h2ec}, //phyinit_io_write: 0x213678, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213778, value : 32'h2ec}, //phyinit_io_write: 0x213679, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213779, value : 32'h2ec}, //phyinit_io_write: 0x213778, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213878, value : 32'h2ec}, //phyinit_io_write: 0x213779, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h213879, value : 32'h2ec}, //phyinit_io_write: 0x213878, 0x2ec
                          '{ step_type : REG_WRITE, reg_addr : 32'h210020, value : 32'h24c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming RxEnDlyTg0/Tg1 to 0x24c
                          '{ step_type : REG_WRITE, reg_addr : 32'h210021, value : 32'h24c}, //phyinit_io_write: 0x210020, 0x24c
                          '{ step_type : REG_WRITE, reg_addr : 32'h211020, value : 32'h24c}, //phyinit_io_write: 0x210021, 0x24c
                          '{ step_type : REG_WRITE, reg_addr : 32'h211021, value : 32'h24c}, //phyinit_io_write: 0x211020, 0x24c
                          '{ step_type : REG_WRITE, reg_addr : 32'h212020, value : 32'h24c}, //phyinit_io_write: 0x211021, 0x24c
                          '{ step_type : REG_WRITE, reg_addr : 32'h212021, value : 32'h24c}, //phyinit_io_write: 0x212020, 0x24c
                          '{ step_type : REG_WRITE, reg_addr : 32'h213020, value : 32'h24c}, //phyinit_io_write: 0x212021, 0x24c
                          '{ step_type : REG_WRITE, reg_addr : 32'h213021, value : 32'h24c}, //phyinit_io_write: 0x213020, 0x24c
                          '{ step_type : REG_WRITE, reg_addr : 32'h210010, value : 32'h1a5}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming RxClkT2UIDlyTg0/Tg1 and RxClkC2UIDlyTg0/Tg1 to 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210011, value : 32'h1a5}, //phyinit_io_write: 0x210010, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210012, value : 32'h1a5}, //phyinit_io_write: 0x210011, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210013, value : 32'h1a5}, //phyinit_io_write: 0x210012, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210110, value : 32'h1a5}, //phyinit_io_write: 0x210013, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210111, value : 32'h1a5}, //phyinit_io_write: 0x210110, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210112, value : 32'h1a5}, //phyinit_io_write: 0x210111, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210113, value : 32'h1a5}, //phyinit_io_write: 0x210112, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210210, value : 32'h1a5}, //phyinit_io_write: 0x210113, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210211, value : 32'h1a5}, //phyinit_io_write: 0x210210, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210212, value : 32'h1a5}, //phyinit_io_write: 0x210211, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210213, value : 32'h1a5}, //phyinit_io_write: 0x210212, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210310, value : 32'h1a5}, //phyinit_io_write: 0x210213, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210311, value : 32'h1a5}, //phyinit_io_write: 0x210310, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210312, value : 32'h1a5}, //phyinit_io_write: 0x210311, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210313, value : 32'h1a5}, //phyinit_io_write: 0x210312, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210410, value : 32'h1a5}, //phyinit_io_write: 0x210313, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210411, value : 32'h1a5}, //phyinit_io_write: 0x210410, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210412, value : 32'h1a5}, //phyinit_io_write: 0x210411, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210413, value : 32'h1a5}, //phyinit_io_write: 0x210412, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210510, value : 32'h1a5}, //phyinit_io_write: 0x210413, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210511, value : 32'h1a5}, //phyinit_io_write: 0x210510, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210512, value : 32'h1a5}, //phyinit_io_write: 0x210511, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210513, value : 32'h1a5}, //phyinit_io_write: 0x210512, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210610, value : 32'h1a5}, //phyinit_io_write: 0x210513, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210611, value : 32'h1a5}, //phyinit_io_write: 0x210610, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210612, value : 32'h1a5}, //phyinit_io_write: 0x210611, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210613, value : 32'h1a5}, //phyinit_io_write: 0x210612, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210710, value : 32'h1a5}, //phyinit_io_write: 0x210613, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210711, value : 32'h1a5}, //phyinit_io_write: 0x210710, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210712, value : 32'h1a5}, //phyinit_io_write: 0x210711, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210713, value : 32'h1a5}, //phyinit_io_write: 0x210712, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210810, value : 32'h1a5}, //phyinit_io_write: 0x210713, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210811, value : 32'h1a5}, //phyinit_io_write: 0x210810, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210812, value : 32'h1a5}, //phyinit_io_write: 0x210811, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h210813, value : 32'h1a5}, //phyinit_io_write: 0x210812, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211010, value : 32'h1a5}, //phyinit_io_write: 0x210813, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211011, value : 32'h1a5}, //phyinit_io_write: 0x211010, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211012, value : 32'h1a5}, //phyinit_io_write: 0x211011, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211013, value : 32'h1a5}, //phyinit_io_write: 0x211012, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211110, value : 32'h1a5}, //phyinit_io_write: 0x211013, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211111, value : 32'h1a5}, //phyinit_io_write: 0x211110, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211112, value : 32'h1a5}, //phyinit_io_write: 0x211111, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211113, value : 32'h1a5}, //phyinit_io_write: 0x211112, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211210, value : 32'h1a5}, //phyinit_io_write: 0x211113, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211211, value : 32'h1a5}, //phyinit_io_write: 0x211210, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211212, value : 32'h1a5}, //phyinit_io_write: 0x211211, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211213, value : 32'h1a5}, //phyinit_io_write: 0x211212, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211310, value : 32'h1a5}, //phyinit_io_write: 0x211213, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211311, value : 32'h1a5}, //phyinit_io_write: 0x211310, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211312, value : 32'h1a5}, //phyinit_io_write: 0x211311, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211313, value : 32'h1a5}, //phyinit_io_write: 0x211312, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211410, value : 32'h1a5}, //phyinit_io_write: 0x211313, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211411, value : 32'h1a5}, //phyinit_io_write: 0x211410, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211412, value : 32'h1a5}, //phyinit_io_write: 0x211411, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211413, value : 32'h1a5}, //phyinit_io_write: 0x211412, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211510, value : 32'h1a5}, //phyinit_io_write: 0x211413, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211511, value : 32'h1a5}, //phyinit_io_write: 0x211510, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211512, value : 32'h1a5}, //phyinit_io_write: 0x211511, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211513, value : 32'h1a5}, //phyinit_io_write: 0x211512, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211610, value : 32'h1a5}, //phyinit_io_write: 0x211513, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211611, value : 32'h1a5}, //phyinit_io_write: 0x211610, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211612, value : 32'h1a5}, //phyinit_io_write: 0x211611, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211613, value : 32'h1a5}, //phyinit_io_write: 0x211612, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211710, value : 32'h1a5}, //phyinit_io_write: 0x211613, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211711, value : 32'h1a5}, //phyinit_io_write: 0x211710, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211712, value : 32'h1a5}, //phyinit_io_write: 0x211711, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211713, value : 32'h1a5}, //phyinit_io_write: 0x211712, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211810, value : 32'h1a5}, //phyinit_io_write: 0x211713, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211811, value : 32'h1a5}, //phyinit_io_write: 0x211810, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211812, value : 32'h1a5}, //phyinit_io_write: 0x211811, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h211813, value : 32'h1a5}, //phyinit_io_write: 0x211812, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212010, value : 32'h1a5}, //phyinit_io_write: 0x211813, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212011, value : 32'h1a5}, //phyinit_io_write: 0x212010, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212012, value : 32'h1a5}, //phyinit_io_write: 0x212011, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212013, value : 32'h1a5}, //phyinit_io_write: 0x212012, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212110, value : 32'h1a5}, //phyinit_io_write: 0x212013, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212111, value : 32'h1a5}, //phyinit_io_write: 0x212110, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212112, value : 32'h1a5}, //phyinit_io_write: 0x212111, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212113, value : 32'h1a5}, //phyinit_io_write: 0x212112, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212210, value : 32'h1a5}, //phyinit_io_write: 0x212113, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212211, value : 32'h1a5}, //phyinit_io_write: 0x212210, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212212, value : 32'h1a5}, //phyinit_io_write: 0x212211, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212213, value : 32'h1a5}, //phyinit_io_write: 0x212212, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212310, value : 32'h1a5}, //phyinit_io_write: 0x212213, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212311, value : 32'h1a5}, //phyinit_io_write: 0x212310, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212312, value : 32'h1a5}, //phyinit_io_write: 0x212311, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212313, value : 32'h1a5}, //phyinit_io_write: 0x212312, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212410, value : 32'h1a5}, //phyinit_io_write: 0x212313, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212411, value : 32'h1a5}, //phyinit_io_write: 0x212410, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212412, value : 32'h1a5}, //phyinit_io_write: 0x212411, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212413, value : 32'h1a5}, //phyinit_io_write: 0x212412, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212510, value : 32'h1a5}, //phyinit_io_write: 0x212413, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212511, value : 32'h1a5}, //phyinit_io_write: 0x212510, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212512, value : 32'h1a5}, //phyinit_io_write: 0x212511, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212513, value : 32'h1a5}, //phyinit_io_write: 0x212512, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212610, value : 32'h1a5}, //phyinit_io_write: 0x212513, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212611, value : 32'h1a5}, //phyinit_io_write: 0x212610, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212612, value : 32'h1a5}, //phyinit_io_write: 0x212611, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212613, value : 32'h1a5}, //phyinit_io_write: 0x212612, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212710, value : 32'h1a5}, //phyinit_io_write: 0x212613, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212711, value : 32'h1a5}, //phyinit_io_write: 0x212710, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212712, value : 32'h1a5}, //phyinit_io_write: 0x212711, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212713, value : 32'h1a5}, //phyinit_io_write: 0x212712, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212810, value : 32'h1a5}, //phyinit_io_write: 0x212713, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212811, value : 32'h1a5}, //phyinit_io_write: 0x212810, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212812, value : 32'h1a5}, //phyinit_io_write: 0x212811, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h212813, value : 32'h1a5}, //phyinit_io_write: 0x212812, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213010, value : 32'h1a5}, //phyinit_io_write: 0x212813, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213011, value : 32'h1a5}, //phyinit_io_write: 0x213010, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213012, value : 32'h1a5}, //phyinit_io_write: 0x213011, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213013, value : 32'h1a5}, //phyinit_io_write: 0x213012, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213110, value : 32'h1a5}, //phyinit_io_write: 0x213013, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213111, value : 32'h1a5}, //phyinit_io_write: 0x213110, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213112, value : 32'h1a5}, //phyinit_io_write: 0x213111, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213113, value : 32'h1a5}, //phyinit_io_write: 0x213112, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213210, value : 32'h1a5}, //phyinit_io_write: 0x213113, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213211, value : 32'h1a5}, //phyinit_io_write: 0x213210, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213212, value : 32'h1a5}, //phyinit_io_write: 0x213211, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213213, value : 32'h1a5}, //phyinit_io_write: 0x213212, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213310, value : 32'h1a5}, //phyinit_io_write: 0x213213, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213311, value : 32'h1a5}, //phyinit_io_write: 0x213310, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213312, value : 32'h1a5}, //phyinit_io_write: 0x213311, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213313, value : 32'h1a5}, //phyinit_io_write: 0x213312, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213410, value : 32'h1a5}, //phyinit_io_write: 0x213313, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213411, value : 32'h1a5}, //phyinit_io_write: 0x213410, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213412, value : 32'h1a5}, //phyinit_io_write: 0x213411, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213413, value : 32'h1a5}, //phyinit_io_write: 0x213412, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213510, value : 32'h1a5}, //phyinit_io_write: 0x213413, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213511, value : 32'h1a5}, //phyinit_io_write: 0x213510, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213512, value : 32'h1a5}, //phyinit_io_write: 0x213511, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213513, value : 32'h1a5}, //phyinit_io_write: 0x213512, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213610, value : 32'h1a5}, //phyinit_io_write: 0x213513, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213611, value : 32'h1a5}, //phyinit_io_write: 0x213610, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213612, value : 32'h1a5}, //phyinit_io_write: 0x213611, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213613, value : 32'h1a5}, //phyinit_io_write: 0x213612, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213710, value : 32'h1a5}, //phyinit_io_write: 0x213613, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213711, value : 32'h1a5}, //phyinit_io_write: 0x213710, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213712, value : 32'h1a5}, //phyinit_io_write: 0x213711, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213713, value : 32'h1a5}, //phyinit_io_write: 0x213712, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213810, value : 32'h1a5}, //phyinit_io_write: 0x213713, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213811, value : 32'h1a5}, //phyinit_io_write: 0x213810, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213812, value : 32'h1a5}, //phyinit_io_write: 0x213811, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h213813, value : 32'h1a5}, //phyinit_io_write: 0x213812, 0x1a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h21000c, value : 32'h67}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming PptWck2DqoCntInvTrn1 to 0xcd
                          '{ step_type : REG_WRITE, reg_addr : 32'h21000d, value : 32'h67}, //phyinit_io_write: 0x21000c, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h210014, value : 32'hcd}, //phyinit_io_write: 0x21000d, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h210015, value : 32'hcd}, //phyinit_io_write: 0x210014, 0xcd
                          '{ step_type : REG_WRITE, reg_addr : 32'h21100c, value : 32'h67}, //phyinit_io_write: 0x210015, 0xcd
                          '{ step_type : REG_WRITE, reg_addr : 32'h21100d, value : 32'h67}, //phyinit_io_write: 0x21100c, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h211014, value : 32'hcd}, //phyinit_io_write: 0x21100d, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h211015, value : 32'hcd}, //phyinit_io_write: 0x211014, 0xcd
                          '{ step_type : REG_WRITE, reg_addr : 32'h21200c, value : 32'h67}, //phyinit_io_write: 0x211015, 0xcd
                          '{ step_type : REG_WRITE, reg_addr : 32'h21200d, value : 32'h67}, //phyinit_io_write: 0x21200c, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h212014, value : 32'hcd}, //phyinit_io_write: 0x21200d, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h212015, value : 32'hcd}, //phyinit_io_write: 0x212014, 0xcd
                          '{ step_type : REG_WRITE, reg_addr : 32'h21300c, value : 32'h67}, //phyinit_io_write: 0x212015, 0xcd
                          '{ step_type : REG_WRITE, reg_addr : 32'h21300d, value : 32'h67}, //phyinit_io_write: 0x21300c, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h213014, value : 32'hcd}, //phyinit_io_write: 0x21300d, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h213015, value : 32'hcd}, //phyinit_io_write: 0x213014, 0xcd
                          '{ step_type : REG_WRITE, reg_addr : 32'h70077, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming HwtCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h220071, value : 32'h55}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming HMRxReplicaLcdlSeed HMRxSeed to 0xc5 HMRxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h200063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC0 Instance0 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h201063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC1 Instance1 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h202063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC2 Instance2 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h203063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC3 Instance3 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h204063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC4 Instance4 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h205063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX0 HMAC5 Instance5 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h207063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC0 Instance7 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h208063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC1 Instance8 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h209063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC2 Instance9 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h20a063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC3 Instance10 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h20b063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC4 Instance11 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h20c063, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=2, Memclk=400MHz, Programming ACX1 HMAC5 Instance12 HMTxLcdlSeed HMTxSeed to 0xc5 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e0063, value : 32'hc5}, //phyinit_io_write: 0x20c063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e0064, value : 32'hc5}, //phyinit_io_write: 0x2e0063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e0087, value : 32'hc5}, //phyinit_io_write: 0x2e0064, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e1063, value : 32'hc5}, //phyinit_io_write: 0x2e0087, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e1064, value : 32'hc5}, //phyinit_io_write: 0x2e1063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e1087, value : 32'hc5}, //phyinit_io_write: 0x2e1064, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e2063, value : 32'hc5}, //phyinit_io_write: 0x2e1087, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e2064, value : 32'hc5}, //phyinit_io_write: 0x2e2063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e2087, value : 32'hc5}, //phyinit_io_write: 0x2e2064, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e3063, value : 32'hc5}, //phyinit_io_write: 0x2e2087, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e3064, value : 32'hc5}, //phyinit_io_write: 0x2e3063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e3087, value : 32'hc5}, //phyinit_io_write: 0x2e3064, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e4063, value : 32'hc5}, //phyinit_io_write: 0x2e3087, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e4064, value : 32'hc5}, //phyinit_io_write: 0x2e4063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e4087, value : 32'hc5}, //phyinit_io_write: 0x2e4064, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e5063, value : 32'hc5}, //phyinit_io_write: 0x2e4087, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e5064, value : 32'hc5}, //phyinit_io_write: 0x2e5063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e5087, value : 32'hc5}, //phyinit_io_write: 0x2e5064, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e6063, value : 32'hc5}, //phyinit_io_write: 0x2e5087, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e6064, value : 32'hc5}, //phyinit_io_write: 0x2e6063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e6087, value : 32'hc5}, //phyinit_io_write: 0x2e6064, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e7063, value : 32'hc5}, //phyinit_io_write: 0x2e6087, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e7064, value : 32'hc5}, //phyinit_io_write: 0x2e7063, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e7087, value : 32'hc5}, //phyinit_io_write: 0x2e7064, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h29080a, value : 32'h2c5}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=2 Programming Seq0bGPR10 to mission mode HMTxLcdlSeed value 0x2c5
                          '{ step_type : REG_WRITE, reg_addr : 32'h29080b, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=2 Programming Seq0bGPR11 to mission mode HMTxLcdlSeed value 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h290815, value : 32'h2c5}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=2 Programming Seq0bGPR21 to mission mode HMTxLcdlSeed value 0x2c5
                          '{ step_type : REG_WRITE, reg_addr : 32'h290816, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=2 Programming Seq0bGPR22 to mission mode HMTxLcdlSeed value 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h21015f, value : 32'hc5}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=2, Memclk=400MHz, Programming RDqRDqsCntrl to 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h21115f, value : 32'hc5}, //phyinit_io_write: 0x21015f, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h21215f, value : 32'hc5}, //phyinit_io_write: 0x21115f, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h21315f, value : 32'hc5}, //phyinit_io_write: 0x21215f, 0xc5
                          '{ step_type : REG_WRITE, reg_addr : 32'h260009, value : 32'h10}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Memclk=400MHz, Programming CPllDacValIn to 0x10
                          '{ step_type : REG_WRITE, reg_addr : 32'h2102a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE0.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2102a1, value : 32'ha}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE0.RxReplicaPathPhase1 to 0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h2102a2, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE0.RxReplicaPathPhase2 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h2102a3, value : 32'hda}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE0.RxReplicaPathPhase3 to 0xda
                          '{ step_type : REG_WRITE, reg_addr : 32'h2102a4, value : 32'h142}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE0.RxReplicaPathPhase4 to 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h2112a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE1.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2112a1, value : 32'ha}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE1.RxReplicaPathPhase1 to 0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h2112a2, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE1.RxReplicaPathPhase2 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h2112a3, value : 32'hda}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE1.RxReplicaPathPhase3 to 0xda
                          '{ step_type : REG_WRITE, reg_addr : 32'h2112a4, value : 32'h142}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE1.RxReplicaPathPhase4 to 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h2122a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE2.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2122a1, value : 32'ha}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE2.RxReplicaPathPhase1 to 0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h2122a2, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE2.RxReplicaPathPhase2 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h2122a3, value : 32'hda}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE2.RxReplicaPathPhase3 to 0xda
                          '{ step_type : REG_WRITE, reg_addr : 32'h2122a4, value : 32'h142}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE2.RxReplicaPathPhase4 to 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h2132a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE3.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2132a1, value : 32'ha}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE3.RxReplicaPathPhase1 to 0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h2132a2, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE3.RxReplicaPathPhase2 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h2132a3, value : 32'hda}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE3.RxReplicaPathPhase3 to 0xda
                          '{ step_type : REG_WRITE, reg_addr : 32'h2132a4, value : 32'h142}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE3.RxReplicaPathPhase4 to 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h2102ad, value : 32'h2}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE0.RxReplicaCtl01::RxReplicaSelPathPhase to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h2112ad, value : 32'h2}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE1.RxReplicaCtl01::RxReplicaSelPathPhase to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h2122ad, value : 32'h2}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE2.RxReplicaCtl01::RxReplicaSelPathPhase to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h2132ad, value : 32'h2}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE3.RxReplicaCtl01::RxReplicaSelPathPhase to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h2102af, value : 32'h46}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE0.RxReplicaCtl03 to 0x46
                          '{ step_type : REG_WRITE, reg_addr : 32'h2112af, value : 32'h46}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE1.RxReplicaCtl03 to 0x46
                          '{ step_type : REG_WRITE, reg_addr : 32'h2122af, value : 32'h46}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE2.RxReplicaCtl03 to 0x46
                          '{ step_type : REG_WRITE, reg_addr : 32'h2132af, value : 32'h46}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming DBYTE3.RxReplicaCtl03 to 0x46
                          '{ step_type : REG_WRITE, reg_addr : 32'h290807, value : 32'h9701}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming Seq0BGPR7 to save ZQCalCodeOvrValPU=0x12e and ZQCalCodeOvrEnPU=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h290808, value : 32'hb681}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=2, Programming Seq0BGPR8 to save ZQCalCodeOvrValPD=0x16d and ZQCalCodeOvrEnPD=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
//[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] End of dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop(), PState=2
// [dwc_ddrphy_phyinit_userCustom_E_setDfiClk] Start of dwc_ddrphy_phyinit_userCustom_E_setDfiClk()
// [dwc_ddrphy_phyinit_userCustom_E_setDfiClk] End of dwc_ddrphy_phyinit_userCustom_E_setDfiClk()
// [dwc_ddrphy_phyinit_F_loadDMEM1D] Start of dwc_ddrphy_phyinit_F_loadDMEM (pstate=2, Train2D=0)
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0088, value : 32'h1}, //[dwc_ddrphy_phyinit_F_loadDMEM] Program csr StartDccmClear to 1 to clear DCCM.
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 8300},
//Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 8300 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0088, value : 32'h0}, //[dwc_ddrphy_phyinit_F_loadDMEM] Program csr StartDccmClear to 0 after DCCM clear is done.
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}, //Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 40 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'h58000, value : 32'h600}, // [dwc_ddrphy_phyinit_WriteOutMem] STARTING. offset 0x58000 size 0x6000, sparse_write=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h58001, value : 32'hc800002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58002, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58004, value : 32'hff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58005, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58009, value : 32'h310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5800f, value : 32'h10000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58010, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58016, value : 32'h50500000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58017, value : 32'h55555050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58018, value : 32'he0e5555},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58019, value : 32'h54540e0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801a, value : 32'h44445454},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801b, value : 32'h50504444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801c, value : 32'h5050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801d, value : 32'h50500000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801e, value : 32'h50505050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801f, value : 32'h5050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58020, value : 32'hac840000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58021, value : 32'hac84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58023, value : 32'h2020000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58024, value : 32'h202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5802a, value : 32'h4040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5802b, value : 32'h404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58032, value : 32'h60600000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58033, value : 32'h6060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58048, value : 32'h23000001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58049, value : 32'h1f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58054, value : 32'h5c0032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58055, value : 32'he000b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58056, value : 32'h164013a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58057, value : 32'h1e801be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58062, value : 32'h6400c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58103, value : 32'h50b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58104, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58108, value : 32'h8080808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58110, value : 32'hef0f4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811b, value : 32'h4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811d, value : 32'h40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811e, value : 32'h180f0e0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811f, value : 32'h4746451e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58120, value : 32'h4a4948},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58121, value : 32'h1000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58125, value : 32'h40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58126, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58129, value : 32'hffffffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5812e, value : 32'h2f059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5812f, value : 32'hffb50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58130, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58131, value : 32'h1f0b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58132, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58133, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58134, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58135, value : 32'hf0b00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58136, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58137, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58138, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58139, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813a, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813b, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813c, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813d, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813e, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813f, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58140, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58141, value : 32'hff740182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58142, value : 32'h800001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58143, value : 32'h1ffbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58144, value : 32'hf0be0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58145, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58146, value : 32'h1f0a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58147, value : 32'hf0a20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58148, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58149, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814a, value : 32'h40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814b, value : 32'h308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814c, value : 32'h560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814e, value : 32'h80000dbc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814f, value : 32'h309},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58150, value : 32'h561},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58151, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58152, value : 32'h80000dcd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58153, value : 32'he0305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58154, value : 32'he0205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58155, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58156, value : 32'h80000dde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58157, value : 32'he0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58158, value : 32'he0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58159, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815a, value : 32'h80000e44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815b, value : 32'he0301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815c, value : 32'he0201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815d, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815e, value : 32'h80000e57},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815f, value : 32'he0302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58160, value : 32'he0202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58161, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58162, value : 32'h80000e6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58163, value : 32'he0303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58164, value : 32'he0203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58165, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58166, value : 32'h80000e7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58167, value : 32'he0304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58168, value : 32'he0204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58169, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816a, value : 32'h80000e90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816b, value : 32'h1ff01ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816c, value : 32'he0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816e, value : 32'h63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816f, value : 32'h64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58170, value : 32'h660},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58172, value : 32'h80000d8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58173, value : 32'h661},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58174, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58175, value : 32'h80000dad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58176, value : 32'he00f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58177, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58178, value : 32'h80000def},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58179, value : 32'he00f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817a, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817b, value : 32'h80000e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817c, value : 32'he00f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817d, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817e, value : 32'h80000e11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817f, value : 32'he00f3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58180, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58181, value : 32'h80000e22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58182, value : 32'he00f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58183, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58184, value : 32'h80000e33},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58185, value : 32'he00f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58186, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58187, value : 32'h80000d9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58188, value : 32'h2011210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58189, value : 32'h1c0a1403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818a, value : 32'hb112e29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818b, value : 32'h1916150d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818c, value : 32'h180f0e0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818d, value : 32'h453a131e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818e, value : 32'h49484746},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818f, value : 32'h2006e4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58190, value : 32'h100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58191, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58192, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58194, value : 32'h2150001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58195, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58196, value : 32'h1010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58197, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58198, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58199, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819a, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819b, value : 32'h6400002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819c, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819d, value : 32'h30215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819e, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819f, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a0, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a1, value : 32'h10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a2, value : 32'habe0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a3, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a4, value : 32'h50320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a5, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c5, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c6, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c7, value : 32'h43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c8, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c9, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ca, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cb, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cc, value : 32'h42b0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cd, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ce, value : 32'h200c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cf, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d0, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d1, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d2, value : 32'h10003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d3, value : 32'h8550002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d4, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d5, value : 32'h40158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d6, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d7, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d8, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d9, value : 32'h10005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581da, value : 32'hc800002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581db, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581dc, value : 32'h601d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581dd, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581de, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581df, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e0, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e1, value : 32'h10ab0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e2, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e3, value : 32'h80258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e4, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e5, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e6, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e7, value : 32'h20009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e8, value : 32'h157c0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e9, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ea, value : 32'ha02ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581eb, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ec, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ed, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ee, value : 32'h2000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ef, value : 32'h19000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f0, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f1, value : 32'hc03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f2, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f3, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f4, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f5, value : 32'h3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f6, value : 32'h21550006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f7, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f8, value : 32'he04b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f9, value : 32'h70003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fa, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fb, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fc, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fd, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fe, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ff, value : 32'h2150004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58200, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58201, value : 32'h4010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58202, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58203, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58204, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58205, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58206, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58207, value : 32'h80006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58208, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58209, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820a, value : 32'h6400006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820b, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820c, value : 32'h80215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820d, value : 32'h2000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820e, value : 32'h30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820f, value : 32'h70004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58210, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58211, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58212, value : 32'he0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58213, value : 32'h70001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58214, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58215, value : 32'habe0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58216, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58217, value : 32'ha0320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58218, value : 32'h30010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58219, value : 32'h40009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5821a, value : 32'h80004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824c, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824d, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824e, value : 32'h20043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824f, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58250, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58251, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58252, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58253, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58254, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58255, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58256, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58257, value : 32'h42b0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58258, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58259, value : 32'h300c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825a, value : 32'h10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825b, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825c, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825d, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825e, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825f, value : 32'h50004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58260, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58261, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58262, value : 32'h8550004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58263, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58264, value : 32'h40158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58265, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58266, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58267, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58268, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58269, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826a, value : 32'h80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826b, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826c, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826d, value : 32'hc800004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826e, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826f, value : 32'h601d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58270, value : 32'h20009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58271, value : 32'h30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58272, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58273, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58274, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58275, value : 32'hb0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58276, value : 32'h70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58277, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58278, value : 32'h10ab0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58279, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827a, value : 32'h70258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827b, value : 32'h3000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827c, value : 32'h30008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827d, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827e, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827f, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58280, value : 32'he0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58281, value : 32'h90003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58282, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58283, value : 32'h157c0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58284, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58285, value : 32'h902ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58286, value : 32'h4000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58287, value : 32'h4000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58288, value : 32'h60002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58289, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828a, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828b, value : 32'h100009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828c, value : 32'hb0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828d, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828e, value : 32'h19000006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828f, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58290, value : 32'hb03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58291, value : 32'h50013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58292, value : 32'h5000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58293, value : 32'h70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58294, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58295, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58296, value : 32'h16000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58297, value : 32'hf0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58298, value : 32'h20006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58299, value : 32'h21550008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829a, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829b, value : 32'he04b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829c, value : 32'h60018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829d, value : 32'h70010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829e, value : 32'h90002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829f, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a0, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a1, value : 32'h60006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a2, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a4, value : 32'h60001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a5, value : 32'h2150007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a6, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a7, value : 32'h8010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a8, value : 32'h80008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582aa, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ab, value : 32'h90007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ac, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ad, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ae, value : 32'ha000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582af, value : 32'h1000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b0, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b1, value : 32'h80002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b2, value : 32'h640000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b3, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b4, value : 32'hc0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b5, value : 32'he000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b6, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b7, value : 32'h30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b8, value : 32'hb0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b9, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ba, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bb, value : 32'h100010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bc, value : 32'h30012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bd, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582be, value : 32'ha0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bf, value : 32'habe000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c0, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c1, value : 32'h120320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c2, value : 32'h140014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c3, value : 32'h70005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c4, value : 32'h40007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c5, value : 32'he000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58300, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58301, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58302, value : 32'h30043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58303, value : 32'h30003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58305, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58306, value : 32'h40003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58307, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58308, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58309, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830a, value : 32'h4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830c, value : 32'h40001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830d, value : 32'h42b0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830e, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830f, value : 32'h500c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58310, value : 32'h50005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58311, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58312, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58313, value : 32'h50004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58314, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58315, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58316, value : 32'h70006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58317, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58318, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58319, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831a, value : 32'h8550006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831b, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831c, value : 32'h80158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831d, value : 32'h90008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831e, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831f, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58320, value : 32'h70005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58321, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58322, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58323, value : 32'ha0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58324, value : 32'h3000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58325, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58326, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58327, value : 32'hc800007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58328, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58329, value : 32'ha01d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832a, value : 32'hc000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832b, value : 32'h40003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832c, value : 32'h30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832d, value : 32'h80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832e, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832f, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58330, value : 32'hd000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58331, value : 32'h4000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58332, value : 32'h60005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58333, value : 32'h60003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58334, value : 32'h10ab0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58335, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58336, value : 32'hd0258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58337, value : 32'hf000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58338, value : 32'h60005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58339, value : 32'h30007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833a, value : 32'h90006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833b, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833c, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833d, value : 32'h10000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833e, value : 32'h60011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833f, value : 32'h80007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58340, value : 32'h60004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58341, value : 32'h157c000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58342, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58343, value : 32'h1002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58344, value : 32'h130011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58345, value : 32'h70006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58346, value : 32'h40009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58347, value : 32'hb0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58348, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58349, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834a, value : 32'h120011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834b, value : 32'h70014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834c, value : 32'ha0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834d, value : 32'h70004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834e, value : 32'h1900000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834f, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58350, value : 32'h1403aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58351, value : 32'h180016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58352, value : 32'h90007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58353, value : 32'h5000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58354, value : 32'he0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58355, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58356, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58357, value : 32'h190017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58358, value : 32'h8001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58359, value : 32'hb000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835a, value : 32'ha0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835b, value : 32'h21550010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835c, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835d, value : 32'h1904b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835e, value : 32'h1d001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835f, value : 32'hb0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58360, value : 32'h7000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58361, value : 32'h12000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58362, value : 32'ha05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58363, value : 32'h50000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58364, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58365, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58366, value : 32'h43416564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58367, value : 32'h63500030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58368, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58369, value : 32'h646f4341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836a, value : 32'h53514465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836b, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836c, value : 32'h4143446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836d, value : 32'h65646f43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836e, value : 32'h314341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836f, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58370, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58371, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58372, value : 32'h30434174},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58373, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58374, value : 32'h4443446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58375, value : 32'h7366664f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58376, value : 32'h43417465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58377, value : 32'h63500031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58378, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58379, value : 32'h66664f44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837a, value : 32'h44746573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837b, value : 32'h50005351},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837c, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837d, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837e, value : 32'h71446564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837f, value : 32'h306e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58380, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58381, value : 32'h43414344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58382, value : 32'h4465646f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58383, value : 32'h316e4c71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58384, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58385, value : 32'h4143446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58386, value : 32'h65646f43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58387, value : 32'h6e4c7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58388, value : 32'h63500032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58389, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838a, value : 32'h646f4341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838b, value : 32'h4c714465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838c, value : 32'h5000336e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838d, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838e, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838f, value : 32'h71446564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58390, value : 32'h346e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58391, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58392, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58393, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58394, value : 32'h4c714474},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58395, value : 32'h5000306e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58396, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58397, value : 32'h664f4443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58398, value : 32'h74657366},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58399, value : 32'h6e4c7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839a, value : 32'h63500031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839b, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839c, value : 32'h66664f44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839d, value : 32'h44746573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839e, value : 32'h326e4c71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839f, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a0, value : 32'h4443446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a1, value : 32'h7366664f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a2, value : 32'h71447465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a3, value : 32'h336e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a4, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a5, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a6, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a7, value : 32'h4c714474},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a8, value : 32'h346e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a9, value : 32'h4050607},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583aa, value : 32'h10203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ab, value : 32'hc0b0a09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ac, value : 32'hb50f0e0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ad, value : 32'h1ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ae, value : 32'h1f0b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583af, value : 32'hb3000100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b0, value : 32'h1f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b1, value : 32'h1f0b400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b2, value : 32'hb0000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b3, value : 32'h300001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b4, value : 32'h7f00300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b5, value : 32'h4000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b6, value : 32'h7f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b7, value : 32'h1fe0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b8, value : 32'h4000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b9, value : 32'h1fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ba, value : 32'h7f01100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bb, value : 32'h21000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bc, value : 32'h1fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bd, value : 32'h1ffbe00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583be, value : 32'hbe000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bf, value : 32'h10001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c0, value : 32'h1f0a700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c1, value : 32'ha2000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c2, value : 32'h20001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c3, value : 32'h2007900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c4, value : 32'h4000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c5, value : 32'h1008b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c6, value : 32'hf05f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c7, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c8, value : 32'h1ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c9, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ca, value : 32'h1ff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cb, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cc, value : 32'hf0b001ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cd, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ce, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cf, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d0, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d1, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d2, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d3, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d4, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d5, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d6, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d7, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d8, value : 32'hf0a70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d9, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583da, value : 32'he000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583db, value : 32'hc000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583dc, value : 32'ha000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583dd, value : 32'h80009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583de, value : 32'h60007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583df, value : 32'h40005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e0, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e1, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e2, value : 32'h110010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e3, value : 32'h130012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e4, value : 32'h150014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e5, value : 32'h170016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e6, value : 32'h190018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e7, value : 32'h1b001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e8, value : 32'h1d001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e9, value : 32'h1f001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ea, value : 32'hef77dbb7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583eb, value : 32'hfbdff7bd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ec, value : 32'hbddfb76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ed, value : 32'hbdffbdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ee, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ef, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f0, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f1, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f2, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f3, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f4, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f5, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f6, value : 32'h1ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f7, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f8, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f9, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fa, value : 32'hf0b90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fb, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fc, value : 32'h1f0ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fd, value : 32'hf0b10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fe, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ff, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58400, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58401, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58402, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58403, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58404, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58405, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58406, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58407, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58408, value : 32'h7f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58409, value : 32'hfe200002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840a, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840b, value : 32'h7f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840c, value : 32'hf01cffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840d, value : 32'hffff0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840e, value : 32'h1fe2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840f, value : 32'hfe2bffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58410, value : 32'hffff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58411, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58412, value : 32'hffb50040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58413, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58414, value : 32'h1f0b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58415, value : 32'hf0b40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58416, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58417, value : 32'h1f0b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58418, value : 32'hf0ba0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58419, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841a, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841b, value : 32'hf0b00002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841c, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841d, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841e, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841f, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58420, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58421, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58422, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58423, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58424, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58425, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58426, value : 32'h7f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58427, value : 32'hfe200002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58428, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58429, value : 32'h7f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842a, value : 32'hf01cffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842b, value : 32'hffff0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842c, value : 32'h1fe2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842d, value : 32'hfe2bffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842e, value : 32'hffff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842f, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58430, value : 32'h40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58431, value : 32'h8840884},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58432, value : 32'h20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58433, value : 32'h10010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58434, value : 32'h10012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58435, value : 32'h1007a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58436, value : 32'h10028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58437, value : 32'h60000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58438, value : 32'h50005000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58439, value : 32'h2008050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843b, value : 32'h60080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843c, value : 32'h3c5a5555},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843d, value : 32'h600000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58440, value : 32'h70},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58441, value : 32'h75},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58442, value : 32'h26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58443, value : 32'ha0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58444, value : 32'ha1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58445, value : 32'ha4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58446, value : 32'ha5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58447, value : 32'ha030201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58448, value : 32'he0d0c0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58449, value : 32'h1413120f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844a, value : 32'h18171615},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844b, value : 32'h1e1c1a19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844c, value : 32'h2221201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844d, value : 32'h2e292825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844e, value : 32'h4746453a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844f, value : 32'h4a4948},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1}, //This allows the firmware unrestricted access to the configuration CSRs.
//[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
// [dwc_ddrphy_phyinit_F_loadDMEM1D] End of dwc_ddrphy_phyinit_F_loadDMEM, Pstate=2
// [dwc_ddrphy_phyinit_G_execFW] Start of dwc_ddrphy_phyinit_G_execFW
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1}, ////     Then rewrite the CSR so that only the StallToMicro remains set (all other fields should be zero).
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h9}, //[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h0}, // [dwc_ddrphy_phyinit_userCustom_G_waitFwDone] Start of dwc_ddrphy_phyinit_userCustom_G_waitFwDone()
// [dwc_ddrphy_phyinit_userCustom_G_waitFwDone] End of dwc_ddrphy_phyinit_userCustom_G_waitFwDone()
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h1}, //// 4.   Halt the microcontroller."
// [dwc_ddrphy_phyinit_G_execFW] End of dwc_ddrphy_phyinit_G_execFW
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}, // [dwc_ddrphy_phyinit_userCustom_H_readMsgBlock] Start of dwc_ddrphy_phyinit_userCustom_H_readMsgBlock()
// [dwc_ddrphy_phyinit_userCustom_H_readMsgBlock] End of dwc_ddrphy_phyinit_userCustom_H_readMsgBlock ()
// 3. If training is required at another frequency, repeat the operations starting at step (E).
// [dwc_ddrphy_phyinit_H_readMsgBlock] End of dwc_ddrphy_phyinit_H_readMsgBlock
//[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Start of dwc_ddrphy_phyinit_I_loadPIEImagePsLoop(), PState=2
                          '{ step_type : REG_WRITE, reg_addr : 32'h260008, value : 32'h4956}, //[dwc_ddrphy_phyinit_programPLL] [phyinit_I_loadPIEImagePsLoop] Pstate=2,  Memclk=400MHz, Programming CpllCtrl5 to 0x4956.
                          '{ step_type : REG_WRITE, reg_addr : 32'h60006, value : 32'h3f0}, //End of dwc_ddrphy_phyinit_programPLL(), PState=2
                          '{ step_type : REG_WRITE, reg_addr : 32'h230015, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h231015, value : 32'h0}, //phyinit_io_write: 0x230015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21007c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21107c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21207c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21307c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21007c, value : 32'h0}, //phyinit_io_write: 0x21307c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21107c, value : 32'h0}, //phyinit_io_write: 0x21007c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21207c, value : 32'h0}, //phyinit_io_write: 0x21107c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21307c, value : 32'h0}, //phyinit_io_write: 0x21207c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h230015, value : 32'h0}, //phyinit_io_write: 0x21307c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h231015, value : 32'h0}, //phyinit_io_write: 0x230015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h270141, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming ACSMWckFreeRunMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h29080c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming GPR12 with Zcalkclkdiv to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h210027, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming RxClkCntl1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h211027, value : 32'h0}, //phyinit_io_write: 0x210027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h212027, value : 32'h0}, //phyinit_io_write: 0x211027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h213027, value : 32'h0}, //phyinit_io_write: 0x212027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h21020f, value : 32'h8}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=2, Programming RxReplicaCtl04 to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h21120f, value : 32'h8}, //phyinit_io_write: 0x21020f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h21220f, value : 32'h8}, //phyinit_io_write: 0x21120f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h21320f, value : 32'h8}, //phyinit_io_write: 0x21220f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e003f, value : 32'h0}, //phyinit_io_write: 0x21320f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e008d, value : 32'h0}, //phyinit_io_write: 0x2e003f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e103f, value : 32'h0}, //phyinit_io_write: 0x2e008d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e108d, value : 32'h0}, //phyinit_io_write: 0x2e103f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e203f, value : 32'h0}, //phyinit_io_write: 0x2e108d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e208d, value : 32'h0}, //phyinit_io_write: 0x2e203f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e303f, value : 32'h0}, //phyinit_io_write: 0x2e208d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e308d, value : 32'h0}, //phyinit_io_write: 0x2e303f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e403f, value : 32'h0}, //phyinit_io_write: 0x2e308d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e408d, value : 32'h0}, //phyinit_io_write: 0x2e403f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e503f, value : 32'h0}, //phyinit_io_write: 0x2e408d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e508d, value : 32'h0}, //phyinit_io_write: 0x2e503f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e603f, value : 32'h0}, //phyinit_io_write: 0x2e508d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e608d, value : 32'h0}, //phyinit_io_write: 0x2e603f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e703f, value : 32'h0}, //phyinit_io_write: 0x2e608d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h2e708d, value : 32'h0}, //phyinit_io_write: 0x2e703f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h290903, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] PState=2, Programming RtrnMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70072, value : 32'h3}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming HwtLpCsEnA to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h29080e, value : 32'h3}, //phyinit_io_write: 0x70072, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h70073, value : 32'h3}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming HwtLpCsEnB to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h29080f, value : 32'h3}, //phyinit_io_write: 0x70073, 0x3
//phyinit_io_write: 0x29080f, 0x3
//[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] End of dwc_ddrphy_phyinit_I_loadPIEImagePsLoop(), PState=2
//[dwc_ddrphy_phyinit_userCustom_customPostTrainPsLoop] End of dwc_ddrphy_phyinit_userCustom_customPostTrainPsLoop(), PState=2
//Start of dwc_ddrphy_phyinit_C_initPhyConfigPsLoop(), PState=3, tck_ps=5000ps
                          '{ step_type : REG_WRITE, reg_addr : 32'h2008b, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, programming PState = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h390801, value : 32'h8692}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming Seq0BGPR1 to 0x8692
                          '{ step_type : REG_WRITE, reg_addr : 32'h390802, value : 32'h0}, //phyinit_io_write: 0x390801, 0x8692
                          '{ step_type : REG_WRITE, reg_addr : 32'h390806, value : 32'h1}, //phyinit_io_write: 0x390802, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3a03ff, value : 32'h4101}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming OdtSeg120 to 0x4101
                          '{ step_type : REG_WRITE, reg_addr : 32'h3a030b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming ZCalCompCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h360008, value : 32'h4962}, //[dwc_ddrphy_phyinit_programPLL] [phyinit_C_initPhyConfigPsLoop] Pstate=3,  Memclk=200MHz, Programming CpllCtrl5 to 0x4962.
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908e0, value : 32'h19}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY0 to 0x19 (0.5us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908e1, value : 32'h4b}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY1 to 0x4b (tZQCal PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908e2, value : 32'h1f4}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY2 to 0x1f4 (10.us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908e3, value : 32'h40}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY3 to 0x40 (dllLock PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908e4, value : 32'h5}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY4 to 0x5 (0.1us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908e5, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY5 to 0x0 (RxReplicaCalWait delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908e6, value : 32'h43}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY6 to 0x43 (Oscillator PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908e7, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY7 to 0x0 (tXDSM_XP PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908ea, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY10 to 0x1 (tPDXCSODTON 20ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908eb, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY11 to 0x1 (20ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908ec, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY12 to 0x3 (50ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h3908ed, value : 32'h14}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming Seq0BDLY13 to 0x14 (tXSR PIE delay, tRFCab delay is 380ns)
                          '{ step_type : REG_WRITE, reg_addr : 32'h320002, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming PclkPtrInitVal to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h360040, value : 32'h3}, //phyinit_io_write: 0x320002, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h320000, value : 32'h2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DfiFreqRatio to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h3100fb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming RxDigStrbEn to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3110fb, value : 32'h0}, //phyinit_io_write: 0x3100fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3120fb, value : 32'h0}, //phyinit_io_write: 0x3110fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3130fb, value : 32'h0}, //phyinit_io_write: 0x3120fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e000b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DxDigStrobeMode HMDBYTE to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e100b, value : 32'h0}, //phyinit_io_write: 0x3e000b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e200b, value : 32'h0}, //phyinit_io_write: 0x3e100b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e300b, value : 32'h0}, //phyinit_io_write: 0x3e200b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e400b, value : 32'h0}, //phyinit_io_write: 0x3e300b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e500b, value : 32'h0}, //phyinit_io_write: 0x3e400b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e600b, value : 32'h0}, //phyinit_io_write: 0x3e500b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e700b, value : 32'h0}, //phyinit_io_write: 0x3e600b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h310024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE0.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h311024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE1.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h312024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE2.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h313024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE3.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h310025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE0.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h311025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE1.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h312025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE2.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h313025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE3.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h310004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE0.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h310003, value : 32'h0}, //phyinit_io_write: 0x310004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h311004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE1.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h311003, value : 32'h0}, //phyinit_io_write: 0x311004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h312004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE2.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h312003, value : 32'h0}, //phyinit_io_write: 0x312004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h313004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE3.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h313003, value : 32'h0}, //phyinit_io_write: 0x313004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3b0004, value : 32'hc8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ZCalClkInfo::ZCalDfiClkTicksPer1uS to 0xc8
                          '{ step_type : REG_WRITE, reg_addr : 32'h3a030c, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h31003e, value : 32'h5}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE RxGainCurrAdjRxReplica to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h31103e, value : 32'h5}, //phyinit_io_write: 0x31003e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h31203e, value : 32'h5}, //phyinit_io_write: 0x31103e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h31303e, value : 32'h5}, //phyinit_io_write: 0x31203e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h320003, value : 32'h1}, //phyinit_io_write: 0x31303e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h32000b, value : 32'h1111}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming CPclkDivRatio to 0x1111
                          '{ step_type : REG_WRITE, reg_addr : 32'h310108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE0.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h311108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE1.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h312108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE2.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h313108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming DBYTE3.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70005, value : 32'h0}, //[phyinit_C_initPhyConfig] Programming EnPhyUpdZQCalUpdate to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h7000f, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming DisableZQupdateOnSnoop to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31000e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h31100e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h31200e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h31300e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h320019, value : 32'h4}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming EnRxDqsTracking::DqsSampNegRxEnSense to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e002c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 0 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e102c, value : 32'h33}, //phyinit_io_write: 0x3e002c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e002d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 0 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e102d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 0 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e202c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 1 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e302c, value : 32'h33}, //phyinit_io_write: 0x3e202c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e202d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 1 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e302d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 1 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e402c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 2 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e502c, value : 32'h33}, //phyinit_io_write: 0x3e402c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e402d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 2 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e502d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 2 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e602c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 3 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e702c, value : 32'h33}, //phyinit_io_write: 0x3e602c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e602d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 3 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e702d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 3 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h300070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC0 Instance0 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h301070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC1 Instance1 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h302070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC2 Instance2 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h303070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC3 Instance3 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h304070, value : 32'hff}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming AC0 HMAC4 Instance4 CS TxImpedanceAC::TxStrenCodePDAC to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h305070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC5 Instance5 TxImpedanceAC::TxStrenCodePD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h307070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC0 Instance7 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h308070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC1 Instance8 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h309070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC2 Instance9 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h30a070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC3 Instance10 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h30b070, value : 32'hff}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming AC1 HMAC4 Instance11 CS TxImpedanceAC::TxStrenCodePDAC to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h30c070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC5 Instance12 TxImpedanceAC::TxStrenCodePD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e002e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 0 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e102e, value : 32'h30}, //phyinit_io_write: 0x3e002e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e002f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 0 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e102f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 0 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e202e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 1 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e302e, value : 32'h30}, //phyinit_io_write: 0x3e202e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e202f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 1 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e302f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 1 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e402e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 2 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e502e, value : 32'h30}, //phyinit_io_write: 0x3e402e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e402f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 2 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e502f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 2 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e602e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 3 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e702e, value : 32'h30}, //phyinit_io_write: 0x3e602e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e602f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 3 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e702f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 3 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h300079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC0 Instance0 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h301079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC1 Instance1 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h302079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC2 Instance2 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h303079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC3 Instance3 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h304079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC4 Instance4 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h305079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC5 DIFF5 OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h307079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC0 Instance7 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h308079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC1 Instance8 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h309079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC2 Instance9 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h30a079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC3 Instance10 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h30b079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC4 Instance11 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h30c079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC5 DIFF12 OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e001c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 0 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e101c, value : 32'h3}, //phyinit_io_write: 0x3e001c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e201c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 1 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e301c, value : 32'h3}, //phyinit_io_write: 0x3e201c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e401c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 2 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e501c, value : 32'h3}, //phyinit_io_write: 0x3e401c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e601c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming HMDBYTE 3 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e701c, value : 32'h3}, //phyinit_io_write: 0x3e601c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h30006d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC0 Instance0 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30106d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC1 Instance1 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30206d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC2 Instance2 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30306d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC3 Instance3 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30406d, value : 32'hf8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC4 Instance4 CS TxSlewAC::TxSlewPDAC to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h30506d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX0 HMAC5 Instance5 TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30706d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC0 Instance7 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30806d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC1 Instance8 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30906d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC2 Instance9 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30a06d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC3 Instance10 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30b06d, value : 32'hf8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC4 Instance11 CS TxSlewAC::TxSlewPDAC to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h30c06d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACX1 HMAC5 Instance12 TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e003e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Programming HMDBYTE RxDQSCtrl::RxDQSDiffSeVrefDACEn to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e103e, value : 32'h0}, //phyinit_io_write: 0x3e003e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e203e, value : 32'h0}, //phyinit_io_write: 0x3e103e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e303e, value : 32'h0}, //phyinit_io_write: 0x3e203e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e403e, value : 32'h0}, //phyinit_io_write: 0x3e303e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e503e, value : 32'h0}, //phyinit_io_write: 0x3e403e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e603e, value : 32'h0}, //phyinit_io_write: 0x3e503e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e703e, value : 32'h0}, //phyinit_io_write: 0x3e603e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h310001, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming WriteLinkEcc to 0
                          '{ step_type : REG_WRITE, reg_addr : 32'h311001, value : 32'h0}, //phyinit_io_write: 0x310001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h312001, value : 32'h0}, //phyinit_io_write: 0x311001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h313001, value : 32'h0}, //phyinit_io_write: 0x312001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h370040, value : 32'h5a}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming PPTTrainSetup::PhyMstrMaxReqToAck to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h370041, value : 32'hf}, //phyinit_io_write: 0x370040, 0x5a
                          '{ step_type : REG_WRITE, reg_addr : 32'h3100a5, value : 32'h1}, //phyinit_io_write: 0x370041, 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h3110a5, value : 32'h1}, //phyinit_io_write: 0x3100a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3120a5, value : 32'h1}, //phyinit_io_write: 0x3110a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3130a5, value : 32'h1}, //phyinit_io_write: 0x3120a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h310209, value : 32'h3232}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Programming RxReplicaRangeVal 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h311209, value : 32'h3232}, //phyinit_io_write: 0x310209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h312209, value : 32'h3232}, //phyinit_io_write: 0x311209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h313209, value : 32'h3232}, //phyinit_io_write: 0x312209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h31020f, value : 32'h6}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Programming RxReplicaCtl04 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h31120f, value : 32'h6}, //phyinit_io_write: 0x31020f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h31220f, value : 32'h6}, //phyinit_io_write: 0x31120f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h31320f, value : 32'h6}, //phyinit_io_write: 0x31220f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h320005, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, DfiFreq=200MHz, Programming PipeCtl[AcInPipeEn]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h310008, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, DfiFreq=200MHz, Programming DBYTE0.LP5DfiDataEnLatency[LP5RLm13]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h311008, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, DfiFreq=200MHz, Programming DBYTE1.LP5DfiDataEnLatency[LP5RLm13]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h312008, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, DfiFreq=200MHz, Programming DBYTE2.LP5DfiDataEnLatency[LP5RLm13]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h313008, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, DfiFreq=200MHz, Programming DBYTE3.LP5DfiDataEnLatency[LP5RLm13]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h37006b, value : 32'h222}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, DfiFreq=200MHz, Programming DfiHandshakeDelays[PhyUpdReqDelay]=0x2 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h370066, value : 32'h20}, //phyinit_io_write: 0x37006b, 0x222
                          '{ step_type : REG_WRITE, reg_addr : 32'h3700eb, value : 32'h222}, //phyinit_io_write: 0x370066, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h3700e6, value : 32'h20}, //phyinit_io_write: 0x3700eb, 0x222
                          '{ step_type : REG_WRITE, reg_addr : 32'h370135, value : 32'h400}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACSMWckWriteFastTogglePulse::ACSMWckWriteFastToggleWidth to 0x19, ACSMWckWriteFastTogglePulse::ACSMWckWriteFastToggleDelay to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h370136, value : 32'h400}, //phyinit_io_write: 0x370135, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h370137, value : 32'h404}, //phyinit_io_write: 0x370136, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h370138, value : 32'h1908}, //phyinit_io_write: 0x370137, 0x404
                          '{ step_type : REG_WRITE, reg_addr : 32'h370139, value : 32'h400}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACSMWckReadFastTogglePulse::ACSMWckReadFastToggleWidth to 0x21, ACSMWckReadFastTogglePulse::ACSMWckReadFastToggleDelay to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h37013a, value : 32'h400}, //phyinit_io_write: 0x370139, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h37013b, value : 32'h404}, //phyinit_io_write: 0x37013a, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h37013c, value : 32'h2108}, //phyinit_io_write: 0x37013b, 0x404
                          '{ step_type : REG_WRITE, reg_addr : 32'h37013d, value : 32'h400}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACSMWckFreqFastTogglePulse::ACSMWckFreqFastToggleWidth to 0x11, ACSMWckFreqFastTogglePulse::ACSMWckFreqFastToggleDelay to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h37013e, value : 32'h400}, //phyinit_io_write: 0x37013d, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h37013f, value : 32'h404}, //phyinit_io_write: 0x37013e, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h370140, value : 32'h1108}, //phyinit_io_write: 0x37013f, 0x404
                          '{ step_type : REG_WRITE, reg_addr : 32'h37012c, value : 32'h80f}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACSMRxValPulse::ACSMRxValDelay to 0xf, ACSMRxValPulse::ACSMRxValWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h37012d, value : 32'h80f}, //phyinit_io_write: 0x37012c, 0x80f
                          '{ step_type : REG_WRITE, reg_addr : 32'h370130, value : 32'h80f}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACSMRdcsPulse::ACSMRdcsDelay to 0xf, ACSMRdcsPulse::ACSMRdcsWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h37012e, value : 32'h807}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACSMTxEnPulse::ACSMTxEnDelay to 0x7, ACSMTxEnPulse::ACSMTxEnWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h37012f, value : 32'h807}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming ACSMWrcsPulse::ACSMWrcsDelay to 0x7, ACSMWrcsPulse::ACSMWrcsWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h330008, value : 32'h0}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming AcPipeEn AC0 to 0. DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h331008, value : 32'h0}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, Programming AcPipeEn AC1 to 0. DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e0013, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Programming csr_EnaRxStrobeEnB to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e1013, value : 32'h1}, //phyinit_io_write: 0x3e0013, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e2013, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Programming csr_EnaRxStrobeEnB to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e3013, value : 32'h1}, //phyinit_io_write: 0x3e2013, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e4013, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Programming csr_EnaRxStrobeEnB to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e5013, value : 32'h1}, //phyinit_io_write: 0x3e4013, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e6013, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Programming csr_EnaRxStrobeEnB to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e7013, value : 32'h1}, //phyinit_io_write: 0x3e6013, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e0002, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Programming HMDBYTE RxDFECtrlDq to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e1002, value : 32'h0}, //phyinit_io_write: 0x3e0002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e2002, value : 32'h0}, //phyinit_io_write: 0x3e1002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e3002, value : 32'h0}, //phyinit_io_write: 0x3e2002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e4002, value : 32'h0}, //phyinit_io_write: 0x3e3002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e5002, value : 32'h0}, //phyinit_io_write: 0x3e4002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e6002, value : 32'h0}, //phyinit_io_write: 0x3e5002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e7002, value : 32'h0}, //phyinit_io_write: 0x3e6002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31010b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=3, Memclk=200MHz, freqThreshold=200MHz, NoRDQS=0 Programming InhibitTxRdPtrInit::DisableRxEnDlyLoad to 0x0, InhibitTxRdPtrInit::DisableTxDqDly to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31110b, value : 32'h0}, //phyinit_io_write: 0x31010b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31210b, value : 32'h0}, //phyinit_io_write: 0x31110b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31310b, value : 32'h0}, //phyinit_io_write: 0x31210b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h300063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC0 Instance0 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h301063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC1 Instance1 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h302063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC2 Instance2 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h303063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC3 Instance3 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h304063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC4 Instance4 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h305063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC5 Instance5 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h307063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC0 Instance7 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h308063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC1 Instance8 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h309063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC2 Instance9 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h30a063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC3 Instance10 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h30b063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC4 Instance11 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h30c063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC5 Instance12 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h39080a, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Programming Seq0BGPR10 to HMTxLcdlSeed Full search value = 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h39080b, value : 32'h2d0}, //phyinit_io_write: 0x39080a, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h390815, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Programming Seq0BGPR21 to ACHMTxLcdlSeed Full search value = 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h390816, value : 32'h2d0}, //phyinit_io_write: 0x390815, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e0063, value : 32'h2d0}, //phyinit_io_write: 0x390816, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e0064, value : 32'h2d0}, //phyinit_io_write: 0x3e0063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e0087, value : 32'h2d0}, //phyinit_io_write: 0x3e0064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e1063, value : 32'h2d0}, //phyinit_io_write: 0x3e0087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e1064, value : 32'h2d0}, //phyinit_io_write: 0x3e1063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e1087, value : 32'h2d0}, //phyinit_io_write: 0x3e1064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e2063, value : 32'h2d0}, //phyinit_io_write: 0x3e1087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e2064, value : 32'h2d0}, //phyinit_io_write: 0x3e2063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e2087, value : 32'h2d0}, //phyinit_io_write: 0x3e2064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e3063, value : 32'h2d0}, //phyinit_io_write: 0x3e2087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e3064, value : 32'h2d0}, //phyinit_io_write: 0x3e3063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e3087, value : 32'h2d0}, //phyinit_io_write: 0x3e3064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e4063, value : 32'h2d0}, //phyinit_io_write: 0x3e3087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e4064, value : 32'h2d0}, //phyinit_io_write: 0x3e4063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e4087, value : 32'h2d0}, //phyinit_io_write: 0x3e4064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e5063, value : 32'h2d0}, //phyinit_io_write: 0x3e4087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e5064, value : 32'h2d0}, //phyinit_io_write: 0x3e5063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e5087, value : 32'h2d0}, //phyinit_io_write: 0x3e5064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e6063, value : 32'h2d0}, //phyinit_io_write: 0x3e5087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e6064, value : 32'h2d0}, //phyinit_io_write: 0x3e6063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e6087, value : 32'h2d0}, //phyinit_io_write: 0x3e6064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e7063, value : 32'h2d0}, //phyinit_io_write: 0x3e6087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e7064, value : 32'h2d0}, //phyinit_io_write: 0x3e7063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e7087, value : 32'h2d0}, //phyinit_io_write: 0x3e7064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0080, value : 32'h7}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming UcclkHclkEnables to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e003c, value : 32'h80}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming RxDQSSeVrefDAC0 to 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e103c, value : 32'h80}, //phyinit_io_write: 0x3e003c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e203c, value : 32'h80}, //phyinit_io_write: 0x3e103c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e303c, value : 32'h80}, //phyinit_io_write: 0x3e203c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e403c, value : 32'h80}, //phyinit_io_write: 0x3e303c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e503c, value : 32'h80}, //phyinit_io_write: 0x3e403c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e603c, value : 32'h80}, //phyinit_io_write: 0x3e503c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e703c, value : 32'h80}, //phyinit_io_write: 0x3e603c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h390817, value : 32'h14}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 3 Seq0BGPR23 to 0x14, NumMemClk_tRFCab=82.0, NumMemClk_7p5ns=1.5, NumMemClk_tXSR=84.0
                          '{ step_type : REG_WRITE, reg_addr : 32'h390818, value : 32'h0}, //phyinit_io_write: 0x390817, 0x14
                          '{ step_type : REG_WRITE, reg_addr : 32'h390819, value : 32'h0}, //phyinit_io_write: 0x390818, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3300eb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 3 AC0 AcLcdlUpdInterval to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3310eb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 3 AC1 AcLcdlUpdInterval to 0x0
//[dwc_ddrphy_phyinit_programDfiMode] Skip DfiMode Programming: Keeping the reset value of 0x3
//End of dwc_ddrphy_phyinit_C_initPhyConfigPsLoop(), Pstate=3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3300d9, value : 32'h40}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming CKXTxDly to 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3300d8, value : 32'h40}, //phyinit_io_write: 0x3300d9, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3301d8, value : 32'h40}, //phyinit_io_write: 0x3300d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3302d8, value : 32'h40}, //phyinit_io_write: 0x3301d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3303d8, value : 32'h40}, //phyinit_io_write: 0x3302d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3304d8, value : 32'h40}, //phyinit_io_write: 0x3303d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3305d8, value : 32'h40}, //phyinit_io_write: 0x3304d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3306d8, value : 32'h40}, //phyinit_io_write: 0x3305d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3308d8, value : 32'h40}, //phyinit_io_write: 0x3306d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3309d8, value : 32'h40}, //phyinit_io_write: 0x3308d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3310d9, value : 32'h40}, //phyinit_io_write: 0x3309d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3310d8, value : 32'h40}, //phyinit_io_write: 0x3310d9, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3311d8, value : 32'h40}, //phyinit_io_write: 0x3310d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3312d8, value : 32'h40}, //phyinit_io_write: 0x3311d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3313d8, value : 32'h40}, //phyinit_io_write: 0x3312d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3314d8, value : 32'h40}, //phyinit_io_write: 0x3313d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3315d8, value : 32'h40}, //phyinit_io_write: 0x3314d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3316d8, value : 32'h40}, //phyinit_io_write: 0x3315d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3318d8, value : 32'h40}, //phyinit_io_write: 0x3316d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h3319d8, value : 32'h40}, //phyinit_io_write: 0x3318d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h310000, value : 32'h5}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming HwtMRL to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h311000, value : 32'h5}, //phyinit_io_write: 0x310000, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h312000, value : 32'h5}, //phyinit_io_write: 0x311000, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h313000, value : 32'h5}, //phyinit_io_write: 0x312000, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h37000d, value : 32'h5}, //phyinit_io_write: 0x313000, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h31002a, value : 32'h200}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming TxWckDlyTg0/Tg1 to 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h31002b, value : 32'h200}, //phyinit_io_write: 0x31002a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h31102a, value : 32'h200}, //phyinit_io_write: 0x31002b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h31102b, value : 32'h200}, //phyinit_io_write: 0x31102a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h31202a, value : 32'h200}, //phyinit_io_write: 0x31102b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h31202b, value : 32'h200}, //phyinit_io_write: 0x31202a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h31302a, value : 32'h200}, //phyinit_io_write: 0x31202b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h31302b, value : 32'h200}, //phyinit_io_write: 0x31302a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h310028, value : 32'h54}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming TxDqsDlyTg0/Tg1 to 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h310029, value : 32'h54}, //phyinit_io_write: 0x310028, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h311028, value : 32'h54}, //phyinit_io_write: 0x310029, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h311029, value : 32'h54}, //phyinit_io_write: 0x311028, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h312028, value : 32'h54}, //phyinit_io_write: 0x311029, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h312029, value : 32'h54}, //phyinit_io_write: 0x312028, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h313028, value : 32'h54}, //phyinit_io_write: 0x312029, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h313029, value : 32'h54}, //phyinit_io_write: 0x313028, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31007a, value : 32'h54}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming TxDqDlyTg0/Tg1 to 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31007b, value : 32'h54}, //phyinit_io_write: 0x31007a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31017a, value : 32'h54}, //phyinit_io_write: 0x31007b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31017b, value : 32'h54}, //phyinit_io_write: 0x31017a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31027a, value : 32'h54}, //phyinit_io_write: 0x31017b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31027b, value : 32'h54}, //phyinit_io_write: 0x31027a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31037a, value : 32'h54}, //phyinit_io_write: 0x31027b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31037b, value : 32'h54}, //phyinit_io_write: 0x31037a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31047a, value : 32'h54}, //phyinit_io_write: 0x31037b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31047b, value : 32'h54}, //phyinit_io_write: 0x31047a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31057a, value : 32'h54}, //phyinit_io_write: 0x31047b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31057b, value : 32'h54}, //phyinit_io_write: 0x31057a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31067a, value : 32'h54}, //phyinit_io_write: 0x31057b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31067b, value : 32'h54}, //phyinit_io_write: 0x31067a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31077a, value : 32'h54}, //phyinit_io_write: 0x31067b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31077b, value : 32'h54}, //phyinit_io_write: 0x31077a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31087a, value : 32'h54}, //phyinit_io_write: 0x31077b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31087b, value : 32'h54}, //phyinit_io_write: 0x31087a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31107a, value : 32'h54}, //phyinit_io_write: 0x31087b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31107b, value : 32'h54}, //phyinit_io_write: 0x31107a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31117a, value : 32'h54}, //phyinit_io_write: 0x31107b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31117b, value : 32'h54}, //phyinit_io_write: 0x31117a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31127a, value : 32'h54}, //phyinit_io_write: 0x31117b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31127b, value : 32'h54}, //phyinit_io_write: 0x31127a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31137a, value : 32'h54}, //phyinit_io_write: 0x31127b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31137b, value : 32'h54}, //phyinit_io_write: 0x31137a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31147a, value : 32'h54}, //phyinit_io_write: 0x31137b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31147b, value : 32'h54}, //phyinit_io_write: 0x31147a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31157a, value : 32'h54}, //phyinit_io_write: 0x31147b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31157b, value : 32'h54}, //phyinit_io_write: 0x31157a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31167a, value : 32'h54}, //phyinit_io_write: 0x31157b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31167b, value : 32'h54}, //phyinit_io_write: 0x31167a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31177a, value : 32'h54}, //phyinit_io_write: 0x31167b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31177b, value : 32'h54}, //phyinit_io_write: 0x31177a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31187a, value : 32'h54}, //phyinit_io_write: 0x31177b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31187b, value : 32'h54}, //phyinit_io_write: 0x31187a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31207a, value : 32'h54}, //phyinit_io_write: 0x31187b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31207b, value : 32'h54}, //phyinit_io_write: 0x31207a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31217a, value : 32'h54}, //phyinit_io_write: 0x31207b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31217b, value : 32'h54}, //phyinit_io_write: 0x31217a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31227a, value : 32'h54}, //phyinit_io_write: 0x31217b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31227b, value : 32'h54}, //phyinit_io_write: 0x31227a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31237a, value : 32'h54}, //phyinit_io_write: 0x31227b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31237b, value : 32'h54}, //phyinit_io_write: 0x31237a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31247a, value : 32'h54}, //phyinit_io_write: 0x31237b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31247b, value : 32'h54}, //phyinit_io_write: 0x31247a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31257a, value : 32'h54}, //phyinit_io_write: 0x31247b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31257b, value : 32'h54}, //phyinit_io_write: 0x31257a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31267a, value : 32'h54}, //phyinit_io_write: 0x31257b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31267b, value : 32'h54}, //phyinit_io_write: 0x31267a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31277a, value : 32'h54}, //phyinit_io_write: 0x31267b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31277b, value : 32'h54}, //phyinit_io_write: 0x31277a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31287a, value : 32'h54}, //phyinit_io_write: 0x31277b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31287b, value : 32'h54}, //phyinit_io_write: 0x31287a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31307a, value : 32'h54}, //phyinit_io_write: 0x31287b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31307b, value : 32'h54}, //phyinit_io_write: 0x31307a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31317a, value : 32'h54}, //phyinit_io_write: 0x31307b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31317b, value : 32'h54}, //phyinit_io_write: 0x31317a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31327a, value : 32'h54}, //phyinit_io_write: 0x31317b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31327b, value : 32'h54}, //phyinit_io_write: 0x31327a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31337a, value : 32'h54}, //phyinit_io_write: 0x31327b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31337b, value : 32'h54}, //phyinit_io_write: 0x31337a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31347a, value : 32'h54}, //phyinit_io_write: 0x31337b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31347b, value : 32'h54}, //phyinit_io_write: 0x31347a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31357a, value : 32'h54}, //phyinit_io_write: 0x31347b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31357b, value : 32'h54}, //phyinit_io_write: 0x31357a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31367a, value : 32'h54}, //phyinit_io_write: 0x31357b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31367b, value : 32'h54}, //phyinit_io_write: 0x31367a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31377a, value : 32'h54}, //phyinit_io_write: 0x31367b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31377b, value : 32'h54}, //phyinit_io_write: 0x31377a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31387a, value : 32'h54}, //phyinit_io_write: 0x31377b, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h31387b, value : 32'h54}, //phyinit_io_write: 0x31387a, 0x54
                          '{ step_type : REG_WRITE, reg_addr : 32'h310078, value : 32'h286}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming RxDigStrbDlyTg0/Tg1 to 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310079, value : 32'h286}, //phyinit_io_write: 0x310078, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310178, value : 32'h286}, //phyinit_io_write: 0x310079, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310179, value : 32'h286}, //phyinit_io_write: 0x310178, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310278, value : 32'h286}, //phyinit_io_write: 0x310179, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310279, value : 32'h286}, //phyinit_io_write: 0x310278, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310378, value : 32'h286}, //phyinit_io_write: 0x310279, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310379, value : 32'h286}, //phyinit_io_write: 0x310378, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310478, value : 32'h286}, //phyinit_io_write: 0x310379, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310479, value : 32'h286}, //phyinit_io_write: 0x310478, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310578, value : 32'h286}, //phyinit_io_write: 0x310479, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310579, value : 32'h286}, //phyinit_io_write: 0x310578, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310678, value : 32'h286}, //phyinit_io_write: 0x310579, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310679, value : 32'h286}, //phyinit_io_write: 0x310678, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310778, value : 32'h286}, //phyinit_io_write: 0x310679, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310779, value : 32'h286}, //phyinit_io_write: 0x310778, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310878, value : 32'h286}, //phyinit_io_write: 0x310779, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310879, value : 32'h286}, //phyinit_io_write: 0x310878, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311078, value : 32'h286}, //phyinit_io_write: 0x310879, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311079, value : 32'h286}, //phyinit_io_write: 0x311078, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311178, value : 32'h286}, //phyinit_io_write: 0x311079, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311179, value : 32'h286}, //phyinit_io_write: 0x311178, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311278, value : 32'h286}, //phyinit_io_write: 0x311179, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311279, value : 32'h286}, //phyinit_io_write: 0x311278, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311378, value : 32'h286}, //phyinit_io_write: 0x311279, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311379, value : 32'h286}, //phyinit_io_write: 0x311378, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311478, value : 32'h286}, //phyinit_io_write: 0x311379, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311479, value : 32'h286}, //phyinit_io_write: 0x311478, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311578, value : 32'h286}, //phyinit_io_write: 0x311479, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311579, value : 32'h286}, //phyinit_io_write: 0x311578, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311678, value : 32'h286}, //phyinit_io_write: 0x311579, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311679, value : 32'h286}, //phyinit_io_write: 0x311678, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311778, value : 32'h286}, //phyinit_io_write: 0x311679, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311779, value : 32'h286}, //phyinit_io_write: 0x311778, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311878, value : 32'h286}, //phyinit_io_write: 0x311779, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h311879, value : 32'h286}, //phyinit_io_write: 0x311878, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312078, value : 32'h286}, //phyinit_io_write: 0x311879, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312079, value : 32'h286}, //phyinit_io_write: 0x312078, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312178, value : 32'h286}, //phyinit_io_write: 0x312079, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312179, value : 32'h286}, //phyinit_io_write: 0x312178, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312278, value : 32'h286}, //phyinit_io_write: 0x312179, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312279, value : 32'h286}, //phyinit_io_write: 0x312278, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312378, value : 32'h286}, //phyinit_io_write: 0x312279, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312379, value : 32'h286}, //phyinit_io_write: 0x312378, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312478, value : 32'h286}, //phyinit_io_write: 0x312379, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312479, value : 32'h286}, //phyinit_io_write: 0x312478, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312578, value : 32'h286}, //phyinit_io_write: 0x312479, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312579, value : 32'h286}, //phyinit_io_write: 0x312578, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312678, value : 32'h286}, //phyinit_io_write: 0x312579, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312679, value : 32'h286}, //phyinit_io_write: 0x312678, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312778, value : 32'h286}, //phyinit_io_write: 0x312679, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312779, value : 32'h286}, //phyinit_io_write: 0x312778, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312878, value : 32'h286}, //phyinit_io_write: 0x312779, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h312879, value : 32'h286}, //phyinit_io_write: 0x312878, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313078, value : 32'h286}, //phyinit_io_write: 0x312879, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313079, value : 32'h286}, //phyinit_io_write: 0x313078, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313178, value : 32'h286}, //phyinit_io_write: 0x313079, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313179, value : 32'h286}, //phyinit_io_write: 0x313178, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313278, value : 32'h286}, //phyinit_io_write: 0x313179, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313279, value : 32'h286}, //phyinit_io_write: 0x313278, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313378, value : 32'h286}, //phyinit_io_write: 0x313279, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313379, value : 32'h286}, //phyinit_io_write: 0x313378, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313478, value : 32'h286}, //phyinit_io_write: 0x313379, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313479, value : 32'h286}, //phyinit_io_write: 0x313478, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313578, value : 32'h286}, //phyinit_io_write: 0x313479, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313579, value : 32'h286}, //phyinit_io_write: 0x313578, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313678, value : 32'h286}, //phyinit_io_write: 0x313579, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313679, value : 32'h286}, //phyinit_io_write: 0x313678, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313778, value : 32'h286}, //phyinit_io_write: 0x313679, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313779, value : 32'h286}, //phyinit_io_write: 0x313778, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313878, value : 32'h286}, //phyinit_io_write: 0x313779, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h313879, value : 32'h286}, //phyinit_io_write: 0x313878, 0x286
                          '{ step_type : REG_WRITE, reg_addr : 32'h310020, value : 32'h1e6}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming RxEnDlyTg0/Tg1 to 0x1e6
                          '{ step_type : REG_WRITE, reg_addr : 32'h310021, value : 32'h1e6}, //phyinit_io_write: 0x310020, 0x1e6
                          '{ step_type : REG_WRITE, reg_addr : 32'h311020, value : 32'h1e6}, //phyinit_io_write: 0x310021, 0x1e6
                          '{ step_type : REG_WRITE, reg_addr : 32'h311021, value : 32'h1e6}, //phyinit_io_write: 0x311020, 0x1e6
                          '{ step_type : REG_WRITE, reg_addr : 32'h312020, value : 32'h1e6}, //phyinit_io_write: 0x311021, 0x1e6
                          '{ step_type : REG_WRITE, reg_addr : 32'h312021, value : 32'h1e6}, //phyinit_io_write: 0x312020, 0x1e6
                          '{ step_type : REG_WRITE, reg_addr : 32'h313020, value : 32'h1e6}, //phyinit_io_write: 0x312021, 0x1e6
                          '{ step_type : REG_WRITE, reg_addr : 32'h313021, value : 32'h1e6}, //phyinit_io_write: 0x313020, 0x1e6
                          '{ step_type : REG_WRITE, reg_addr : 32'h310010, value : 32'h202}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming RxClkT2UIDlyTg0/Tg1 and RxClkC2UIDlyTg0/Tg1 to 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310011, value : 32'h202}, //phyinit_io_write: 0x310010, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310012, value : 32'h202}, //phyinit_io_write: 0x310011, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310013, value : 32'h202}, //phyinit_io_write: 0x310012, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310110, value : 32'h202}, //phyinit_io_write: 0x310013, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310111, value : 32'h202}, //phyinit_io_write: 0x310110, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310112, value : 32'h202}, //phyinit_io_write: 0x310111, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310113, value : 32'h202}, //phyinit_io_write: 0x310112, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310210, value : 32'h202}, //phyinit_io_write: 0x310113, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310211, value : 32'h202}, //phyinit_io_write: 0x310210, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310212, value : 32'h202}, //phyinit_io_write: 0x310211, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310213, value : 32'h202}, //phyinit_io_write: 0x310212, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310310, value : 32'h202}, //phyinit_io_write: 0x310213, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310311, value : 32'h202}, //phyinit_io_write: 0x310310, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310312, value : 32'h202}, //phyinit_io_write: 0x310311, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310313, value : 32'h202}, //phyinit_io_write: 0x310312, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310410, value : 32'h202}, //phyinit_io_write: 0x310313, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310411, value : 32'h202}, //phyinit_io_write: 0x310410, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310412, value : 32'h202}, //phyinit_io_write: 0x310411, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310413, value : 32'h202}, //phyinit_io_write: 0x310412, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310510, value : 32'h202}, //phyinit_io_write: 0x310413, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310511, value : 32'h202}, //phyinit_io_write: 0x310510, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310512, value : 32'h202}, //phyinit_io_write: 0x310511, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310513, value : 32'h202}, //phyinit_io_write: 0x310512, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310610, value : 32'h202}, //phyinit_io_write: 0x310513, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310611, value : 32'h202}, //phyinit_io_write: 0x310610, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310612, value : 32'h202}, //phyinit_io_write: 0x310611, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310613, value : 32'h202}, //phyinit_io_write: 0x310612, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310710, value : 32'h202}, //phyinit_io_write: 0x310613, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310711, value : 32'h202}, //phyinit_io_write: 0x310710, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310712, value : 32'h202}, //phyinit_io_write: 0x310711, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310713, value : 32'h202}, //phyinit_io_write: 0x310712, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310810, value : 32'h202}, //phyinit_io_write: 0x310713, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310811, value : 32'h202}, //phyinit_io_write: 0x310810, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310812, value : 32'h202}, //phyinit_io_write: 0x310811, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h310813, value : 32'h202}, //phyinit_io_write: 0x310812, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311010, value : 32'h202}, //phyinit_io_write: 0x310813, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311011, value : 32'h202}, //phyinit_io_write: 0x311010, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311012, value : 32'h202}, //phyinit_io_write: 0x311011, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311013, value : 32'h202}, //phyinit_io_write: 0x311012, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311110, value : 32'h202}, //phyinit_io_write: 0x311013, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311111, value : 32'h202}, //phyinit_io_write: 0x311110, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311112, value : 32'h202}, //phyinit_io_write: 0x311111, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311113, value : 32'h202}, //phyinit_io_write: 0x311112, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311210, value : 32'h202}, //phyinit_io_write: 0x311113, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311211, value : 32'h202}, //phyinit_io_write: 0x311210, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311212, value : 32'h202}, //phyinit_io_write: 0x311211, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311213, value : 32'h202}, //phyinit_io_write: 0x311212, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311310, value : 32'h202}, //phyinit_io_write: 0x311213, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311311, value : 32'h202}, //phyinit_io_write: 0x311310, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311312, value : 32'h202}, //phyinit_io_write: 0x311311, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311313, value : 32'h202}, //phyinit_io_write: 0x311312, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311410, value : 32'h202}, //phyinit_io_write: 0x311313, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311411, value : 32'h202}, //phyinit_io_write: 0x311410, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311412, value : 32'h202}, //phyinit_io_write: 0x311411, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311413, value : 32'h202}, //phyinit_io_write: 0x311412, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311510, value : 32'h202}, //phyinit_io_write: 0x311413, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311511, value : 32'h202}, //phyinit_io_write: 0x311510, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311512, value : 32'h202}, //phyinit_io_write: 0x311511, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311513, value : 32'h202}, //phyinit_io_write: 0x311512, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311610, value : 32'h202}, //phyinit_io_write: 0x311513, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311611, value : 32'h202}, //phyinit_io_write: 0x311610, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311612, value : 32'h202}, //phyinit_io_write: 0x311611, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311613, value : 32'h202}, //phyinit_io_write: 0x311612, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311710, value : 32'h202}, //phyinit_io_write: 0x311613, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311711, value : 32'h202}, //phyinit_io_write: 0x311710, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311712, value : 32'h202}, //phyinit_io_write: 0x311711, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311713, value : 32'h202}, //phyinit_io_write: 0x311712, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311810, value : 32'h202}, //phyinit_io_write: 0x311713, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311811, value : 32'h202}, //phyinit_io_write: 0x311810, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311812, value : 32'h202}, //phyinit_io_write: 0x311811, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h311813, value : 32'h202}, //phyinit_io_write: 0x311812, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312010, value : 32'h202}, //phyinit_io_write: 0x311813, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312011, value : 32'h202}, //phyinit_io_write: 0x312010, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312012, value : 32'h202}, //phyinit_io_write: 0x312011, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312013, value : 32'h202}, //phyinit_io_write: 0x312012, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312110, value : 32'h202}, //phyinit_io_write: 0x312013, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312111, value : 32'h202}, //phyinit_io_write: 0x312110, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312112, value : 32'h202}, //phyinit_io_write: 0x312111, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312113, value : 32'h202}, //phyinit_io_write: 0x312112, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312210, value : 32'h202}, //phyinit_io_write: 0x312113, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312211, value : 32'h202}, //phyinit_io_write: 0x312210, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312212, value : 32'h202}, //phyinit_io_write: 0x312211, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312213, value : 32'h202}, //phyinit_io_write: 0x312212, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312310, value : 32'h202}, //phyinit_io_write: 0x312213, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312311, value : 32'h202}, //phyinit_io_write: 0x312310, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312312, value : 32'h202}, //phyinit_io_write: 0x312311, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312313, value : 32'h202}, //phyinit_io_write: 0x312312, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312410, value : 32'h202}, //phyinit_io_write: 0x312313, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312411, value : 32'h202}, //phyinit_io_write: 0x312410, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312412, value : 32'h202}, //phyinit_io_write: 0x312411, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312413, value : 32'h202}, //phyinit_io_write: 0x312412, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312510, value : 32'h202}, //phyinit_io_write: 0x312413, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312511, value : 32'h202}, //phyinit_io_write: 0x312510, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312512, value : 32'h202}, //phyinit_io_write: 0x312511, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312513, value : 32'h202}, //phyinit_io_write: 0x312512, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312610, value : 32'h202}, //phyinit_io_write: 0x312513, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312611, value : 32'h202}, //phyinit_io_write: 0x312610, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312612, value : 32'h202}, //phyinit_io_write: 0x312611, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312613, value : 32'h202}, //phyinit_io_write: 0x312612, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312710, value : 32'h202}, //phyinit_io_write: 0x312613, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312711, value : 32'h202}, //phyinit_io_write: 0x312710, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312712, value : 32'h202}, //phyinit_io_write: 0x312711, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312713, value : 32'h202}, //phyinit_io_write: 0x312712, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312810, value : 32'h202}, //phyinit_io_write: 0x312713, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312811, value : 32'h202}, //phyinit_io_write: 0x312810, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312812, value : 32'h202}, //phyinit_io_write: 0x312811, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h312813, value : 32'h202}, //phyinit_io_write: 0x312812, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313010, value : 32'h202}, //phyinit_io_write: 0x312813, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313011, value : 32'h202}, //phyinit_io_write: 0x313010, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313012, value : 32'h202}, //phyinit_io_write: 0x313011, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313013, value : 32'h202}, //phyinit_io_write: 0x313012, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313110, value : 32'h202}, //phyinit_io_write: 0x313013, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313111, value : 32'h202}, //phyinit_io_write: 0x313110, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313112, value : 32'h202}, //phyinit_io_write: 0x313111, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313113, value : 32'h202}, //phyinit_io_write: 0x313112, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313210, value : 32'h202}, //phyinit_io_write: 0x313113, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313211, value : 32'h202}, //phyinit_io_write: 0x313210, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313212, value : 32'h202}, //phyinit_io_write: 0x313211, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313213, value : 32'h202}, //phyinit_io_write: 0x313212, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313310, value : 32'h202}, //phyinit_io_write: 0x313213, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313311, value : 32'h202}, //phyinit_io_write: 0x313310, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313312, value : 32'h202}, //phyinit_io_write: 0x313311, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313313, value : 32'h202}, //phyinit_io_write: 0x313312, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313410, value : 32'h202}, //phyinit_io_write: 0x313313, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313411, value : 32'h202}, //phyinit_io_write: 0x313410, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313412, value : 32'h202}, //phyinit_io_write: 0x313411, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313413, value : 32'h202}, //phyinit_io_write: 0x313412, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313510, value : 32'h202}, //phyinit_io_write: 0x313413, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313511, value : 32'h202}, //phyinit_io_write: 0x313510, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313512, value : 32'h202}, //phyinit_io_write: 0x313511, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313513, value : 32'h202}, //phyinit_io_write: 0x313512, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313610, value : 32'h202}, //phyinit_io_write: 0x313513, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313611, value : 32'h202}, //phyinit_io_write: 0x313610, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313612, value : 32'h202}, //phyinit_io_write: 0x313611, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313613, value : 32'h202}, //phyinit_io_write: 0x313612, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313710, value : 32'h202}, //phyinit_io_write: 0x313613, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313711, value : 32'h202}, //phyinit_io_write: 0x313710, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313712, value : 32'h202}, //phyinit_io_write: 0x313711, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313713, value : 32'h202}, //phyinit_io_write: 0x313712, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313810, value : 32'h202}, //phyinit_io_write: 0x313713, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313811, value : 32'h202}, //phyinit_io_write: 0x313810, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313812, value : 32'h202}, //phyinit_io_write: 0x313811, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h313813, value : 32'h202}, //phyinit_io_write: 0x313812, 0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h31000c, value : 32'h34}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming PptWck2DqoCntInvTrn1 to 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h31000d, value : 32'h34}, //phyinit_io_write: 0x31000c, 0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h310014, value : 32'h67}, //phyinit_io_write: 0x31000d, 0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h310015, value : 32'h67}, //phyinit_io_write: 0x310014, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h31100c, value : 32'h34}, //phyinit_io_write: 0x310015, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h31100d, value : 32'h34}, //phyinit_io_write: 0x31100c, 0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h311014, value : 32'h67}, //phyinit_io_write: 0x31100d, 0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h311015, value : 32'h67}, //phyinit_io_write: 0x311014, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h31200c, value : 32'h34}, //phyinit_io_write: 0x311015, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h31200d, value : 32'h34}, //phyinit_io_write: 0x31200c, 0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h312014, value : 32'h67}, //phyinit_io_write: 0x31200d, 0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h312015, value : 32'h67}, //phyinit_io_write: 0x312014, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h31300c, value : 32'h34}, //phyinit_io_write: 0x312015, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h31300d, value : 32'h34}, //phyinit_io_write: 0x31300c, 0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h313014, value : 32'h67}, //phyinit_io_write: 0x31300d, 0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h313015, value : 32'h67}, //phyinit_io_write: 0x313014, 0x67
                          '{ step_type : REG_WRITE, reg_addr : 32'h70077, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming HwtCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h320071, value : 32'h44}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming HMRxReplicaLcdlSeed HMRxSeed to 0xd0 HMRxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h300063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC0 Instance0 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h301063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC1 Instance1 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h302063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC2 Instance2 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h303063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC3 Instance3 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h304063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC4 Instance4 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h305063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX0 HMAC5 Instance5 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h307063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC0 Instance7 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h308063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC1 Instance8 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h309063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC2 Instance9 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h30a063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC3 Instance10 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h30b063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC4 Instance11 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h30c063, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=3, Memclk=200MHz, Programming ACX1 HMAC5 Instance12 HMTxLcdlSeed HMTxSeed to 0xd0 HMTxSeedIs1UI 0x1 
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e0063, value : 32'h2d0}, //phyinit_io_write: 0x30c063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e0064, value : 32'h2d0}, //phyinit_io_write: 0x3e0063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e0087, value : 32'h2d0}, //phyinit_io_write: 0x3e0064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e1063, value : 32'h2d0}, //phyinit_io_write: 0x3e0087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e1064, value : 32'h2d0}, //phyinit_io_write: 0x3e1063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e1087, value : 32'h2d0}, //phyinit_io_write: 0x3e1064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e2063, value : 32'h2d0}, //phyinit_io_write: 0x3e1087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e2064, value : 32'h2d0}, //phyinit_io_write: 0x3e2063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e2087, value : 32'h2d0}, //phyinit_io_write: 0x3e2064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e3063, value : 32'h2d0}, //phyinit_io_write: 0x3e2087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e3064, value : 32'h2d0}, //phyinit_io_write: 0x3e3063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e3087, value : 32'h2d0}, //phyinit_io_write: 0x3e3064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e4063, value : 32'h2d0}, //phyinit_io_write: 0x3e3087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e4064, value : 32'h2d0}, //phyinit_io_write: 0x3e4063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e4087, value : 32'h2d0}, //phyinit_io_write: 0x3e4064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e5063, value : 32'h2d0}, //phyinit_io_write: 0x3e4087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e5064, value : 32'h2d0}, //phyinit_io_write: 0x3e5063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e5087, value : 32'h2d0}, //phyinit_io_write: 0x3e5064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e6063, value : 32'h2d0}, //phyinit_io_write: 0x3e5087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e6064, value : 32'h2d0}, //phyinit_io_write: 0x3e6063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e6087, value : 32'h2d0}, //phyinit_io_write: 0x3e6064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e7063, value : 32'h2d0}, //phyinit_io_write: 0x3e6087, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e7064, value : 32'h2d0}, //phyinit_io_write: 0x3e7063, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e7087, value : 32'h2d0}, //phyinit_io_write: 0x3e7064, 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h39080a, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=3 Programming Seq0bGPR10 to mission mode HMTxLcdlSeed value 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h39080b, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=3 Programming Seq0bGPR11 to mission mode HMTxLcdlSeed value 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h390815, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=3 Programming Seq0bGPR21 to mission mode HMTxLcdlSeed value 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h390816, value : 32'h2d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=3 Programming Seq0bGPR22 to mission mode HMTxLcdlSeed value 0x2d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31015f, value : 32'h14d0}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=3, Memclk=200MHz, Programming RDqRDqsCntrl to 0x14d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31115f, value : 32'h14d0}, //phyinit_io_write: 0x31015f, 0x14d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31215f, value : 32'h14d0}, //phyinit_io_write: 0x31115f, 0x14d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31315f, value : 32'h14d0}, //phyinit_io_write: 0x31215f, 0x14d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h360009, value : 32'h10}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Memclk=200MHz, Programming CPllDacValIn to 0x10
                          '{ step_type : REG_WRITE, reg_addr : 32'h3102a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE0.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3102a1, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE0.RxReplicaPathPhase1 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h3102a2, value : 32'h142}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE0.RxReplicaPathPhase2 to 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h3102a3, value : 32'h1ff}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE0.RxReplicaPathPhase3 to 0x1ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h3102a4, value : 32'h1ff}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE0.RxReplicaPathPhase4 to 0x1ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h3112a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE1.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3112a1, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE1.RxReplicaPathPhase1 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h3112a2, value : 32'h142}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE1.RxReplicaPathPhase2 to 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h3112a3, value : 32'h1ff}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE1.RxReplicaPathPhase3 to 0x1ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h3112a4, value : 32'h1ff}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE1.RxReplicaPathPhase4 to 0x1ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h3122a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE2.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3122a1, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE2.RxReplicaPathPhase1 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h3122a2, value : 32'h142}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE2.RxReplicaPathPhase2 to 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h3122a3, value : 32'h1ff}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE2.RxReplicaPathPhase3 to 0x1ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h3122a4, value : 32'h1ff}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE2.RxReplicaPathPhase4 to 0x1ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h3132a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE3.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3132a1, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE3.RxReplicaPathPhase1 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h3132a2, value : 32'h142}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE3.RxReplicaPathPhase2 to 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h3132a3, value : 32'h1ff}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE3.RxReplicaPathPhase3 to 0x1ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h3132a4, value : 32'h1ff}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE3.RxReplicaPathPhase4 to 0x1ff
                          '{ step_type : REG_WRITE, reg_addr : 32'h3102ad, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE0.RxReplicaCtl01::RxReplicaSelPathPhase to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3112ad, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE1.RxReplicaCtl01::RxReplicaSelPathPhase to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3122ad, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE2.RxReplicaCtl01::RxReplicaSelPathPhase to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3132ad, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE3.RxReplicaCtl01::RxReplicaSelPathPhase to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h3102af, value : 32'h23}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE0.RxReplicaCtl03 to 0x23
                          '{ step_type : REG_WRITE, reg_addr : 32'h3112af, value : 32'h23}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE1.RxReplicaCtl03 to 0x23
                          '{ step_type : REG_WRITE, reg_addr : 32'h3122af, value : 32'h23}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE2.RxReplicaCtl03 to 0x23
                          '{ step_type : REG_WRITE, reg_addr : 32'h3132af, value : 32'h23}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming DBYTE3.RxReplicaCtl03 to 0x23
                          '{ step_type : REG_WRITE, reg_addr : 32'h390807, value : 32'h9701}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming Seq0BGPR7 to save ZQCalCodeOvrValPU=0x12e and ZQCalCodeOvrEnPU=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h390808, value : 32'hb681}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=3, Programming Seq0BGPR8 to save ZQCalCodeOvrValPD=0x16d and ZQCalCodeOvrEnPD=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
//[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] End of dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop(), PState=3
// [dwc_ddrphy_phyinit_userCustom_E_setDfiClk] Start of dwc_ddrphy_phyinit_userCustom_E_setDfiClk()
// [dwc_ddrphy_phyinit_userCustom_E_setDfiClk] End of dwc_ddrphy_phyinit_userCustom_E_setDfiClk()
// [dwc_ddrphy_phyinit_F_loadDMEM1D] Start of dwc_ddrphy_phyinit_F_loadDMEM (pstate=3, Train2D=0)
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0088, value : 32'h1}, //[dwc_ddrphy_phyinit_F_loadDMEM] Program csr StartDccmClear to 1 to clear DCCM.
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 8300},
//Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 8300 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0088, value : 32'h0}, //[dwc_ddrphy_phyinit_F_loadDMEM] Program csr StartDccmClear to 0 after DCCM clear is done.
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}, //Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 40 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'h58000, value : 32'h600}, // [dwc_ddrphy_phyinit_WriteOutMem] STARTING. offset 0x58000 size 0x6000, sparse_write=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h58001, value : 32'h6400003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58002, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58004, value : 32'hff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58005, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58009, value : 32'h310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5800f, value : 32'h10000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58010, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58016, value : 32'h20200000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58017, value : 32'h22222020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58018, value : 32'he0e2222},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58019, value : 32'h54540e0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801a, value : 32'h44445454},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801b, value : 32'h50504444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801c, value : 32'h5050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801d, value : 32'h50500000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801e, value : 32'h50505050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801f, value : 32'h5050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58020, value : 32'hac840000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58021, value : 32'hac84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58023, value : 32'h2020000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58024, value : 32'h202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5802a, value : 32'h4040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5802b, value : 32'h404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58032, value : 32'h60600000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58033, value : 32'h6060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58048, value : 32'hf000001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58049, value : 32'hf},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58054, value : 32'h5c0032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58055, value : 32'he000b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58056, value : 32'h164013a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58057, value : 32'h1e801be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58062, value : 32'h6400c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58103, value : 32'h50b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58104, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58108, value : 32'h8080808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58110, value : 32'hef0f4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811b, value : 32'h4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811d, value : 32'h40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811e, value : 32'h180f0e0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811f, value : 32'h4746451e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58120, value : 32'h4a4948},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58121, value : 32'h1000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58125, value : 32'h40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58126, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58129, value : 32'hffffffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5812e, value : 32'h2f059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5812f, value : 32'hffb50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58130, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58131, value : 32'h1f0b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58132, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58133, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58134, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58135, value : 32'hf0b00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58136, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58137, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58138, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58139, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813a, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813b, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813c, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813d, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813e, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813f, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58140, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58141, value : 32'hff740182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58142, value : 32'h800001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58143, value : 32'h1ffbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58144, value : 32'hf0be0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58145, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58146, value : 32'h1f0a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58147, value : 32'hf0a20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58148, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58149, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814a, value : 32'h40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814b, value : 32'h308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814c, value : 32'h560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814e, value : 32'h80000dbc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814f, value : 32'h309},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58150, value : 32'h561},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58151, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58152, value : 32'h80000dcd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58153, value : 32'he0305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58154, value : 32'he0205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58155, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58156, value : 32'h80000dde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58157, value : 32'he0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58158, value : 32'he0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58159, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815a, value : 32'h80000e44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815b, value : 32'he0301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815c, value : 32'he0201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815d, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815e, value : 32'h80000e57},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815f, value : 32'he0302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58160, value : 32'he0202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58161, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58162, value : 32'h80000e6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58163, value : 32'he0303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58164, value : 32'he0203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58165, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58166, value : 32'h80000e7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58167, value : 32'he0304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58168, value : 32'he0204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58169, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816a, value : 32'h80000e90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816b, value : 32'h1ff01ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816c, value : 32'he0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816e, value : 32'h63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816f, value : 32'h64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58170, value : 32'h660},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58172, value : 32'h80000d8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58173, value : 32'h661},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58174, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58175, value : 32'h80000dad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58176, value : 32'he00f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58177, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58178, value : 32'h80000def},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58179, value : 32'he00f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817a, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817b, value : 32'h80000e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817c, value : 32'he00f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817d, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817e, value : 32'h80000e11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817f, value : 32'he00f3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58180, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58181, value : 32'h80000e22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58182, value : 32'he00f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58183, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58184, value : 32'h80000e33},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58185, value : 32'he00f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58186, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58187, value : 32'h80000d9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58188, value : 32'h2011210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58189, value : 32'h1c0a1403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818a, value : 32'hb112e29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818b, value : 32'h1916150d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818c, value : 32'h180f0e0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818d, value : 32'h453a131e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818e, value : 32'h49484746},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818f, value : 32'h2006e4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58190, value : 32'h100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58191, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58192, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58194, value : 32'h2150001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58195, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58196, value : 32'h1010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58197, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58198, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58199, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819a, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819b, value : 32'h6400002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819c, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819d, value : 32'h30215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819e, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819f, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a0, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a1, value : 32'h10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a2, value : 32'habe0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a3, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a4, value : 32'h50320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a5, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c5, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c6, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c7, value : 32'h43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c8, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c9, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ca, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cb, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cc, value : 32'h42b0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cd, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ce, value : 32'h200c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cf, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d0, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d1, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d2, value : 32'h10003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d3, value : 32'h8550002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d4, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d5, value : 32'h40158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d6, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d7, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d8, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d9, value : 32'h10005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581da, value : 32'hc800002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581db, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581dc, value : 32'h601d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581dd, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581de, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581df, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e0, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e1, value : 32'h10ab0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e2, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e3, value : 32'h80258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e4, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e5, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e6, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e7, value : 32'h20009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e8, value : 32'h157c0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e9, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ea, value : 32'ha02ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581eb, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ec, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ed, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ee, value : 32'h2000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ef, value : 32'h19000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f0, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f1, value : 32'hc03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f2, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f3, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f4, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f5, value : 32'h3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f6, value : 32'h21550006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f7, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f8, value : 32'he04b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f9, value : 32'h70003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fa, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fb, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fc, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fd, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fe, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ff, value : 32'h2150004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58200, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58201, value : 32'h4010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58202, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58203, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58204, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58205, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58206, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58207, value : 32'h80006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58208, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58209, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820a, value : 32'h6400006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820b, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820c, value : 32'h80215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820d, value : 32'h2000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820e, value : 32'h30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820f, value : 32'h70004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58210, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58211, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58212, value : 32'he0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58213, value : 32'h70001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58214, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58215, value : 32'habe0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58216, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58217, value : 32'ha0320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58218, value : 32'h30010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58219, value : 32'h40009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5821a, value : 32'h80004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824c, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824d, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824e, value : 32'h20043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824f, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58250, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58251, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58252, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58253, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58254, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58255, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58256, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58257, value : 32'h42b0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58258, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58259, value : 32'h300c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825a, value : 32'h10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825b, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825c, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825d, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825e, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825f, value : 32'h50004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58260, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58261, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58262, value : 32'h8550004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58263, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58264, value : 32'h40158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58265, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58266, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58267, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58268, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58269, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826a, value : 32'h80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826b, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826c, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826d, value : 32'hc800004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826e, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826f, value : 32'h601d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58270, value : 32'h20009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58271, value : 32'h30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58272, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58273, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58274, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58275, value : 32'hb0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58276, value : 32'h70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58277, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58278, value : 32'h10ab0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58279, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827a, value : 32'h70258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827b, value : 32'h3000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827c, value : 32'h30008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827d, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827e, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827f, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58280, value : 32'he0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58281, value : 32'h90003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58282, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58283, value : 32'h157c0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58284, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58285, value : 32'h902ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58286, value : 32'h4000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58287, value : 32'h4000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58288, value : 32'h60002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58289, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828a, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828b, value : 32'h100009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828c, value : 32'hb0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828d, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828e, value : 32'h19000006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828f, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58290, value : 32'hb03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58291, value : 32'h50013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58292, value : 32'h5000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58293, value : 32'h70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58294, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58295, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58296, value : 32'h16000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58297, value : 32'hf0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58298, value : 32'h20006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58299, value : 32'h21550008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829a, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829b, value : 32'he04b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829c, value : 32'h60018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829d, value : 32'h70010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829e, value : 32'h90002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829f, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a0, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a1, value : 32'h60006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a2, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a4, value : 32'h60001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a5, value : 32'h2150007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a6, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a7, value : 32'h8010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a8, value : 32'h80008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582aa, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ab, value : 32'h90007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ac, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ad, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ae, value : 32'ha000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582af, value : 32'h1000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b0, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b1, value : 32'h80002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b2, value : 32'h640000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b3, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b4, value : 32'hc0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b5, value : 32'he000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b6, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b7, value : 32'h30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b8, value : 32'hb0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b9, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ba, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bb, value : 32'h100010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bc, value : 32'h30012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bd, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582be, value : 32'ha0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bf, value : 32'habe000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c0, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c1, value : 32'h120320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c2, value : 32'h140014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c3, value : 32'h70005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c4, value : 32'h40007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c5, value : 32'he000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58300, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58301, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58302, value : 32'h30043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58303, value : 32'h30003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58305, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58306, value : 32'h40003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58307, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58308, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58309, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830a, value : 32'h4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830c, value : 32'h40001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830d, value : 32'h42b0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830e, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830f, value : 32'h500c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58310, value : 32'h50005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58311, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58312, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58313, value : 32'h50004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58314, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58315, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58316, value : 32'h70006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58317, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58318, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58319, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831a, value : 32'h8550006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831b, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831c, value : 32'h80158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831d, value : 32'h90008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831e, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831f, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58320, value : 32'h70005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58321, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58322, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58323, value : 32'ha0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58324, value : 32'h3000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58325, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58326, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58327, value : 32'hc800007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58328, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58329, value : 32'ha01d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832a, value : 32'hc000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832b, value : 32'h40003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832c, value : 32'h30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832d, value : 32'h80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832e, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832f, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58330, value : 32'hd000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58331, value : 32'h4000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58332, value : 32'h60005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58333, value : 32'h60003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58334, value : 32'h10ab0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58335, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58336, value : 32'hd0258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58337, value : 32'hf000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58338, value : 32'h60005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58339, value : 32'h30007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833a, value : 32'h90006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833b, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833c, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833d, value : 32'h10000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833e, value : 32'h60011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833f, value : 32'h80007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58340, value : 32'h60004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58341, value : 32'h157c000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58342, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58343, value : 32'h1002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58344, value : 32'h130011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58345, value : 32'h70006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58346, value : 32'h40009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58347, value : 32'hb0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58348, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58349, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834a, value : 32'h120011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834b, value : 32'h70014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834c, value : 32'ha0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834d, value : 32'h70004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834e, value : 32'h1900000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834f, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58350, value : 32'h1403aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58351, value : 32'h180016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58352, value : 32'h90007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58353, value : 32'h5000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58354, value : 32'he0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58355, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58356, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58357, value : 32'h190017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58358, value : 32'h8001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58359, value : 32'hb000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835a, value : 32'ha0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835b, value : 32'h21550010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835c, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835d, value : 32'h1904b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835e, value : 32'h1d001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835f, value : 32'hb0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58360, value : 32'h7000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58361, value : 32'h12000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58362, value : 32'ha05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58363, value : 32'h50000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58364, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58365, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58366, value : 32'h43416564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58367, value : 32'h63500030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58368, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58369, value : 32'h646f4341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836a, value : 32'h53514465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836b, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836c, value : 32'h4143446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836d, value : 32'h65646f43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836e, value : 32'h314341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836f, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58370, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58371, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58372, value : 32'h30434174},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58373, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58374, value : 32'h4443446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58375, value : 32'h7366664f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58376, value : 32'h43417465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58377, value : 32'h63500031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58378, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58379, value : 32'h66664f44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837a, value : 32'h44746573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837b, value : 32'h50005351},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837c, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837d, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837e, value : 32'h71446564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837f, value : 32'h306e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58380, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58381, value : 32'h43414344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58382, value : 32'h4465646f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58383, value : 32'h316e4c71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58384, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58385, value : 32'h4143446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58386, value : 32'h65646f43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58387, value : 32'h6e4c7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58388, value : 32'h63500032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58389, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838a, value : 32'h646f4341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838b, value : 32'h4c714465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838c, value : 32'h5000336e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838d, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838e, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838f, value : 32'h71446564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58390, value : 32'h346e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58391, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58392, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58393, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58394, value : 32'h4c714474},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58395, value : 32'h5000306e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58396, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58397, value : 32'h664f4443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58398, value : 32'h74657366},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58399, value : 32'h6e4c7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839a, value : 32'h63500031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839b, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839c, value : 32'h66664f44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839d, value : 32'h44746573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839e, value : 32'h326e4c71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839f, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a0, value : 32'h4443446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a1, value : 32'h7366664f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a2, value : 32'h71447465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a3, value : 32'h336e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a4, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a5, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a6, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a7, value : 32'h4c714474},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a8, value : 32'h346e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a9, value : 32'h4050607},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583aa, value : 32'h10203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ab, value : 32'hc0b0a09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ac, value : 32'hb50f0e0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ad, value : 32'h1ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ae, value : 32'h1f0b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583af, value : 32'hb3000100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b0, value : 32'h1f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b1, value : 32'h1f0b400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b2, value : 32'hb0000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b3, value : 32'h300001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b4, value : 32'h7f00300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b5, value : 32'h4000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b6, value : 32'h7f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b7, value : 32'h1fe0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b8, value : 32'h4000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b9, value : 32'h1fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ba, value : 32'h7f01100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bb, value : 32'h21000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bc, value : 32'h1fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bd, value : 32'h1ffbe00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583be, value : 32'hbe000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bf, value : 32'h10001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c0, value : 32'h1f0a700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c1, value : 32'ha2000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c2, value : 32'h20001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c3, value : 32'h2007900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c4, value : 32'h4000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c5, value : 32'h1008b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c6, value : 32'hf05f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c7, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c8, value : 32'h1ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c9, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ca, value : 32'h1ff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cb, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cc, value : 32'hf0b001ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cd, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ce, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cf, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d0, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d1, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d2, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d3, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d4, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d5, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d6, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d7, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d8, value : 32'hf0a70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d9, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583da, value : 32'he000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583db, value : 32'hc000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583dc, value : 32'ha000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583dd, value : 32'h80009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583de, value : 32'h60007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583df, value : 32'h40005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e0, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e1, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e2, value : 32'h110010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e3, value : 32'h130012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e4, value : 32'h150014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e5, value : 32'h170016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e6, value : 32'h190018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e7, value : 32'h1b001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e8, value : 32'h1d001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e9, value : 32'h1f001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ea, value : 32'hef77dbb7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583eb, value : 32'hfbdff7bd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ec, value : 32'hbddfb76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ed, value : 32'hbdffbdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ee, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ef, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f0, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f1, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f2, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f3, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f4, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f5, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f6, value : 32'h1ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f7, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f8, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f9, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fa, value : 32'hf0b90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fb, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fc, value : 32'h1f0ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fd, value : 32'hf0b10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fe, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ff, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58400, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58401, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58402, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58403, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58404, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58405, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58406, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58407, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58408, value : 32'h7f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58409, value : 32'hfe200002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840a, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840b, value : 32'h7f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840c, value : 32'hf01cffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840d, value : 32'hffff0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840e, value : 32'h1fe2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840f, value : 32'hfe2bffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58410, value : 32'hffff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58411, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58412, value : 32'hffb50040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58413, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58414, value : 32'h1f0b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58415, value : 32'hf0b40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58416, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58417, value : 32'h1f0b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58418, value : 32'hf0ba0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58419, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841a, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841b, value : 32'hf0b00002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841c, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841d, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841e, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841f, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58420, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58421, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58422, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58423, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58424, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58425, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58426, value : 32'h7f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58427, value : 32'hfe200002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58428, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58429, value : 32'h7f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842a, value : 32'hf01cffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842b, value : 32'hffff0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842c, value : 32'h1fe2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842d, value : 32'hfe2bffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842e, value : 32'hffff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842f, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58430, value : 32'h40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58431, value : 32'h8840884},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58432, value : 32'h20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58433, value : 32'h10010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58434, value : 32'h10012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58435, value : 32'h1007a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58436, value : 32'h10028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58437, value : 32'h60000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58438, value : 32'h50005000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58439, value : 32'h2008050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843b, value : 32'h60080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843c, value : 32'h3c5a5555},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843d, value : 32'h600000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58440, value : 32'h70},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58441, value : 32'h75},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58442, value : 32'h26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58443, value : 32'ha0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58444, value : 32'ha1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58445, value : 32'ha4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58446, value : 32'ha5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58447, value : 32'ha030201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58448, value : 32'he0d0c0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58449, value : 32'h1413120f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844a, value : 32'h18171615},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844b, value : 32'h1e1c1a19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844c, value : 32'h2221201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844d, value : 32'h2e292825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844e, value : 32'h4746453a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844f, value : 32'h4a4948},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1}, //This allows the firmware unrestricted access to the configuration CSRs.
//[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
// [dwc_ddrphy_phyinit_F_loadDMEM1D] End of dwc_ddrphy_phyinit_F_loadDMEM, Pstate=3
// [dwc_ddrphy_phyinit_G_execFW] Start of dwc_ddrphy_phyinit_G_execFW
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1}, ////     Then rewrite the CSR so that only the StallToMicro remains set (all other fields should be zero).
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h9}, //[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h0}, // [dwc_ddrphy_phyinit_userCustom_G_waitFwDone] Start of dwc_ddrphy_phyinit_userCustom_G_waitFwDone()
// [dwc_ddrphy_phyinit_userCustom_G_waitFwDone] End of dwc_ddrphy_phyinit_userCustom_G_waitFwDone()
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h1}, //// 4.   Halt the microcontroller."
// [dwc_ddrphy_phyinit_G_execFW] End of dwc_ddrphy_phyinit_G_execFW
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}, // [dwc_ddrphy_phyinit_userCustom_H_readMsgBlock] Start of dwc_ddrphy_phyinit_userCustom_H_readMsgBlock()
// [dwc_ddrphy_phyinit_userCustom_H_readMsgBlock] End of dwc_ddrphy_phyinit_userCustom_H_readMsgBlock ()
// 3. If training is required at another frequency, repeat the operations starting at step (E).
// [dwc_ddrphy_phyinit_H_readMsgBlock] End of dwc_ddrphy_phyinit_H_readMsgBlock
//[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Start of dwc_ddrphy_phyinit_I_loadPIEImagePsLoop(), PState=3
                          '{ step_type : REG_WRITE, reg_addr : 32'h360008, value : 32'h4822}, //[dwc_ddrphy_phyinit_programPLL] [phyinit_I_loadPIEImagePsLoop] Pstate=3,  Memclk=200MHz, Programming CpllCtrl5 to 0x4822.
                          '{ step_type : REG_WRITE, reg_addr : 32'h60006, value : 32'h3f0}, //End of dwc_ddrphy_phyinit_programPLL(), PState=3
                          '{ step_type : REG_WRITE, reg_addr : 32'h330015, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h331015, value : 32'h0}, //phyinit_io_write: 0x330015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31007c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31107c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31207c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31307c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31007c, value : 32'h0}, //phyinit_io_write: 0x31307c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31107c, value : 32'h0}, //phyinit_io_write: 0x31007c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31207c, value : 32'h0}, //phyinit_io_write: 0x31107c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31307c, value : 32'h0}, //phyinit_io_write: 0x31207c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h330015, value : 32'h0}, //phyinit_io_write: 0x31307c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h331015, value : 32'h0}, //phyinit_io_write: 0x330015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h370141, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming ACSMWckFreeRunMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h39080c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming GPR12 with Zcalkclkdiv to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h310027, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming RxClkCntl1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h311027, value : 32'h0}, //phyinit_io_write: 0x310027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h312027, value : 32'h0}, //phyinit_io_write: 0x311027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h313027, value : 32'h0}, //phyinit_io_write: 0x312027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31020f, value : 32'h8}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=3, Programming RxReplicaCtl04 to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h31120f, value : 32'h8}, //phyinit_io_write: 0x31020f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h31220f, value : 32'h8}, //phyinit_io_write: 0x31120f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h31320f, value : 32'h8}, //phyinit_io_write: 0x31220f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e003f, value : 32'h0}, //phyinit_io_write: 0x31320f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e008d, value : 32'h0}, //phyinit_io_write: 0x3e003f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e103f, value : 32'h0}, //phyinit_io_write: 0x3e008d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e108d, value : 32'h0}, //phyinit_io_write: 0x3e103f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e203f, value : 32'h0}, //phyinit_io_write: 0x3e108d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e208d, value : 32'h0}, //phyinit_io_write: 0x3e203f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e303f, value : 32'h0}, //phyinit_io_write: 0x3e208d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e308d, value : 32'h0}, //phyinit_io_write: 0x3e303f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e403f, value : 32'h0}, //phyinit_io_write: 0x3e308d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e408d, value : 32'h0}, //phyinit_io_write: 0x3e403f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e503f, value : 32'h0}, //phyinit_io_write: 0x3e408d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e508d, value : 32'h0}, //phyinit_io_write: 0x3e503f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e603f, value : 32'h0}, //phyinit_io_write: 0x3e508d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e608d, value : 32'h0}, //phyinit_io_write: 0x3e603f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e703f, value : 32'h0}, //phyinit_io_write: 0x3e608d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h3e708d, value : 32'h0}, //phyinit_io_write: 0x3e703f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h390903, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] PState=3, Programming RtrnMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70072, value : 32'h3}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming HwtLpCsEnA to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h39080e, value : 32'h3}, //phyinit_io_write: 0x70072, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h70073, value : 32'h3}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming HwtLpCsEnB to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h39080f, value : 32'h3}, //phyinit_io_write: 0x70073, 0x3
//phyinit_io_write: 0x39080f, 0x3
//[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] End of dwc_ddrphy_phyinit_I_loadPIEImagePsLoop(), PState=3
//[dwc_ddrphy_phyinit_userCustom_customPostTrainPsLoop] End of dwc_ddrphy_phyinit_userCustom_customPostTrainPsLoop(), PState=3
//Start of dwc_ddrphy_phyinit_C_initPhyConfigPsLoop(), PState=0, tck_ps=1250ps
                          '{ step_type : REG_WRITE, reg_addr : 32'h2008b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, programming PState = 0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90801, value : 32'hc0a2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming Seq0BGPR1 to 0xc0a2
                          '{ step_type : REG_WRITE, reg_addr : 32'h90802, value : 32'h0}, //phyinit_io_write: 0x90801, 0xc0a2
                          '{ step_type : REG_WRITE, reg_addr : 32'h90806, value : 32'h1}, //phyinit_io_write: 0x90802, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'ha03ff, value : 32'h4101}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming OdtSeg120 to 0x4101
                          '{ step_type : REG_WRITE, reg_addr : 32'ha030b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming ZCalCompCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h60008, value : 32'h2e9a}, //[dwc_ddrphy_phyinit_programPLL] [phyinit_C_initPhyConfigPsLoop] Pstate=0,  Memclk=800MHz, Programming CpllCtrl5 to 0x2e9a.
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e0, value : 32'h64}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY0 to 0x64 (0.5us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e1, value : 32'h12c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY1 to 0x12c (tZQCal PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e2, value : 32'h7d0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY2 to 0x7d0 (10.us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e3, value : 32'h58}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY3 to 0x58 (dllLock PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e4, value : 32'h14}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY4 to 0x14 (0.1us PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e5, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY5 to 0x0 (RxReplicaCalWait delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e6, value : 32'h43}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY6 to 0x43 (Oscillator PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e7, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY7 to 0x0 (tXDSM_XP PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908ea, value : 32'h4}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY10 to 0x4 (tPDXCSODTON 20ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908eb, value : 32'h4}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY11 to 0x4 (20ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908ec, value : 32'ha}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY12 to 0xa (50ns PIE delay)
                          '{ step_type : REG_WRITE, reg_addr : 32'h908ed, value : 32'h4e}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming Seq0BDLY13 to 0x4e (tXSR PIE delay, tRFCab delay is 380ns)
                          '{ step_type : REG_WRITE, reg_addr : 32'h20002, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming PclkPtrInitVal to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h60040, value : 32'h3}, //phyinit_io_write: 0x20002, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h20000, value : 32'h2}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DfiFreqRatio to 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h100fb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming RxDigStrbEn to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h110fb, value : 32'h0}, //phyinit_io_write: 0x100fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h120fb, value : 32'h0}, //phyinit_io_write: 0x110fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h130fb, value : 32'h0}, //phyinit_io_write: 0x120fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he000b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DxDigStrobeMode HMDBYTE to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he100b, value : 32'h0}, //phyinit_io_write: 0xe000b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he200b, value : 32'h0}, //phyinit_io_write: 0xe100b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he300b, value : 32'h0}, //phyinit_io_write: 0xe200b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he400b, value : 32'h0}, //phyinit_io_write: 0xe300b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he500b, value : 32'h0}, //phyinit_io_write: 0xe400b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he600b, value : 32'h0}, //phyinit_io_write: 0xe500b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he700b, value : 32'h0}, //phyinit_io_write: 0xe600b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE0.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE1.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h12024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE2.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h13024, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE3.DqsPreambleControl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE0.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h11025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE1.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h12025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE2.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h13025, value : 32'h2c}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE3.DbyteRxDqsModeCntrl to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h10004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE0.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10003, value : 32'h0}, //phyinit_io_write: 0x10004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE1.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11003, value : 32'h0}, //phyinit_io_write: 0x11004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h12004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE2.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h12003, value : 32'h0}, //phyinit_io_write: 0x12004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h13004, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE3.DxDfiClkDis to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h13003, value : 32'h0}, //phyinit_io_write: 0x13004, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb0004, value : 32'h320}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ZCalClkInfo::ZCalDfiClkTicksPer1uS to 0x320
                          '{ step_type : REG_WRITE, reg_addr : 32'ha030c, value : 32'h0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003e, value : 32'h5}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE RxGainCurrAdjRxReplica to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103e, value : 32'h5}, //phyinit_io_write: 0x1003e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203e, value : 32'h5}, //phyinit_io_write: 0x1103e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303e, value : 32'h5}, //phyinit_io_write: 0x1203e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h20003, value : 32'h1}, //phyinit_io_write: 0x1303e, 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h2000b, value : 32'h1111}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming CPclkDivRatio to 0x1111
                          '{ step_type : REG_WRITE, reg_addr : 32'h10108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE0.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE1.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h12108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE2.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h13108, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming DBYTE3.DMIPinPresent::RdDbiEnabled to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70005, value : 32'h0}, //[phyinit_C_initPhyConfig] Programming EnPhyUpdZQCalUpdate to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h7000f, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming DisableZQupdateOnSnoop to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1000e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h1100e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h1200e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h1300e, value : 32'h1300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming TrackingModeCntrl to 0x1300
                          '{ step_type : REG_WRITE, reg_addr : 32'h20019, value : 32'h4}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming EnRxDqsTracking::DqsSampNegRxEnSense to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he002c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 0 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he102c, value : 32'h33}, //phyinit_io_write: 0xe002c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'he002d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 0 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he102d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 0 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he202c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 1 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he302c, value : 32'h33}, //phyinit_io_write: 0xe202c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'he202d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 1 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he302d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 1 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he402c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 2 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he502c, value : 32'h33}, //phyinit_io_write: 0xe402c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'he402d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 2 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he502d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 2 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he602c, value : 32'h33}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 3 TxImpedanceDq::TxStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he702c, value : 32'h33}, //phyinit_io_write: 0xe602c, 0x33
                          '{ step_type : REG_WRITE, reg_addr : 32'he602d, value : 32'h303}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 3 TxImpedanceDqs::TxStrenCodeDqsPDC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he702d, value : 32'h3333}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 3 WCK TxImpedanceDqs::TxStrenCodeDqsPDT/C to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h70, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC0 Instance0 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC1 Instance1 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h2070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC2 Instance2 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h3070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC3 Instance3 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h4070, value : 32'hff}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming AC0 HMAC4 Instance4 CS TxImpedanceAC::TxStrenCodePDAC to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'h5070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC5 Instance5 TxImpedanceAC::TxStrenCodePD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h7070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC0 Instance7 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h8070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC1 Instance8 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h9070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC2 Instance9 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'ha070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC3 Instance10 SE TxImpedanceAC::TxStrenCodePDAC to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'hb070, value : 32'hff}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming AC1 HMAC4 Instance11 CS TxImpedanceAC::TxStrenCodePDAC to 0xff
                          '{ step_type : REG_WRITE, reg_addr : 32'hc070, value : 32'h77}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC5 Instance12 TxImpedanceAC::TxStrenCodePD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'he002e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 0 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he102e, value : 32'h30}, //phyinit_io_write: 0xe002e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'he002f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 0 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he102f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 0 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'he202e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 1 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he302e, value : 32'h30}, //phyinit_io_write: 0xe202e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'he202f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 1 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he302f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 1 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'he402e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 2 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he502e, value : 32'h30}, //phyinit_io_write: 0xe402e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'he402f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 2 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he502f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 2 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'he602e, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 3 OdtImpedanceDq::OdtStrenCodeDqPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he702e, value : 32'h30}, //phyinit_io_write: 0xe602e, 0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'he602f, value : 32'h3300}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 3 OdtImpedanceDqs::OdtStrenCodeDqsPD to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he702f, value : 32'h7700}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 3 WCK OdtImpedanceDqs::OdtStrenCodeWckPD to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h79, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC0 Instance0 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h1079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC1 Instance1 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h2079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC2 Instance2 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h3079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC3 Instance3 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h4079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC4 Instance4 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h5079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC5 DIFF5 OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h7079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC0 Instance7 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h8079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC1 Instance8 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h9079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC2 Instance9 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'ha079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC3 Instance10 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'hb079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC4 Instance11 SE OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'hc079, value : 32'h30}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC5 DIFF12 OdtImpedanceAC::OdtStrenCodePDAC to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he001c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 0 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he101c, value : 32'h3}, //phyinit_io_write: 0xe001c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he201c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 1 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he301c, value : 32'h3}, //phyinit_io_write: 0xe201c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he401c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 2 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he501c, value : 32'h3}, //phyinit_io_write: 0xe401c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'he601c, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming HMDBYTE 3 TxDQSlew::TxDQSlewPD to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he701c, value : 32'h3}, //phyinit_io_write: 0xe601c, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h6d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC0 Instance0 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h106d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC1 Instance1 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h206d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC2 Instance2 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h306d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC3 Instance3 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h406d, value : 32'hf8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC4 Instance4 CS TxSlewAC::TxSlewPDAC to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h506d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX0 HMAC5 Instance5 TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h706d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC0 Instance7 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h806d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC1 Instance8 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h906d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC2 Instance9 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'ha06d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC3 Instance10 SE TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb06d, value : 32'hf8}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC4 Instance11 CS TxSlewAC::TxSlewPDAC to 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'hc06d, value : 32'h3}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACX1 HMAC5 Instance12 TxSlewAC::TxSlewPDAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he003e, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Programming HMDBYTE RxDQSCtrl::RxDQSDiffSeVrefDACEn to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he103e, value : 32'h0}, //phyinit_io_write: 0xe003e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he203e, value : 32'h0}, //phyinit_io_write: 0xe103e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he303e, value : 32'h0}, //phyinit_io_write: 0xe203e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he403e, value : 32'h0}, //phyinit_io_write: 0xe303e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he503e, value : 32'h0}, //phyinit_io_write: 0xe403e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he603e, value : 32'h0}, //phyinit_io_write: 0xe503e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he703e, value : 32'h0}, //phyinit_io_write: 0xe603e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10001, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming WriteLinkEcc to 0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11001, value : 32'h0}, //phyinit_io_write: 0x10001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h12001, value : 32'h0}, //phyinit_io_write: 0x11001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h13001, value : 32'h0}, //phyinit_io_write: 0x12001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70040, value : 32'h5a}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming PPTTrainSetup::PhyMstrMaxReqToAck to 0x5
                          '{ step_type : REG_WRITE, reg_addr : 32'h70041, value : 32'hf}, //phyinit_io_write: 0x70040, 0x5a
                          '{ step_type : REG_WRITE, reg_addr : 32'h100a5, value : 32'h1}, //phyinit_io_write: 0x70041, 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h110a5, value : 32'h1}, //phyinit_io_write: 0x100a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h120a5, value : 32'h1}, //phyinit_io_write: 0x110a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h130a5, value : 32'h1}, //phyinit_io_write: 0x120a5, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h10209, value : 32'h3232}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Programming RxReplicaRangeVal 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h11209, value : 32'h3232}, //phyinit_io_write: 0x10209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h12209, value : 32'h3232}, //phyinit_io_write: 0x11209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h13209, value : 32'h3232}, //phyinit_io_write: 0x12209, 0x3232
                          '{ step_type : REG_WRITE, reg_addr : 32'h1020f, value : 32'h6}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Programming RxReplicaCtl04 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h1120f, value : 32'h6}, //phyinit_io_write: 0x1020f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h1220f, value : 32'h6}, //phyinit_io_write: 0x1120f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h1320f, value : 32'h6}, //phyinit_io_write: 0x1220f, 0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h20005, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, DfiFreq=800MHz, Programming PipeCtl[AcInPipeEn]=0x0 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h10008, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, DfiFreq=800MHz, Programming DBYTE0.LP5DfiDataEnLatency[LP5RLm13]=0x1 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h11008, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, DfiFreq=800MHz, Programming DBYTE1.LP5DfiDataEnLatency[LP5RLm13]=0x1 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h12008, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, DfiFreq=800MHz, Programming DBYTE2.LP5DfiDataEnLatency[LP5RLm13]=0x1 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h13008, value : 32'h1}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, DfiFreq=800MHz, Programming DBYTE3.LP5DfiDataEnLatency[LP5RLm13]=0x1 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h7006b, value : 32'h222}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, DfiFreq=800MHz, Programming DfiHandshakeDelays[PhyUpdReqDelay]=0x2 DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h70066, value : 32'h20}, //phyinit_io_write: 0x7006b, 0x222
                          '{ step_type : REG_WRITE, reg_addr : 32'h700eb, value : 32'h222}, //phyinit_io_write: 0x70066, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h700e6, value : 32'h20}, //phyinit_io_write: 0x700eb, 0x222
                          '{ step_type : REG_WRITE, reg_addr : 32'h70135, value : 32'h100c}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACSMWckWriteFastTogglePulse::ACSMWckWriteFastToggleWidth to 0x19, ACSMWckWriteFastTogglePulse::ACSMWckWriteFastToggleDelay to 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h70136, value : 32'h100c}, //phyinit_io_write: 0x70135, 0x100c
                          '{ step_type : REG_WRITE, reg_addr : 32'h70137, value : 32'h41c}, //phyinit_io_write: 0x70136, 0x100c
                          '{ step_type : REG_WRITE, reg_addr : 32'h70138, value : 32'h1920}, //phyinit_io_write: 0x70137, 0x41c
                          '{ step_type : REG_WRITE, reg_addr : 32'h70139, value : 32'h1018}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACSMWckReadFastTogglePulse::ACSMWckReadFastToggleWidth to 0x2d, ACSMWckReadFastTogglePulse::ACSMWckReadFastToggleDelay to 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h7013a, value : 32'h1018}, //phyinit_io_write: 0x70139, 0x1018
                          '{ step_type : REG_WRITE, reg_addr : 32'h7013b, value : 32'h428}, //phyinit_io_write: 0x7013a, 0x1018
                          '{ step_type : REG_WRITE, reg_addr : 32'h7013c, value : 32'h2d2c}, //phyinit_io_write: 0x7013b, 0x428
                          '{ step_type : REG_WRITE, reg_addr : 32'h7013d, value : 32'h1004}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACSMWckFreqFastTogglePulse::ACSMWckFreqFastToggleWidth to 0x11, ACSMWckFreqFastTogglePulse::ACSMWckFreqFastToggleDelay to 0x18
                          '{ step_type : REG_WRITE, reg_addr : 32'h7013e, value : 32'h1004}, //phyinit_io_write: 0x7013d, 0x1004
                          '{ step_type : REG_WRITE, reg_addr : 32'h7013f, value : 32'h414}, //phyinit_io_write: 0x7013e, 0x1004
                          '{ step_type : REG_WRITE, reg_addr : 32'h70140, value : 32'h1118}, //phyinit_io_write: 0x7013f, 0x414
                          '{ step_type : REG_WRITE, reg_addr : 32'h7012c, value : 32'h837}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACSMRxValPulse::ACSMRxValDelay to 0x37, ACSMRxValPulse::ACSMRxValWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h7012d, value : 32'h837}, //phyinit_io_write: 0x7012c, 0x837
                          '{ step_type : REG_WRITE, reg_addr : 32'h70130, value : 32'h837}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACSMRdcsPulse::ACSMRdcsDelay to 0x37, ACSMRdcsPulse::ACSMRdcsWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h7012e, value : 32'h81f}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACSMTxEnPulse::ACSMTxEnDelay to 0x1f, ACSMTxEnPulse::ACSMTxEnWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h7012f, value : 32'h81f}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming ACSMWrcsPulse::ACSMWrcsDelay to 0x1f, ACSMWrcsPulse::ACSMWrcsWidth to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h30008, value : 32'h0}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming AcPipeEn AC0 to 0. DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h31008, value : 32'h0}, //[dwc_ddrphy_phyinit_ACSM_delay] [phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, Programming AcPipeEn AC1 to 0. DFI ratio is 2
                          '{ step_type : REG_WRITE, reg_addr : 32'he0013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he1013, value : 32'h0}, //phyinit_io_write: 0xe0013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he2013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he3013, value : 32'h0}, //phyinit_io_write: 0xe2013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he4013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he5013, value : 32'h0}, //phyinit_io_write: 0xe4013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he6013, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Programming csr_EnaRxStrobeEnB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he7013, value : 32'h0}, //phyinit_io_write: 0xe6013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h5e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC0 Instance0 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h15e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC1 Instance1 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h25e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC2 Instance2 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h35e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC3 Instance3 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h45e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC4 Instance4 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h55e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC5 Instance5 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h75e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC0 Instance7 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h85e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC1 Instance8 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h95e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC2 Instance9 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'ha5e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC3 Instance10 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'hb5e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC4 Instance11 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'hc5e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC5 Instance12 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he05e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming HMDBYTE0 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he15e3, value : 32'h4}, //phyinit_io_write: 0xe05e3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he25e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming HMDBYTE1 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he35e3, value : 32'h4}, //phyinit_io_write: 0xe25e3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he45e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming HMDBYTE2 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he55e3, value : 32'h4}, //phyinit_io_write: 0xe45e3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he65e3, value : 32'h4}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming HMDBYTE3 PclkDCALcdlAddDlySampEn to 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'he75e3, value : 32'h4}, //phyinit_io_write: 0xe65e3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h50a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC0 Instance0 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h150a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC1 Instance1 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h250a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC2 Instance2 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h350a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC3 Instance3 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h450a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC4 Instance4 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h550a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX0 HMAC5 Instance5 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h750a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC0 Instance7 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h850a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC1 Instance8 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h950a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC2 Instance9 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'ha50a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC3 Instance10 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb50a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC4 Instance11 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hc50a, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming ACX1 HMAC5 Instance12 PclkDCASampDelayLCDLAC to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1080b, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming DBYTE0 PclkDCASampDelayLCDLDB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1180b, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming DBYTE1 PclkDCASampDelayLCDLDB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1280b, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming DBYTE2 PclkDCASampDelayLCDLDB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1380b, value : 32'h0}, //[dwc_ddrphy_phyinit_programPclkDca] Programming DBYTE3 PclkDCASampDelayLCDLDB to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30803, value : 32'h106a}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming PclkDCAStaticCtr0AC to 0x106a
                          '{ step_type : REG_WRITE, reg_addr : 32'h31803, value : 32'h106a}, //phyinit_io_write: 0x30803, 0x106a
                          '{ step_type : REG_WRITE, reg_addr : 32'h10803, value : 32'h106a}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming PclkDCAStaticCtr0DB to 0x106a
                          '{ step_type : REG_WRITE, reg_addr : 32'h11803, value : 32'h106a}, //phyinit_io_write: 0x10803, 0x106a
                          '{ step_type : REG_WRITE, reg_addr : 32'h12803, value : 32'h106a}, //phyinit_io_write: 0x11803, 0x106a
                          '{ step_type : REG_WRITE, reg_addr : 32'h13803, value : 32'h106a}, //phyinit_io_write: 0x12803, 0x106a
                          '{ step_type : REG_WRITE, reg_addr : 32'h503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC0 Instance0 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC1 Instance1 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h2503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC2 Instance2 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h3503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC3 Instance3 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h4503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC4 Instance4 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h5503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC5 Instance5 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h7503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC0 Instance7 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h8503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC1 Instance8 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h9503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC2 Instance9 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'ha503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC3 Instance10 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'hb503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC4 Instance11 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'hc503, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC5 Instance12 PclkDCAStaticCtrl1AC to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h10c03, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming PclkDCAStaticCtrl1DB to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h11c03, value : 32'h1f}, //phyinit_io_write: 0x10c03, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h12c03, value : 32'h1f}, //phyinit_io_write: 0x11c03, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h13c03, value : 32'h1f}, //phyinit_io_write: 0x12c03, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC0 Instance0 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h1110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC1 Instance1 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h2110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC2 Instance2 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h3110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC3 Instance3 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h4110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC4 Instance4 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h5110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX0 HMAC5 Instance5 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h7110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC0 Instance7 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h8110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC1 Instance8 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h9110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC2 Instance9 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'ha110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC3 Instance10 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'hb110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC4 Instance11 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'hc110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming ACX1 HMAC5 Instance12 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'he0110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming HMDBYTE0 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'he1110, value : 32'h1f}, //phyinit_io_write: 0xe0110, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'he2110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming HMDBYTE1 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'he3110, value : 32'h1f}, //phyinit_io_write: 0xe2110, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'he4110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming HMDBYTE2 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'he5110, value : 32'h1f}, //phyinit_io_write: 0xe4110, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'he6110, value : 32'h1f}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming HMDBYTE3 PclkDCATxLcdlPhase to 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'he7110, value : 32'h1f}, //phyinit_io_write: 0xe6110, 0x1f
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e8, value : 32'h13}, //[dwc_ddrphy_phyinit_programPclkDca] Pstate=0, Programming Seq0BDLY9 to 64
                          '{ step_type : REG_WRITE, reg_addr : 32'h908e9, value : 32'h40}, //phyinit_io_write: 0x908e8, 0x13
                          '{ step_type : REG_WRITE, reg_addr : 32'he0002, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Programming HMDBYTE RxDFECtrlDq to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he1002, value : 32'h0}, //phyinit_io_write: 0xe0002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he2002, value : 32'h0}, //phyinit_io_write: 0xe1002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he3002, value : 32'h0}, //phyinit_io_write: 0xe2002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he4002, value : 32'h0}, //phyinit_io_write: 0xe3002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he5002, value : 32'h0}, //phyinit_io_write: 0xe4002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he6002, value : 32'h0}, //phyinit_io_write: 0xe5002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'he7002, value : 32'h0}, //phyinit_io_write: 0xe6002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1010b, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Pstate=0, Memclk=800MHz, freqThreshold=200MHz, NoRDQS=0 Programming InhibitTxRdPtrInit::DisableRxEnDlyLoad to 0x0, InhibitTxRdPtrInit::DisableTxDqDly to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1110b, value : 32'h0}, //phyinit_io_write: 0x1010b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1210b, value : 32'h0}, //phyinit_io_write: 0x1110b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1310b, value : 32'h0}, //phyinit_io_write: 0x1210b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h63, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC0 Instance0 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h1063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC1 Instance1 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h2063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC2 Instance2 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h3063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC3 Instance3 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h4063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC4 Instance4 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h5063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC5 Instance5 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h7063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC0 Instance7 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h8063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC1 Instance8 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h9063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC2 Instance9 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'ha063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC3 Instance10 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'hb063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC4 Instance11 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'hc063, value : 32'h68}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC5 Instance12 HMTxLcdlSeed HMTxSeed to 0x68 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h9080a, value : 32'h268}, //[dwc_ddrphy_phyinit_programLCDLSeed] Programming Seq0BGPR10 to HMTxLcdlSeed Full search value = 0x268
                          '{ step_type : REG_WRITE, reg_addr : 32'h9080b, value : 32'h68}, //phyinit_io_write: 0x9080a, 0x268
                          '{ step_type : REG_WRITE, reg_addr : 32'h90815, value : 32'h268}, //[dwc_ddrphy_phyinit_programLCDLSeed] Programming Seq0BGPR21 to ACHMTxLcdlSeed Full search value = 0x268
                          '{ step_type : REG_WRITE, reg_addr : 32'h90816, value : 32'h68}, //phyinit_io_write: 0x90815, 0x268
                          '{ step_type : REG_WRITE, reg_addr : 32'he0063, value : 32'h68}, //phyinit_io_write: 0x90816, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he0064, value : 32'h68}, //phyinit_io_write: 0xe0063, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he0087, value : 32'h68}, //phyinit_io_write: 0xe0064, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he1063, value : 32'h68}, //phyinit_io_write: 0xe0087, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he1064, value : 32'h68}, //phyinit_io_write: 0xe1063, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he1087, value : 32'h68}, //phyinit_io_write: 0xe1064, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he2063, value : 32'h68}, //phyinit_io_write: 0xe1087, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he2064, value : 32'h68}, //phyinit_io_write: 0xe2063, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he2087, value : 32'h68}, //phyinit_io_write: 0xe2064, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he3063, value : 32'h68}, //phyinit_io_write: 0xe2087, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he3064, value : 32'h68}, //phyinit_io_write: 0xe3063, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he3087, value : 32'h68}, //phyinit_io_write: 0xe3064, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he4063, value : 32'h68}, //phyinit_io_write: 0xe3087, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he4064, value : 32'h68}, //phyinit_io_write: 0xe4063, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he4087, value : 32'h68}, //phyinit_io_write: 0xe4064, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he5063, value : 32'h68}, //phyinit_io_write: 0xe4087, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he5064, value : 32'h68}, //phyinit_io_write: 0xe5063, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he5087, value : 32'h68}, //phyinit_io_write: 0xe5064, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he6063, value : 32'h68}, //phyinit_io_write: 0xe5087, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he6064, value : 32'h68}, //phyinit_io_write: 0xe6063, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he6087, value : 32'h68}, //phyinit_io_write: 0xe6064, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he7063, value : 32'h68}, //phyinit_io_write: 0xe6087, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he7064, value : 32'h68}, //phyinit_io_write: 0xe7063, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'he7087, value : 32'h68}, //phyinit_io_write: 0xe7064, 0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0080, value : 32'h7}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming UcclkHclkEnables to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'he003c, value : 32'h80}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming RxDQSSeVrefDAC0 to 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'he103c, value : 32'h80}, //phyinit_io_write: 0xe003c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'he203c, value : 32'h80}, //phyinit_io_write: 0xe103c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'he303c, value : 32'h80}, //phyinit_io_write: 0xe203c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'he403c, value : 32'h80}, //phyinit_io_write: 0xe303c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'he503c, value : 32'h80}, //phyinit_io_write: 0xe403c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'he603c, value : 32'h80}, //phyinit_io_write: 0xe503c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'he703c, value : 32'h80}, //phyinit_io_write: 0xe603c, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h90817, value : 32'h53}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 0 Seq0BGPR23 to 0x53, NumMemClk_tRFCab=328.0, NumMemClk_7p5ns=6.0, NumMemClk_tXSR=334.0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90818, value : 32'h0}, //phyinit_io_write: 0x90817, 0x53
                          '{ step_type : REG_WRITE, reg_addr : 32'h90819, value : 32'h0}, //phyinit_io_write: 0x90818, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h300eb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 0 AC0 AcLcdlUpdInterval to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h310eb, value : 32'h0}, //[dwc_ddrphy_phyinit_C_initPhyConfigPsLoop] Programming PState 0 AC1 AcLcdlUpdInterval to 0x0
//[dwc_ddrphy_phyinit_programDfiMode] Skip DfiMode Programming: Keeping the reset value of 0x3
//End of dwc_ddrphy_phyinit_C_initPhyConfigPsLoop(), Pstate=0
                          '{ step_type : REG_WRITE, reg_addr : 32'h300d9, value : 32'h40}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming CKXTxDly to 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h300d8, value : 32'h40}, //phyinit_io_write: 0x300d9, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h301d8, value : 32'h40}, //phyinit_io_write: 0x300d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h302d8, value : 32'h40}, //phyinit_io_write: 0x301d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h303d8, value : 32'h40}, //phyinit_io_write: 0x302d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h304d8, value : 32'h40}, //phyinit_io_write: 0x303d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h305d8, value : 32'h40}, //phyinit_io_write: 0x304d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h306d8, value : 32'h40}, //phyinit_io_write: 0x305d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h308d8, value : 32'h40}, //phyinit_io_write: 0x306d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h309d8, value : 32'h40}, //phyinit_io_write: 0x308d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h310d9, value : 32'h40}, //phyinit_io_write: 0x309d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h310d8, value : 32'h40}, //phyinit_io_write: 0x310d9, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h311d8, value : 32'h40}, //phyinit_io_write: 0x310d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h312d8, value : 32'h40}, //phyinit_io_write: 0x311d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h313d8, value : 32'h40}, //phyinit_io_write: 0x312d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h314d8, value : 32'h40}, //phyinit_io_write: 0x313d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h315d8, value : 32'h40}, //phyinit_io_write: 0x314d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h316d8, value : 32'h40}, //phyinit_io_write: 0x315d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h318d8, value : 32'h40}, //phyinit_io_write: 0x316d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h319d8, value : 32'h40}, //phyinit_io_write: 0x318d8, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h10000, value : 32'h7}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming HwtMRL to 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h11000, value : 32'h7}, //phyinit_io_write: 0x10000, 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h12000, value : 32'h7}, //phyinit_io_write: 0x11000, 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h13000, value : 32'h7}, //phyinit_io_write: 0x12000, 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h7000d, value : 32'h7}, //phyinit_io_write: 0x13000, 0x7
                          '{ step_type : REG_WRITE, reg_addr : 32'h1002a, value : 32'h200}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming TxWckDlyTg0/Tg1 to 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h1002b, value : 32'h200}, //phyinit_io_write: 0x1002a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102a, value : 32'h200}, //phyinit_io_write: 0x1002b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h1102b, value : 32'h200}, //phyinit_io_write: 0x1102a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h1202a, value : 32'h200}, //phyinit_io_write: 0x1102b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h1202b, value : 32'h200}, //phyinit_io_write: 0x1202a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h1302a, value : 32'h200}, //phyinit_io_write: 0x1202b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h1302b, value : 32'h200}, //phyinit_io_write: 0x1302a, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h10028, value : 32'hed}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming TxDqsDlyTg0/Tg1 to 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h10029, value : 32'hed}, //phyinit_io_write: 0x10028, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h11028, value : 32'hed}, //phyinit_io_write: 0x10029, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h11029, value : 32'hed}, //phyinit_io_write: 0x11028, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h12028, value : 32'hed}, //phyinit_io_write: 0x11029, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h12029, value : 32'hed}, //phyinit_io_write: 0x12028, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h13028, value : 32'hed}, //phyinit_io_write: 0x12029, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h13029, value : 32'hed}, //phyinit_io_write: 0x13028, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1007a, value : 32'hed}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming TxDqDlyTg0/Tg1 to 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1007b, value : 32'hed}, //phyinit_io_write: 0x1007a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1017a, value : 32'hed}, //phyinit_io_write: 0x1007b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1017b, value : 32'hed}, //phyinit_io_write: 0x1017a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1027a, value : 32'hed}, //phyinit_io_write: 0x1017b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1027b, value : 32'hed}, //phyinit_io_write: 0x1027a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1037a, value : 32'hed}, //phyinit_io_write: 0x1027b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1037b, value : 32'hed}, //phyinit_io_write: 0x1037a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1047a, value : 32'hed}, //phyinit_io_write: 0x1037b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1047b, value : 32'hed}, //phyinit_io_write: 0x1047a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1057a, value : 32'hed}, //phyinit_io_write: 0x1047b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1057b, value : 32'hed}, //phyinit_io_write: 0x1057a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1067a, value : 32'hed}, //phyinit_io_write: 0x1057b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1067b, value : 32'hed}, //phyinit_io_write: 0x1067a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1077a, value : 32'hed}, //phyinit_io_write: 0x1067b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1077b, value : 32'hed}, //phyinit_io_write: 0x1077a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1087a, value : 32'hed}, //phyinit_io_write: 0x1077b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1087b, value : 32'hed}, //phyinit_io_write: 0x1087a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1107a, value : 32'hed}, //phyinit_io_write: 0x1087b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1107b, value : 32'hed}, //phyinit_io_write: 0x1107a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1117a, value : 32'hed}, //phyinit_io_write: 0x1107b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1117b, value : 32'hed}, //phyinit_io_write: 0x1117a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1127a, value : 32'hed}, //phyinit_io_write: 0x1117b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1127b, value : 32'hed}, //phyinit_io_write: 0x1127a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1137a, value : 32'hed}, //phyinit_io_write: 0x1127b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1137b, value : 32'hed}, //phyinit_io_write: 0x1137a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1147a, value : 32'hed}, //phyinit_io_write: 0x1137b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1147b, value : 32'hed}, //phyinit_io_write: 0x1147a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1157a, value : 32'hed}, //phyinit_io_write: 0x1147b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1157b, value : 32'hed}, //phyinit_io_write: 0x1157a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1167a, value : 32'hed}, //phyinit_io_write: 0x1157b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1167b, value : 32'hed}, //phyinit_io_write: 0x1167a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1177a, value : 32'hed}, //phyinit_io_write: 0x1167b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1177b, value : 32'hed}, //phyinit_io_write: 0x1177a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1187a, value : 32'hed}, //phyinit_io_write: 0x1177b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1187b, value : 32'hed}, //phyinit_io_write: 0x1187a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1207a, value : 32'hed}, //phyinit_io_write: 0x1187b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1207b, value : 32'hed}, //phyinit_io_write: 0x1207a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1217a, value : 32'hed}, //phyinit_io_write: 0x1207b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1217b, value : 32'hed}, //phyinit_io_write: 0x1217a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1227a, value : 32'hed}, //phyinit_io_write: 0x1217b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1227b, value : 32'hed}, //phyinit_io_write: 0x1227a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1237a, value : 32'hed}, //phyinit_io_write: 0x1227b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1237b, value : 32'hed}, //phyinit_io_write: 0x1237a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1247a, value : 32'hed}, //phyinit_io_write: 0x1237b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1247b, value : 32'hed}, //phyinit_io_write: 0x1247a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1257a, value : 32'hed}, //phyinit_io_write: 0x1247b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1257b, value : 32'hed}, //phyinit_io_write: 0x1257a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1267a, value : 32'hed}, //phyinit_io_write: 0x1257b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1267b, value : 32'hed}, //phyinit_io_write: 0x1267a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1277a, value : 32'hed}, //phyinit_io_write: 0x1267b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1277b, value : 32'hed}, //phyinit_io_write: 0x1277a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1287a, value : 32'hed}, //phyinit_io_write: 0x1277b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1287b, value : 32'hed}, //phyinit_io_write: 0x1287a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1307a, value : 32'hed}, //phyinit_io_write: 0x1287b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1307b, value : 32'hed}, //phyinit_io_write: 0x1307a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1317a, value : 32'hed}, //phyinit_io_write: 0x1307b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1317b, value : 32'hed}, //phyinit_io_write: 0x1317a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1327a, value : 32'hed}, //phyinit_io_write: 0x1317b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1327b, value : 32'hed}, //phyinit_io_write: 0x1327a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1337a, value : 32'hed}, //phyinit_io_write: 0x1327b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1337b, value : 32'hed}, //phyinit_io_write: 0x1337a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1347a, value : 32'hed}, //phyinit_io_write: 0x1337b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1347b, value : 32'hed}, //phyinit_io_write: 0x1347a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1357a, value : 32'hed}, //phyinit_io_write: 0x1347b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1357b, value : 32'hed}, //phyinit_io_write: 0x1357a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1367a, value : 32'hed}, //phyinit_io_write: 0x1357b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1367b, value : 32'hed}, //phyinit_io_write: 0x1367a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1377a, value : 32'hed}, //phyinit_io_write: 0x1367b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1377b, value : 32'hed}, //phyinit_io_write: 0x1377a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1387a, value : 32'hed}, //phyinit_io_write: 0x1377b, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h1387b, value : 32'hed}, //phyinit_io_write: 0x1387a, 0xed
                          '{ step_type : REG_WRITE, reg_addr : 32'h10078, value : 32'h3b9}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming RxDigStrbDlyTg0/Tg1 to 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10079, value : 32'h3b9}, //phyinit_io_write: 0x10078, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10178, value : 32'h3b9}, //phyinit_io_write: 0x10079, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10179, value : 32'h3b9}, //phyinit_io_write: 0x10178, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10278, value : 32'h3b9}, //phyinit_io_write: 0x10179, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10279, value : 32'h3b9}, //phyinit_io_write: 0x10278, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10378, value : 32'h3b9}, //phyinit_io_write: 0x10279, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10379, value : 32'h3b9}, //phyinit_io_write: 0x10378, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10478, value : 32'h3b9}, //phyinit_io_write: 0x10379, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10479, value : 32'h3b9}, //phyinit_io_write: 0x10478, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10578, value : 32'h3b9}, //phyinit_io_write: 0x10479, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10579, value : 32'h3b9}, //phyinit_io_write: 0x10578, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10678, value : 32'h3b9}, //phyinit_io_write: 0x10579, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10679, value : 32'h3b9}, //phyinit_io_write: 0x10678, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10778, value : 32'h3b9}, //phyinit_io_write: 0x10679, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10779, value : 32'h3b9}, //phyinit_io_write: 0x10778, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10878, value : 32'h3b9}, //phyinit_io_write: 0x10779, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10879, value : 32'h3b9}, //phyinit_io_write: 0x10878, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11078, value : 32'h3b9}, //phyinit_io_write: 0x10879, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11079, value : 32'h3b9}, //phyinit_io_write: 0x11078, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11178, value : 32'h3b9}, //phyinit_io_write: 0x11079, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11179, value : 32'h3b9}, //phyinit_io_write: 0x11178, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11278, value : 32'h3b9}, //phyinit_io_write: 0x11179, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11279, value : 32'h3b9}, //phyinit_io_write: 0x11278, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11378, value : 32'h3b9}, //phyinit_io_write: 0x11279, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11379, value : 32'h3b9}, //phyinit_io_write: 0x11378, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11478, value : 32'h3b9}, //phyinit_io_write: 0x11379, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11479, value : 32'h3b9}, //phyinit_io_write: 0x11478, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11578, value : 32'h3b9}, //phyinit_io_write: 0x11479, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11579, value : 32'h3b9}, //phyinit_io_write: 0x11578, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11678, value : 32'h3b9}, //phyinit_io_write: 0x11579, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11679, value : 32'h3b9}, //phyinit_io_write: 0x11678, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11778, value : 32'h3b9}, //phyinit_io_write: 0x11679, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11779, value : 32'h3b9}, //phyinit_io_write: 0x11778, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11878, value : 32'h3b9}, //phyinit_io_write: 0x11779, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h11879, value : 32'h3b9}, //phyinit_io_write: 0x11878, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12078, value : 32'h3b9}, //phyinit_io_write: 0x11879, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12079, value : 32'h3b9}, //phyinit_io_write: 0x12078, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12178, value : 32'h3b9}, //phyinit_io_write: 0x12079, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12179, value : 32'h3b9}, //phyinit_io_write: 0x12178, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12278, value : 32'h3b9}, //phyinit_io_write: 0x12179, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12279, value : 32'h3b9}, //phyinit_io_write: 0x12278, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12378, value : 32'h3b9}, //phyinit_io_write: 0x12279, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12379, value : 32'h3b9}, //phyinit_io_write: 0x12378, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12478, value : 32'h3b9}, //phyinit_io_write: 0x12379, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12479, value : 32'h3b9}, //phyinit_io_write: 0x12478, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12578, value : 32'h3b9}, //phyinit_io_write: 0x12479, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12579, value : 32'h3b9}, //phyinit_io_write: 0x12578, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12678, value : 32'h3b9}, //phyinit_io_write: 0x12579, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12679, value : 32'h3b9}, //phyinit_io_write: 0x12678, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12778, value : 32'h3b9}, //phyinit_io_write: 0x12679, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12779, value : 32'h3b9}, //phyinit_io_write: 0x12778, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12878, value : 32'h3b9}, //phyinit_io_write: 0x12779, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h12879, value : 32'h3b9}, //phyinit_io_write: 0x12878, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13078, value : 32'h3b9}, //phyinit_io_write: 0x12879, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13079, value : 32'h3b9}, //phyinit_io_write: 0x13078, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13178, value : 32'h3b9}, //phyinit_io_write: 0x13079, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13179, value : 32'h3b9}, //phyinit_io_write: 0x13178, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13278, value : 32'h3b9}, //phyinit_io_write: 0x13179, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13279, value : 32'h3b9}, //phyinit_io_write: 0x13278, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13378, value : 32'h3b9}, //phyinit_io_write: 0x13279, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13379, value : 32'h3b9}, //phyinit_io_write: 0x13378, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13478, value : 32'h3b9}, //phyinit_io_write: 0x13379, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13479, value : 32'h3b9}, //phyinit_io_write: 0x13478, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13578, value : 32'h3b9}, //phyinit_io_write: 0x13479, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13579, value : 32'h3b9}, //phyinit_io_write: 0x13578, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13678, value : 32'h3b9}, //phyinit_io_write: 0x13579, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13679, value : 32'h3b9}, //phyinit_io_write: 0x13678, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13778, value : 32'h3b9}, //phyinit_io_write: 0x13679, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13779, value : 32'h3b9}, //phyinit_io_write: 0x13778, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13878, value : 32'h3b9}, //phyinit_io_write: 0x13779, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h13879, value : 32'h3b9}, //phyinit_io_write: 0x13878, 0x3b9
                          '{ step_type : REG_WRITE, reg_addr : 32'h10020, value : 32'h319}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming RxEnDlyTg0/Tg1 to 0x319
                          '{ step_type : REG_WRITE, reg_addr : 32'h10021, value : 32'h319}, //phyinit_io_write: 0x10020, 0x319
                          '{ step_type : REG_WRITE, reg_addr : 32'h11020, value : 32'h319}, //phyinit_io_write: 0x10021, 0x319
                          '{ step_type : REG_WRITE, reg_addr : 32'h11021, value : 32'h319}, //phyinit_io_write: 0x11020, 0x319
                          '{ step_type : REG_WRITE, reg_addr : 32'h12020, value : 32'h319}, //phyinit_io_write: 0x11021, 0x319
                          '{ step_type : REG_WRITE, reg_addr : 32'h12021, value : 32'h319}, //phyinit_io_write: 0x12020, 0x319
                          '{ step_type : REG_WRITE, reg_addr : 32'h13020, value : 32'h319}, //phyinit_io_write: 0x12021, 0x319
                          '{ step_type : REG_WRITE, reg_addr : 32'h13021, value : 32'h319}, //phyinit_io_write: 0x13020, 0x319
                          '{ step_type : REG_WRITE, reg_addr : 32'h10010, value : 32'h12b}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming RxClkT2UIDlyTg0/Tg1 and RxClkC2UIDlyTg0/Tg1 to 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10011, value : 32'h12b}, //phyinit_io_write: 0x10010, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10012, value : 32'h12b}, //phyinit_io_write: 0x10011, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10013, value : 32'h12b}, //phyinit_io_write: 0x10012, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10110, value : 32'h12b}, //phyinit_io_write: 0x10013, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10111, value : 32'h12b}, //phyinit_io_write: 0x10110, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10112, value : 32'h12b}, //phyinit_io_write: 0x10111, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10113, value : 32'h12b}, //phyinit_io_write: 0x10112, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10210, value : 32'h12b}, //phyinit_io_write: 0x10113, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10211, value : 32'h12b}, //phyinit_io_write: 0x10210, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10212, value : 32'h12b}, //phyinit_io_write: 0x10211, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10213, value : 32'h12b}, //phyinit_io_write: 0x10212, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10310, value : 32'h12b}, //phyinit_io_write: 0x10213, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10311, value : 32'h12b}, //phyinit_io_write: 0x10310, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10312, value : 32'h12b}, //phyinit_io_write: 0x10311, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10313, value : 32'h12b}, //phyinit_io_write: 0x10312, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10410, value : 32'h12b}, //phyinit_io_write: 0x10313, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10411, value : 32'h12b}, //phyinit_io_write: 0x10410, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10412, value : 32'h12b}, //phyinit_io_write: 0x10411, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10413, value : 32'h12b}, //phyinit_io_write: 0x10412, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10510, value : 32'h12b}, //phyinit_io_write: 0x10413, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10511, value : 32'h12b}, //phyinit_io_write: 0x10510, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10512, value : 32'h12b}, //phyinit_io_write: 0x10511, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10513, value : 32'h12b}, //phyinit_io_write: 0x10512, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10610, value : 32'h12b}, //phyinit_io_write: 0x10513, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10611, value : 32'h12b}, //phyinit_io_write: 0x10610, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10612, value : 32'h12b}, //phyinit_io_write: 0x10611, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10613, value : 32'h12b}, //phyinit_io_write: 0x10612, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10710, value : 32'h12b}, //phyinit_io_write: 0x10613, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10711, value : 32'h12b}, //phyinit_io_write: 0x10710, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10712, value : 32'h12b}, //phyinit_io_write: 0x10711, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10713, value : 32'h12b}, //phyinit_io_write: 0x10712, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10810, value : 32'h12b}, //phyinit_io_write: 0x10713, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10811, value : 32'h12b}, //phyinit_io_write: 0x10810, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10812, value : 32'h12b}, //phyinit_io_write: 0x10811, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h10813, value : 32'h12b}, //phyinit_io_write: 0x10812, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11010, value : 32'h12b}, //phyinit_io_write: 0x10813, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11011, value : 32'h12b}, //phyinit_io_write: 0x11010, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11012, value : 32'h12b}, //phyinit_io_write: 0x11011, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11013, value : 32'h12b}, //phyinit_io_write: 0x11012, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11110, value : 32'h12b}, //phyinit_io_write: 0x11013, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11111, value : 32'h12b}, //phyinit_io_write: 0x11110, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11112, value : 32'h12b}, //phyinit_io_write: 0x11111, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11113, value : 32'h12b}, //phyinit_io_write: 0x11112, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11210, value : 32'h12b}, //phyinit_io_write: 0x11113, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11211, value : 32'h12b}, //phyinit_io_write: 0x11210, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11212, value : 32'h12b}, //phyinit_io_write: 0x11211, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11213, value : 32'h12b}, //phyinit_io_write: 0x11212, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11310, value : 32'h12b}, //phyinit_io_write: 0x11213, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11311, value : 32'h12b}, //phyinit_io_write: 0x11310, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11312, value : 32'h12b}, //phyinit_io_write: 0x11311, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11313, value : 32'h12b}, //phyinit_io_write: 0x11312, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11410, value : 32'h12b}, //phyinit_io_write: 0x11313, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11411, value : 32'h12b}, //phyinit_io_write: 0x11410, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11412, value : 32'h12b}, //phyinit_io_write: 0x11411, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11413, value : 32'h12b}, //phyinit_io_write: 0x11412, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11510, value : 32'h12b}, //phyinit_io_write: 0x11413, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11511, value : 32'h12b}, //phyinit_io_write: 0x11510, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11512, value : 32'h12b}, //phyinit_io_write: 0x11511, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11513, value : 32'h12b}, //phyinit_io_write: 0x11512, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11610, value : 32'h12b}, //phyinit_io_write: 0x11513, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11611, value : 32'h12b}, //phyinit_io_write: 0x11610, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11612, value : 32'h12b}, //phyinit_io_write: 0x11611, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11613, value : 32'h12b}, //phyinit_io_write: 0x11612, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11710, value : 32'h12b}, //phyinit_io_write: 0x11613, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11711, value : 32'h12b}, //phyinit_io_write: 0x11710, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11712, value : 32'h12b}, //phyinit_io_write: 0x11711, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11713, value : 32'h12b}, //phyinit_io_write: 0x11712, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11810, value : 32'h12b}, //phyinit_io_write: 0x11713, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11811, value : 32'h12b}, //phyinit_io_write: 0x11810, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11812, value : 32'h12b}, //phyinit_io_write: 0x11811, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h11813, value : 32'h12b}, //phyinit_io_write: 0x11812, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12010, value : 32'h12b}, //phyinit_io_write: 0x11813, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12011, value : 32'h12b}, //phyinit_io_write: 0x12010, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12012, value : 32'h12b}, //phyinit_io_write: 0x12011, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12013, value : 32'h12b}, //phyinit_io_write: 0x12012, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12110, value : 32'h12b}, //phyinit_io_write: 0x12013, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12111, value : 32'h12b}, //phyinit_io_write: 0x12110, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12112, value : 32'h12b}, //phyinit_io_write: 0x12111, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12113, value : 32'h12b}, //phyinit_io_write: 0x12112, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12210, value : 32'h12b}, //phyinit_io_write: 0x12113, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12211, value : 32'h12b}, //phyinit_io_write: 0x12210, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12212, value : 32'h12b}, //phyinit_io_write: 0x12211, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12213, value : 32'h12b}, //phyinit_io_write: 0x12212, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12310, value : 32'h12b}, //phyinit_io_write: 0x12213, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12311, value : 32'h12b}, //phyinit_io_write: 0x12310, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12312, value : 32'h12b}, //phyinit_io_write: 0x12311, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12313, value : 32'h12b}, //phyinit_io_write: 0x12312, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12410, value : 32'h12b}, //phyinit_io_write: 0x12313, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12411, value : 32'h12b}, //phyinit_io_write: 0x12410, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12412, value : 32'h12b}, //phyinit_io_write: 0x12411, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12413, value : 32'h12b}, //phyinit_io_write: 0x12412, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12510, value : 32'h12b}, //phyinit_io_write: 0x12413, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12511, value : 32'h12b}, //phyinit_io_write: 0x12510, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12512, value : 32'h12b}, //phyinit_io_write: 0x12511, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12513, value : 32'h12b}, //phyinit_io_write: 0x12512, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12610, value : 32'h12b}, //phyinit_io_write: 0x12513, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12611, value : 32'h12b}, //phyinit_io_write: 0x12610, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12612, value : 32'h12b}, //phyinit_io_write: 0x12611, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12613, value : 32'h12b}, //phyinit_io_write: 0x12612, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12710, value : 32'h12b}, //phyinit_io_write: 0x12613, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12711, value : 32'h12b}, //phyinit_io_write: 0x12710, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12712, value : 32'h12b}, //phyinit_io_write: 0x12711, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12713, value : 32'h12b}, //phyinit_io_write: 0x12712, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12810, value : 32'h12b}, //phyinit_io_write: 0x12713, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12811, value : 32'h12b}, //phyinit_io_write: 0x12810, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12812, value : 32'h12b}, //phyinit_io_write: 0x12811, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h12813, value : 32'h12b}, //phyinit_io_write: 0x12812, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13010, value : 32'h12b}, //phyinit_io_write: 0x12813, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13011, value : 32'h12b}, //phyinit_io_write: 0x13010, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13012, value : 32'h12b}, //phyinit_io_write: 0x13011, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13013, value : 32'h12b}, //phyinit_io_write: 0x13012, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13110, value : 32'h12b}, //phyinit_io_write: 0x13013, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13111, value : 32'h12b}, //phyinit_io_write: 0x13110, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13112, value : 32'h12b}, //phyinit_io_write: 0x13111, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13113, value : 32'h12b}, //phyinit_io_write: 0x13112, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13210, value : 32'h12b}, //phyinit_io_write: 0x13113, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13211, value : 32'h12b}, //phyinit_io_write: 0x13210, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13212, value : 32'h12b}, //phyinit_io_write: 0x13211, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13213, value : 32'h12b}, //phyinit_io_write: 0x13212, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13310, value : 32'h12b}, //phyinit_io_write: 0x13213, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13311, value : 32'h12b}, //phyinit_io_write: 0x13310, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13312, value : 32'h12b}, //phyinit_io_write: 0x13311, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13313, value : 32'h12b}, //phyinit_io_write: 0x13312, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13410, value : 32'h12b}, //phyinit_io_write: 0x13313, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13411, value : 32'h12b}, //phyinit_io_write: 0x13410, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13412, value : 32'h12b}, //phyinit_io_write: 0x13411, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13413, value : 32'h12b}, //phyinit_io_write: 0x13412, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13510, value : 32'h12b}, //phyinit_io_write: 0x13413, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13511, value : 32'h12b}, //phyinit_io_write: 0x13510, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13512, value : 32'h12b}, //phyinit_io_write: 0x13511, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13513, value : 32'h12b}, //phyinit_io_write: 0x13512, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13610, value : 32'h12b}, //phyinit_io_write: 0x13513, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13611, value : 32'h12b}, //phyinit_io_write: 0x13610, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13612, value : 32'h12b}, //phyinit_io_write: 0x13611, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13613, value : 32'h12b}, //phyinit_io_write: 0x13612, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13710, value : 32'h12b}, //phyinit_io_write: 0x13613, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13711, value : 32'h12b}, //phyinit_io_write: 0x13710, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13712, value : 32'h12b}, //phyinit_io_write: 0x13711, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13713, value : 32'h12b}, //phyinit_io_write: 0x13712, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13810, value : 32'h12b}, //phyinit_io_write: 0x13713, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13811, value : 32'h12b}, //phyinit_io_write: 0x13810, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13812, value : 32'h12b}, //phyinit_io_write: 0x13811, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h13813, value : 32'h12b}, //phyinit_io_write: 0x13812, 0x12b
                          '{ step_type : REG_WRITE, reg_addr : 32'h1000c, value : 32'hcc}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming PptWck2DqoCntInvTrn1 to 0x198
                          '{ step_type : REG_WRITE, reg_addr : 32'h1000d, value : 32'hcc}, //phyinit_io_write: 0x1000c, 0xcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h10014, value : 32'h198}, //phyinit_io_write: 0x1000d, 0xcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h10015, value : 32'h198}, //phyinit_io_write: 0x10014, 0x198
                          '{ step_type : REG_WRITE, reg_addr : 32'h1100c, value : 32'hcc}, //phyinit_io_write: 0x10015, 0x198
                          '{ step_type : REG_WRITE, reg_addr : 32'h1100d, value : 32'hcc}, //phyinit_io_write: 0x1100c, 0xcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h11014, value : 32'h198}, //phyinit_io_write: 0x1100d, 0xcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h11015, value : 32'h198}, //phyinit_io_write: 0x11014, 0x198
                          '{ step_type : REG_WRITE, reg_addr : 32'h1200c, value : 32'hcc}, //phyinit_io_write: 0x11015, 0x198
                          '{ step_type : REG_WRITE, reg_addr : 32'h1200d, value : 32'hcc}, //phyinit_io_write: 0x1200c, 0xcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h12014, value : 32'h198}, //phyinit_io_write: 0x1200d, 0xcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h12015, value : 32'h198}, //phyinit_io_write: 0x12014, 0x198
                          '{ step_type : REG_WRITE, reg_addr : 32'h1300c, value : 32'hcc}, //phyinit_io_write: 0x12015, 0x198
                          '{ step_type : REG_WRITE, reg_addr : 32'h1300d, value : 32'hcc}, //phyinit_io_write: 0x1300c, 0xcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h13014, value : 32'h198}, //phyinit_io_write: 0x1300d, 0xcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h13015, value : 32'h198}, //phyinit_io_write: 0x13014, 0x198
                          '{ step_type : REG_WRITE, reg_addr : 32'h70077, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming HwtCtrl to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h20071, value : 32'h66}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming HMRxReplicaLcdlSeed HMRxSeed to 0x62 HMRxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h63, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC0 Instance0 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h1063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC1 Instance1 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h2063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC2 Instance2 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h3063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC3 Instance3 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h4063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC4 Instance4 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h5063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX0 HMAC5 Instance5 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h7063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC0 Instance7 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h8063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC1 Instance8 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'h9063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC2 Instance9 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'ha063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC3 Instance10 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'hb063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC4 Instance11 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'hc063, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] LcdlSeed Pstate=0, Memclk=800MHz, Programming ACX1 HMAC5 Instance12 HMTxLcdlSeed HMTxSeed to 0x62 HMTxSeedIs1UI 0x0 
                          '{ step_type : REG_WRITE, reg_addr : 32'he0063, value : 32'h62}, //phyinit_io_write: 0xc063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he0064, value : 32'h62}, //phyinit_io_write: 0xe0063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he0087, value : 32'h62}, //phyinit_io_write: 0xe0064, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he1063, value : 32'h62}, //phyinit_io_write: 0xe0087, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he1064, value : 32'h62}, //phyinit_io_write: 0xe1063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he1087, value : 32'h62}, //phyinit_io_write: 0xe1064, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he2063, value : 32'h62}, //phyinit_io_write: 0xe1087, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he2064, value : 32'h62}, //phyinit_io_write: 0xe2063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he2087, value : 32'h62}, //phyinit_io_write: 0xe2064, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he3063, value : 32'h62}, //phyinit_io_write: 0xe2087, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he3064, value : 32'h62}, //phyinit_io_write: 0xe3063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he3087, value : 32'h62}, //phyinit_io_write: 0xe3064, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he4063, value : 32'h62}, //phyinit_io_write: 0xe3087, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he4064, value : 32'h62}, //phyinit_io_write: 0xe4063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he4087, value : 32'h62}, //phyinit_io_write: 0xe4064, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he5063, value : 32'h62}, //phyinit_io_write: 0xe4087, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he5064, value : 32'h62}, //phyinit_io_write: 0xe5063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he5087, value : 32'h62}, //phyinit_io_write: 0xe5064, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he6063, value : 32'h62}, //phyinit_io_write: 0xe5087, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he6064, value : 32'h62}, //phyinit_io_write: 0xe6063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he6087, value : 32'h62}, //phyinit_io_write: 0xe6064, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he7063, value : 32'h62}, //phyinit_io_write: 0xe6087, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he7064, value : 32'h62}, //phyinit_io_write: 0xe7063, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'he7087, value : 32'h62}, //phyinit_io_write: 0xe7064, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'h9080a, value : 32'h262}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=0 Programming Seq0bGPR10 to mission mode HMTxLcdlSeed value 0x262
                          '{ step_type : REG_WRITE, reg_addr : 32'h9080b, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=0 Programming Seq0bGPR11 to mission mode HMTxLcdlSeed value 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'h90815, value : 32'h262}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=0 Programming Seq0bGPR21 to mission mode HMTxLcdlSeed value 0x262
                          '{ step_type : REG_WRITE, reg_addr : 32'h90816, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=0 Programming Seq0bGPR22 to mission mode HMTxLcdlSeed value 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'h1015f, value : 32'h62}, //[dwc_ddrphy_phyinit_programLCDLSeed] Pstate=0, Memclk=800MHz, Programming RDqRDqsCntrl to 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'h1115f, value : 32'h62}, //phyinit_io_write: 0x1015f, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'h1215f, value : 32'h62}, //phyinit_io_write: 0x1115f, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'h1315f, value : 32'h62}, //phyinit_io_write: 0x1215f, 0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'h60009, value : 32'h10}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Memclk=800MHz, Programming CPllDacValIn to 0x10
                          '{ step_type : REG_WRITE, reg_addr : 32'h102a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE0.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h102a1, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE0.RxReplicaPathPhase1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h102a2, value : 32'ha}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE0.RxReplicaPathPhase2 to 0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h102a3, value : 32'h3e}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE0.RxReplicaPathPhase3 to 0x3e
                          '{ step_type : REG_WRITE, reg_addr : 32'h102a4, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE0.RxReplicaPathPhase4 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h112a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE1.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h112a1, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE1.RxReplicaPathPhase1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h112a2, value : 32'ha}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE1.RxReplicaPathPhase2 to 0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h112a3, value : 32'h3e}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE1.RxReplicaPathPhase3 to 0x3e
                          '{ step_type : REG_WRITE, reg_addr : 32'h112a4, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE1.RxReplicaPathPhase4 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h122a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE2.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h122a1, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE2.RxReplicaPathPhase1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h122a2, value : 32'ha}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE2.RxReplicaPathPhase2 to 0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h122a3, value : 32'h3e}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE2.RxReplicaPathPhase3 to 0x3e
                          '{ step_type : REG_WRITE, reg_addr : 32'h122a4, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE2.RxReplicaPathPhase4 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h132a0, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE3.RxReplicaPathPhase0 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h132a1, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE3.RxReplicaPathPhase1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h132a2, value : 32'ha}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE3.RxReplicaPathPhase2 to 0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h132a3, value : 32'h3e}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE3.RxReplicaPathPhase3 to 0x3e
                          '{ step_type : REG_WRITE, reg_addr : 32'h132a4, value : 32'h72}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE3.RxReplicaPathPhase4 to 0x72
                          '{ step_type : REG_WRITE, reg_addr : 32'h102ad, value : 32'h3}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE0.RxReplicaCtl01::RxReplicaSelPathPhase to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h112ad, value : 32'h3}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE1.RxReplicaCtl01::RxReplicaSelPathPhase to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h122ad, value : 32'h3}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE2.RxReplicaCtl01::RxReplicaSelPathPhase to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h132ad, value : 32'h3}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE3.RxReplicaCtl01::RxReplicaSelPathPhase to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h102af, value : 32'h4c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE0.RxReplicaCtl03 to 0x4c
                          '{ step_type : REG_WRITE, reg_addr : 32'h112af, value : 32'h4c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE1.RxReplicaCtl03 to 0x4c
                          '{ step_type : REG_WRITE, reg_addr : 32'h122af, value : 32'h4c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE2.RxReplicaCtl03 to 0x4c
                          '{ step_type : REG_WRITE, reg_addr : 32'h132af, value : 32'h4c}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming DBYTE3.RxReplicaCtl03 to 0x4c
                          '{ step_type : REG_WRITE, reg_addr : 32'h90807, value : 32'h9701}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming Seq0BGPR7 to save ZQCalCodeOvrValPU=0x12e and ZQCalCodeOvrEnPU=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h90808, value : 32'hb681}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Pstate=0, Programming Seq0BGPR8 to save ZQCalCodeOvrValPD=0x16d and ZQCalCodeOvrEnPD=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1003f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1103f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1203f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h1}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h1303f, value : 32'h0}, //[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] Programming TtcfControl[TtcfForceSendAll] to 0x0
//[dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop] End of dwc_ddrphy_phyinit_progCsrSkipTrainPsLoop(), PState=0
// [dwc_ddrphy_phyinit_userCustom_E_setDfiClk] Start of dwc_ddrphy_phyinit_userCustom_E_setDfiClk()
// [dwc_ddrphy_phyinit_userCustom_E_setDfiClk] End of dwc_ddrphy_phyinit_userCustom_E_setDfiClk()
// [dwc_ddrphy_phyinit_F_loadDMEM1D] Start of dwc_ddrphy_phyinit_F_loadDMEM (pstate=0, Train2D=0)
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0088, value : 32'h1}, //[dwc_ddrphy_phyinit_F_loadDMEM] Program csr StartDccmClear to 1 to clear DCCM.
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 8300},
//Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 8300 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0088, value : 32'h0}, //[dwc_ddrphy_phyinit_F_loadDMEM] Program csr StartDccmClear to 0 after DCCM clear is done.
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}, //Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 40 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'h58000, value : 32'h600}, // [dwc_ddrphy_phyinit_WriteOutMem] STARTING. offset 0x58000 size 0x6000, sparse_write=1
                          '{ step_type : REG_WRITE, reg_addr : 32'h58001, value : 32'h19000020},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58002, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58004, value : 32'hff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58005, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58009, value : 32'h310},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5800f, value : 32'h10000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58010, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58016, value : 32'hb0b00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58017, value : 32'hbbbbb0b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58018, value : 32'he0ebbbb},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58019, value : 32'h54540e0e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801a, value : 32'h44445454},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801b, value : 32'h50504444},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801c, value : 32'h5050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801d, value : 32'h50500000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801e, value : 32'h50505050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5801f, value : 32'h5050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58020, value : 32'hac840000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58021, value : 32'hac84},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58023, value : 32'h2020000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58024, value : 32'h202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5802a, value : 32'h4040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5802b, value : 32'h404},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58032, value : 32'h60600000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58033, value : 32'h6060},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58048, value : 32'h3b000001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58049, value : 32'h37},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58054, value : 32'h5c0032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58055, value : 32'he000b6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58056, value : 32'h164013a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58057, value : 32'h1e801be},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58062, value : 32'h6400c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58103, value : 32'h50b0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58104, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58108, value : 32'h8080808},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58110, value : 32'hef0f4f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811b, value : 32'h4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811d, value : 32'h40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811e, value : 32'h180f0e0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5811f, value : 32'h4746451e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58120, value : 32'h4a4948},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58121, value : 32'h1000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58125, value : 32'h40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58126, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58129, value : 32'hffffffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5812e, value : 32'h2f059},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5812f, value : 32'hffb50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58130, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58131, value : 32'h1f0b5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58132, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58133, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58134, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58135, value : 32'hf0b00000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58136, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58137, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58138, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58139, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813a, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813b, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813c, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813d, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813e, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5813f, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58140, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58141, value : 32'hff740182},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58142, value : 32'h800001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58143, value : 32'h1ffbe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58144, value : 32'hf0be0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58145, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58146, value : 32'h1f0a7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58147, value : 32'hf0a20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58148, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58149, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814a, value : 32'h40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814b, value : 32'h308},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814c, value : 32'h560},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814e, value : 32'h80000dbc},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5814f, value : 32'h309},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58150, value : 32'h561},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58151, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58152, value : 32'h80000dcd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58153, value : 32'he0305},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58154, value : 32'he0205},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58155, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58156, value : 32'h80000dde},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58157, value : 32'he0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58158, value : 32'he0200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58159, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815a, value : 32'h80000e44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815b, value : 32'he0301},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815c, value : 32'he0201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815d, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815e, value : 32'h80000e57},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5815f, value : 32'he0302},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58160, value : 32'he0202},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58161, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58162, value : 32'h80000e6a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58163, value : 32'he0303},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58164, value : 32'he0203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58165, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58166, value : 32'h80000e7d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58167, value : 32'he0304},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58168, value : 32'he0204},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58169, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816a, value : 32'h80000e90},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816b, value : 32'h1ff01ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816c, value : 32'he0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816e, value : 32'h63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5816f, value : 32'h64},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58170, value : 32'h660},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58172, value : 32'h80000d8f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58173, value : 32'h661},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58174, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58175, value : 32'h80000dad},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58176, value : 32'he00f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58177, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58178, value : 32'h80000def},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58179, value : 32'he00f1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817a, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817b, value : 32'h80000e00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817c, value : 32'he00f2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817d, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817e, value : 32'h80000e11},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5817f, value : 32'he00f3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58180, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58181, value : 32'h80000e22},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58182, value : 32'he00f4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58183, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58184, value : 32'h80000e33},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58185, value : 32'he00f5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58186, value : 32'h3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58187, value : 32'h80000d9e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58188, value : 32'h2011210},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58189, value : 32'h1c0a1403},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818a, value : 32'hb112e29},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818b, value : 32'h1916150d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818c, value : 32'h180f0e0c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818d, value : 32'h453a131e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818e, value : 32'h49484746},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5818f, value : 32'h2006e4a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58190, value : 32'h100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58191, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58192, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58194, value : 32'h2150001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58195, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58196, value : 32'h1010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58197, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58198, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58199, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819a, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819b, value : 32'h6400002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819c, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819d, value : 32'h30215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819e, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5819f, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a0, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a1, value : 32'h10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a2, value : 32'habe0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a3, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a4, value : 32'h50320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581a5, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c5, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c6, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c7, value : 32'h43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c8, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581c9, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ca, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cb, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cc, value : 32'h42b0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cd, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ce, value : 32'h200c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581cf, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d0, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d1, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d2, value : 32'h10003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d3, value : 32'h8550002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d4, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d5, value : 32'h40158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d6, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d7, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d8, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581d9, value : 32'h10005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581da, value : 32'hc800002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581db, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581dc, value : 32'h601d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581dd, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581de, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581df, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e0, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e1, value : 32'h10ab0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e2, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e3, value : 32'h80258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e4, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e5, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e6, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e7, value : 32'h20009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e8, value : 32'h157c0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581e9, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ea, value : 32'ha02ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581eb, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ec, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ed, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ee, value : 32'h2000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ef, value : 32'h19000004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f0, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f1, value : 32'hc03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f2, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f3, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f4, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f5, value : 32'h3000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f6, value : 32'h21550006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f7, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f8, value : 32'he04b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581f9, value : 32'h70003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fa, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fb, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fc, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fd, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581fe, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h581ff, value : 32'h2150004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58200, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58201, value : 32'h4010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58202, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58203, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58204, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58205, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58206, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58207, value : 32'h80006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58208, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58209, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820a, value : 32'h6400006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820b, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820c, value : 32'h80215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820d, value : 32'h2000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820e, value : 32'h30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5820f, value : 32'h70004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58210, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58211, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58212, value : 32'he0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58213, value : 32'h70001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58214, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58215, value : 32'habe0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58216, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58217, value : 32'ha0320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58218, value : 32'h30010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58219, value : 32'h40009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5821a, value : 32'h80004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824c, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824d, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824e, value : 32'h20043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5824f, value : 32'h2},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58250, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58251, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58252, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58253, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58254, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58255, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58256, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58257, value : 32'h42b0003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58258, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58259, value : 32'h300c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825a, value : 32'h10004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825b, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825c, value : 32'h30002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825d, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825e, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5825f, value : 32'h50004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58260, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58261, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58262, value : 32'h8550004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58263, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58264, value : 32'h40158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58265, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58266, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58267, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58268, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58269, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826a, value : 32'h80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826b, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826c, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826d, value : 32'hc800004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826e, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5826f, value : 32'h601d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58270, value : 32'h20009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58271, value : 32'h30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58272, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58273, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58274, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58275, value : 32'hb0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58276, value : 32'h70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58277, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58278, value : 32'h10ab0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58279, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827a, value : 32'h70258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827b, value : 32'h3000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827c, value : 32'h30008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827d, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827e, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5827f, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58280, value : 32'he0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58281, value : 32'h90003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58282, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58283, value : 32'h157c0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58284, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58285, value : 32'h902ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58286, value : 32'h4000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58287, value : 32'h4000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58288, value : 32'h60002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58289, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828a, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828b, value : 32'h100009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828c, value : 32'hb0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828d, value : 32'h20004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828e, value : 32'h19000006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5828f, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58290, value : 32'hb03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58291, value : 32'h50013},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58292, value : 32'h5000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58293, value : 32'h70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58294, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58295, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58296, value : 32'h16000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58297, value : 32'hf0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58298, value : 32'h20006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58299, value : 32'h21550008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829a, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829b, value : 32'he04b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829c, value : 32'h60018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829d, value : 32'h70010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829e, value : 32'h90002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5829f, value : 32'h2150028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a0, value : 32'h85000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a1, value : 32'h60006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a2, value : 32'h6},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a4, value : 32'h60001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a5, value : 32'h2150007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a6, value : 32'h85042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a7, value : 32'h8010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582a8, value : 32'h80008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582aa, value : 32'h20000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ab, value : 32'h90007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ac, value : 32'h640042b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ad, value : 32'h190010b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ae, value : 32'ha000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582af, value : 32'h1000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b0, value : 32'h30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b1, value : 32'h80002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b2, value : 32'h640000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b3, value : 32'h1900855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b4, value : 32'hc0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b5, value : 32'he000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b6, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b7, value : 32'h30004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b8, value : 32'hb0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582b9, value : 32'habe0855},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582ba, value : 32'h2b00215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bb, value : 32'h100010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bc, value : 32'h30012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bd, value : 32'h50003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582be, value : 32'ha0004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582bf, value : 32'habe000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c0, value : 32'h2b00c80},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c1, value : 32'h120320},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c2, value : 32'h140014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c3, value : 32'h70005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c4, value : 32'h40007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h582c5, value : 32'he000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58300, value : 32'h280000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58301, value : 32'h50215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58302, value : 32'h30043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58303, value : 32'h30003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58305, value : 32'h10000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58306, value : 32'h40003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58307, value : 32'h42b0215},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58308, value : 32'h850043},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58309, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830a, value : 32'h4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830c, value : 32'h40001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830d, value : 32'h42b0005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830e, value : 32'h850640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5830f, value : 32'h500c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58310, value : 32'h50005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58311, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58312, value : 32'h10002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58313, value : 32'h50004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58314, value : 32'h8550640},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58315, value : 32'h10b00c8},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58316, value : 32'h70006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58317, value : 32'h10007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58318, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58319, value : 32'h40002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831a, value : 32'h8550006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831b, value : 32'h10b0abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831c, value : 32'h80158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831d, value : 32'h90008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831e, value : 32'h20002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5831f, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58320, value : 32'h70005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58321, value : 32'hc800abe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58322, value : 32'h1900158},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58323, value : 32'ha0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58324, value : 32'h3000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58325, value : 32'h40004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58326, value : 32'h50002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58327, value : 32'hc800007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58328, value : 32'h1900e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58329, value : 32'ha01d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832a, value : 32'hc000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832b, value : 32'h40003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832c, value : 32'h30005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832d, value : 32'h80005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832e, value : 32'h10ab0e95},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5832f, value : 32'h21501d3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58330, value : 32'hd000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58331, value : 32'h4000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58332, value : 32'h60005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58333, value : 32'h60003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58334, value : 32'h10ab0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58335, value : 32'h21512c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58336, value : 32'hd0258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58337, value : 32'hf000e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58338, value : 32'h60005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58339, value : 32'h30007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833a, value : 32'h90006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833b, value : 32'h157c12c0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833c, value : 32'h2b00258},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833d, value : 32'h10000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833e, value : 32'h60011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5833f, value : 32'h80007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58340, value : 32'h60004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58341, value : 32'h157c000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58342, value : 32'h2b01770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58343, value : 32'h1002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58344, value : 32'h130011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58345, value : 32'h70006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58346, value : 32'h40009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58347, value : 32'hb0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58348, value : 32'h19001770},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58349, value : 32'h32002ee},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834a, value : 32'h120011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834b, value : 32'h70014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834c, value : 32'ha0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834d, value : 32'h70004},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834e, value : 32'h1900000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5834f, value : 32'h3201d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58350, value : 32'h1403aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58351, value : 32'h180016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58352, value : 32'h90007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58353, value : 32'h5000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58354, value : 32'he0009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58355, value : 32'h21551d4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58356, value : 32'h42b03aa},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58357, value : 32'h190017},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58358, value : 32'h8001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58359, value : 32'hb000a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835a, value : 32'ha0006},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835b, value : 32'h21550010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835c, value : 32'h42b2580},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835d, value : 32'h1904b0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835e, value : 32'h1d001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5835f, value : 32'hb0008},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58360, value : 32'h7000c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58361, value : 32'h12000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58362, value : 32'ha05},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58363, value : 32'h50000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58364, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58365, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58366, value : 32'h43416564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58367, value : 32'h63500030},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58368, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58369, value : 32'h646f4341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836a, value : 32'h53514465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836b, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836c, value : 32'h4143446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836d, value : 32'h65646f43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836e, value : 32'h314341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5836f, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58370, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58371, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58372, value : 32'h30434174},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58373, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58374, value : 32'h4443446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58375, value : 32'h7366664f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58376, value : 32'h43417465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58377, value : 32'h63500031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58378, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58379, value : 32'h66664f44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837a, value : 32'h44746573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837b, value : 32'h50005351},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837c, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837d, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837e, value : 32'h71446564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5837f, value : 32'h306e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58380, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58381, value : 32'h43414344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58382, value : 32'h4465646f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58383, value : 32'h316e4c71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58384, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58385, value : 32'h4143446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58386, value : 32'h65646f43},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58387, value : 32'h6e4c7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58388, value : 32'h63500032},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58389, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838a, value : 32'h646f4341},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838b, value : 32'h4c714465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838c, value : 32'h5000336e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838d, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838e, value : 32'h6f434143},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5838f, value : 32'h71446564},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58390, value : 32'h346e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58391, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58392, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58393, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58394, value : 32'h4c714474},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58395, value : 32'h5000306e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58396, value : 32'h446b6c63},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58397, value : 32'h664f4443},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58398, value : 32'h74657366},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58399, value : 32'h6e4c7144},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839a, value : 32'h63500031},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839b, value : 32'h43446b6c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839c, value : 32'h66664f44},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839d, value : 32'h44746573},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839e, value : 32'h326e4c71},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5839f, value : 32'h6c635000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a0, value : 32'h4443446b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a1, value : 32'h7366664f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a2, value : 32'h71447465},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a3, value : 32'h336e4c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a4, value : 32'h6b6c6350},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a5, value : 32'h4f444344},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a6, value : 32'h65736666},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a7, value : 32'h4c714474},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a8, value : 32'h346e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583a9, value : 32'h4050607},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583aa, value : 32'h10203},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ab, value : 32'hc0b0a09},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ac, value : 32'hb50f0e0d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ad, value : 32'h1ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ae, value : 32'h1f0b500},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583af, value : 32'hb3000100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b0, value : 32'h1f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b1, value : 32'h1f0b400},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b2, value : 32'hb0000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b3, value : 32'h300001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b4, value : 32'h7f00300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b5, value : 32'h4000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b6, value : 32'h7f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b7, value : 32'h1fe0300},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b8, value : 32'h4000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583b9, value : 32'h1fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ba, value : 32'h7f01100},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bb, value : 32'h21000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bc, value : 32'h1fe},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bd, value : 32'h1ffbe00},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583be, value : 32'hbe000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583bf, value : 32'h10001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c0, value : 32'h1f0a700},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c1, value : 32'ha2000000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c2, value : 32'h20001f0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c3, value : 32'h2007900},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c4, value : 32'h4000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c5, value : 32'h1008b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c6, value : 32'hf05f0000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c7, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c8, value : 32'h1ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583c9, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ca, value : 32'h1ff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cb, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cc, value : 32'hf0b001ff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cd, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ce, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583cf, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d0, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d1, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d2, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d3, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d4, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d5, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d6, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d7, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d8, value : 32'hf0a70002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583d9, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583da, value : 32'he000f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583db, value : 32'hc000d},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583dc, value : 32'ha000b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583dd, value : 32'h80009},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583de, value : 32'h60007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583df, value : 32'h40005},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e0, value : 32'h20003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e1, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e2, value : 32'h110010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e3, value : 32'h130012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e4, value : 32'h150014},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e5, value : 32'h170016},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e6, value : 32'h190018},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e7, value : 32'h1b001a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e8, value : 32'h1d001c},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583e9, value : 32'h1f001e},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ea, value : 32'hef77dbb7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583eb, value : 32'hfbdff7bd},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ec, value : 32'hbddfb76f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ed, value : 32'hbdffbdef},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ee, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ef, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f0, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f1, value : 32'h200},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f2, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f3, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f4, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f5, value : 32'h10},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f6, value : 32'h1ffb5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f7, value : 32'hf0b30001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f8, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583f9, value : 32'h1f0b4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fa, value : 32'hf0b90000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fb, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fc, value : 32'h1f0ba},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fd, value : 32'hf0b10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583fe, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h583ff, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58400, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58401, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58402, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58403, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58404, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58405, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58406, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58407, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58408, value : 32'h7f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58409, value : 32'hfe200002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840a, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840b, value : 32'h7f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840c, value : 32'hf01cffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840d, value : 32'hffff0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840e, value : 32'h1fe2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5840f, value : 32'hfe2bffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58410, value : 32'hffff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58411, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58412, value : 32'hffb50040},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58413, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58414, value : 32'h1f0b3},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58415, value : 32'hf0b40000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58416, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58417, value : 32'h1f0b9},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58418, value : 32'hf0ba0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58419, value : 32'h10001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841a, value : 32'h1f0b1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841b, value : 32'hf0b00002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841c, value : 32'h300001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841d, value : 32'h7f003},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841e, value : 32'hf0040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5841f, value : 32'h7},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58420, value : 32'h1fe03},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58421, value : 32'hfe040000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58422, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58423, value : 32'h7f011},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58424, value : 32'hfe210000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58425, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58426, value : 32'h7f010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58427, value : 32'hfe200002},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58428, value : 32'h20001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58429, value : 32'h7f01b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842a, value : 32'hf01cffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842b, value : 32'hffff0007},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842c, value : 32'h1fe2a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842d, value : 32'hfe2bffff},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842e, value : 32'hffff0001},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5842f, value : 32'h20079},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58430, value : 32'h40},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58431, value : 32'h8840884},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58432, value : 32'h20},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58433, value : 32'h10010},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58434, value : 32'h10012},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58435, value : 32'h1007a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58436, value : 32'h10028},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58437, value : 32'h60000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58438, value : 32'h50005000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58439, value : 32'h2008050},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843b, value : 32'h60080},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843c, value : 32'h3c5a5555},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5843d, value : 32'h600000},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58440, value : 32'h70},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58441, value : 32'h75},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58442, value : 32'h26},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58443, value : 32'ha0},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58444, value : 32'ha1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58445, value : 32'ha4},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58446, value : 32'ha5},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58447, value : 32'ha030201},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58448, value : 32'he0d0c0b},
                          '{ step_type : REG_WRITE, reg_addr : 32'h58449, value : 32'h1413120f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844a, value : 32'h18171615},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844b, value : 32'h1e1c1a19},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844c, value : 32'h2221201f},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844d, value : 32'h2e292825},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844e, value : 32'h4746453a},
                          '{ step_type : REG_WRITE, reg_addr : 32'h5844f, value : 32'h4a4948},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1}, //This allows the firmware unrestricted access to the configuration CSRs.
//[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
// [dwc_ddrphy_phyinit_F_loadDMEM1D] End of dwc_ddrphy_phyinit_F_loadDMEM, Pstate=0
// [dwc_ddrphy_phyinit_G_execFW] Start of dwc_ddrphy_phyinit_G_execFW
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1}, ////     Then rewrite the CSR so that only the StallToMicro remains set (all other fields should be zero).
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h9}, //[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h0}, // [dwc_ddrphy_phyinit_userCustom_G_waitFwDone] Start of dwc_ddrphy_phyinit_userCustom_G_waitFwDone()
// [dwc_ddrphy_phyinit_userCustom_G_waitFwDone] End of dwc_ddrphy_phyinit_userCustom_G_waitFwDone()
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0099, value : 32'h1}, //// 4.   Halt the microcontroller."
// [dwc_ddrphy_phyinit_G_execFW] End of dwc_ddrphy_phyinit_G_execFW
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}, // [dwc_ddrphy_phyinit_userCustom_H_readMsgBlock] Start of dwc_ddrphy_phyinit_userCustom_H_readMsgBlock()
// [dwc_ddrphy_phyinit_userCustom_H_readMsgBlock] End of dwc_ddrphy_phyinit_userCustom_H_readMsgBlock ()
// 3. If training is required at another frequency, repeat the operations starting at step (E).
// [dwc_ddrphy_phyinit_H_readMsgBlock] End of dwc_ddrphy_phyinit_H_readMsgBlock
//[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Start of dwc_ddrphy_phyinit_I_loadPIEImagePsLoop(), PState=0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb0310, value : 32'h1}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming ZCalRun to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'hb0311, value : 32'h1},
                          '{ step_type : REG_WRITE, reg_addr : 32'h60008, value : 32'h2d56}, //[dwc_ddrphy_phyinit_programPLL] [phyinit_I_loadPIEImagePsLoop] Pstate=0,  Memclk=800MHz, Programming CpllCtrl5 to 0x2d56.
                          '{ step_type : REG_WRITE, reg_addr : 32'h60006, value : 32'h3f0}, //End of dwc_ddrphy_phyinit_programPLL(), PState=0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30015, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31015, value : 32'h0}, //phyinit_io_write: 0x30015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1007c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1107c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1207c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1307c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming SingleEndedMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1007c, value : 32'h0}, //phyinit_io_write: 0x1307c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1107c, value : 32'h0}, //phyinit_io_write: 0x1007c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1207c, value : 32'h0}, //phyinit_io_write: 0x1107c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1307c, value : 32'h0}, //phyinit_io_write: 0x1207c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h30015, value : 32'h0}, //phyinit_io_write: 0x1307c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h31015, value : 32'h0}, //phyinit_io_write: 0x30015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70141, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming ACSMWckFreeRunMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hb0001, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming ZcalClkDiv to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h9080c, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming GPR12 with Zcalkclkdiv to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h10027, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming RxClkCntl1 to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h11027, value : 32'h0}, //phyinit_io_write: 0x10027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h12027, value : 32'h0}, //phyinit_io_write: 0x11027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h13027, value : 32'h0}, //phyinit_io_write: 0x12027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h1020f, value : 32'h8}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Pstate=0, Programming RxReplicaCtl04 to 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h1120f, value : 32'h8}, //phyinit_io_write: 0x1020f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h1220f, value : 32'h8}, //phyinit_io_write: 0x1120f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h1320f, value : 32'h8}, //phyinit_io_write: 0x1220f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'he003f, value : 32'h1}, //phyinit_io_write: 0x1320f, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'he008d, value : 32'h1}, //phyinit_io_write: 0xe003f, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he103f, value : 32'h1}, //phyinit_io_write: 0xe008d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he108d, value : 32'h1}, //phyinit_io_write: 0xe103f, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he203f, value : 32'h1}, //phyinit_io_write: 0xe108d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he208d, value : 32'h1}, //phyinit_io_write: 0xe203f, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he303f, value : 32'h1}, //phyinit_io_write: 0xe208d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he308d, value : 32'h1}, //phyinit_io_write: 0xe303f, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he403f, value : 32'h1}, //phyinit_io_write: 0xe308d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he408d, value : 32'h1}, //phyinit_io_write: 0xe403f, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he503f, value : 32'h1}, //phyinit_io_write: 0xe408d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he508d, value : 32'h1}, //phyinit_io_write: 0xe503f, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he603f, value : 32'h1}, //phyinit_io_write: 0xe508d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he608d, value : 32'h1}, //phyinit_io_write: 0xe603f, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he703f, value : 32'h1}, //phyinit_io_write: 0xe608d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'he708d, value : 32'h1}, //phyinit_io_write: 0xe703f, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h90903, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] PState=0, Programming RtrnMode to 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70072, value : 32'h3}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming HwtLpCsEnA to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h9080e, value : 32'h3}, //phyinit_io_write: 0x70072, 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h70073, value : 32'h3}, //[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] Programming HwtLpCsEnB to 0x3
                          '{ step_type : REG_WRITE, reg_addr : 32'h9080f, value : 32'h3}, //phyinit_io_write: 0x70073, 0x3
//phyinit_io_write: 0x9080f, 0x3
//[dwc_ddrphy_phyinit_I_loadPIEImagePsLoop] End of dwc_ddrphy_phyinit_I_loadPIEImagePsLoop(), PState=0
//[dwc_ddrphy_phyinit_userCustom_customPostTrainPsLoop] End of dwc_ddrphy_phyinit_userCustom_customPostTrainPsLoop(), PState=0
//[dwc_ddrphy_phyinit_I_loadPIEImage] Start of dwc_ddrphy_phyinit_I_loadPIEImage() prog_csr=1
                          '{ step_type : WAIT_DFI, reg_addr : 0, value : 40},
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h0}, //Calling  [dwc_ddrphy_phyinit_userCustom_wait] to wait 40 DfiClks;
                          '{ step_type : REG_WRITE, reg_addr : 32'h41000, value : 32'h0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41001, value : 32'h0}, //phyinit_io_write: 0x41000, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41002, value : 32'h0}, //phyinit_io_write: 0x41001, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41003, value : 32'h0}, //phyinit_io_write: 0x41002, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41454, value : 32'hc028}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 16
                          '{ step_type : REG_WRITE, reg_addr : 32'h41455, value : 32'h100000}, //phyinit_io_write: 0x41454, 0xc028
                          '{ step_type : REG_WRITE, reg_addr : 32'h41456, value : 32'h0}, //phyinit_io_write: 0x41455, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41457, value : 32'h0}, //phyinit_io_write: 0x41456, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41458, value : 32'h0}, //phyinit_io_write: 0x41457, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41459, value : 32'h4000000}, //phyinit_io_write: 0x41458, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4145a, value : 32'h0}, //phyinit_io_write: 0x41459, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4145b, value : 32'h0}, //phyinit_io_write: 0x4145a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4145c, value : 32'h0}, //phyinit_io_write: 0x4145b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4145d, value : 32'h0}, //phyinit_io_write: 0x4145c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4145e, value : 32'h0}, //phyinit_io_write: 0x4145d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4145f, value : 32'h0}, //phyinit_io_write: 0x4145e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41460, value : 32'hc858}, //phyinit_io_write: 0x4145f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41461, value : 32'h100000}, //phyinit_io_write: 0x41460, 0xc858
                          '{ step_type : REG_WRITE, reg_addr : 32'h41462, value : 32'he088}, //phyinit_io_write: 0x41461, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41463, value : 32'h100000}, //phyinit_io_write: 0x41462, 0xe088
                          '{ step_type : REG_WRITE, reg_addr : 32'h41464, value : 32'he038}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41465, value : 32'h100000}, //phyinit_io_write: 0x41464, 0xe038
                          '{ step_type : REG_WRITE, reg_addr : 32'h41466, value : 32'hc858}, //phyinit_io_write: 0x41465, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41467, value : 32'h100000}, //phyinit_io_write: 0x41466, 0xc858
                          '{ step_type : REG_WRITE, reg_addr : 32'h41468, value : 32'hc088}, //phyinit_io_write: 0x41467, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41469, value : 32'h100000}, //phyinit_io_write: 0x41468, 0xc088
                          '{ step_type : REG_WRITE, reg_addr : 32'h4146a, value : 32'h0}, //phyinit_io_write: 0x41469, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4146b, value : 32'h0}, //phyinit_io_write: 0x4146a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4146c, value : 32'hc028}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 16
                          '{ step_type : REG_WRITE, reg_addr : 32'h4146d, value : 32'h100000}, //phyinit_io_write: 0x4146c, 0xc028
                          '{ step_type : REG_WRITE, reg_addr : 32'h4146e, value : 32'h0}, //phyinit_io_write: 0x4146d, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4146f, value : 32'h0}, //phyinit_io_write: 0x4146e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41470, value : 32'h0}, //phyinit_io_write: 0x4146f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41471, value : 32'h4000000}, //phyinit_io_write: 0x41470, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41472, value : 32'h0}, //phyinit_io_write: 0x41471, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41473, value : 32'h0}, //phyinit_io_write: 0x41472, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41474, value : 32'h0}, //phyinit_io_write: 0x41473, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41475, value : 32'h0}, //phyinit_io_write: 0x41474, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41476, value : 32'h0}, //phyinit_io_write: 0x41475, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41477, value : 32'h0}, //phyinit_io_write: 0x41476, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41478, value : 32'hc858}, //phyinit_io_write: 0x41477, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41479, value : 32'h100000}, //phyinit_io_write: 0x41478, 0xc858
                          '{ step_type : REG_WRITE, reg_addr : 32'h4147a, value : 32'he208}, //phyinit_io_write: 0x41479, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4147b, value : 32'h100000}, //phyinit_io_write: 0x4147a, 0xe208
                          '{ step_type : REG_WRITE, reg_addr : 32'h4147c, value : 32'he038}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4147d, value : 32'h100000}, //phyinit_io_write: 0x4147c, 0xe038
                          '{ step_type : REG_WRITE, reg_addr : 32'h4147e, value : 32'hc858}, //phyinit_io_write: 0x4147d, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4147f, value : 32'h100000}, //phyinit_io_write: 0x4147e, 0xc858
                          '{ step_type : REG_WRITE, reg_addr : 32'h41480, value : 32'hc208}, //phyinit_io_write: 0x4147f, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41481, value : 32'h100000}, //phyinit_io_write: 0x41480, 0xc208
                          '{ step_type : REG_WRITE, reg_addr : 32'h41482, value : 32'h0}, //phyinit_io_write: 0x41481, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41483, value : 32'h0}, //phyinit_io_write: 0x41482, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41484, value : 32'hc040}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41485, value : 32'h100000}, //phyinit_io_write: 0x41484, 0xc040
                          '{ step_type : REG_WRITE, reg_addr : 32'h41486, value : 32'h0}, //phyinit_io_write: 0x41485, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41487, value : 32'h100000}, //phyinit_io_write: 0x41486, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41488, value : 32'hc068}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41489, value : 32'h100000}, //phyinit_io_write: 0x41488, 0xc068
                          '{ step_type : REG_WRITE, reg_addr : 32'h4148a, value : 32'h0}, //phyinit_io_write: 0x41489, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4148b, value : 32'h0}, //phyinit_io_write: 0x4148a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4148c, value : 32'hce58}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4148d, value : 32'h100000}, //phyinit_io_write: 0x4148c, 0xce58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4148e, value : 32'hc208}, //phyinit_io_write: 0x4148d, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4148f, value : 32'h100000}, //phyinit_io_write: 0x4148e, 0xc208
                          '{ step_type : REG_WRITE, reg_addr : 32'h41490, value : 32'h0}, //phyinit_io_write: 0x4148f, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41491, value : 32'h0}, //phyinit_io_write: 0x41490, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41492, value : 32'h0}, //phyinit_io_write: 0x41491, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41493, value : 32'h0}, //phyinit_io_write: 0x41492, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41494, value : 32'hc370}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41495, value : 32'h100000}, //phyinit_io_write: 0x41494, 0xc370
                          '{ step_type : REG_WRITE, reg_addr : 32'h41496, value : 32'h0}, //phyinit_io_write: 0x41495, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41497, value : 32'h0}, //phyinit_io_write: 0x41496, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41498, value : 32'hd2d8}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 100
                          '{ step_type : REG_WRITE, reg_addr : 32'h41499, value : 32'h100000}, //phyinit_io_write: 0x41498, 0xd2d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4149a, value : 32'he008}, //phyinit_io_write: 0x41499, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4149b, value : 32'h100000}, //phyinit_io_write: 0x4149a, 0xe008
                          '{ step_type : REG_WRITE, reg_addr : 32'h4149c, value : 32'h0}, //phyinit_io_write: 0x4149b, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4149d, value : 32'h7b000000}, //phyinit_io_write: 0x4149c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4149e, value : 32'h0}, //phyinit_io_write: 0x4149d, 0x7b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4149f, value : 32'h0}, //phyinit_io_write: 0x4149e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a0, value : 32'hc0f0}, //phyinit_io_write: 0x4149f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a1, value : 32'h100000}, //phyinit_io_write: 0x414a0, 0xc0f0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a2, value : 32'hcfd8}, //phyinit_io_write: 0x414a1, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a3, value : 32'h100000}, //phyinit_io_write: 0x414a2, 0xcfd8
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a4, value : 32'hc008}, //phyinit_io_write: 0x414a3, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a5, value : 32'h100000}, //phyinit_io_write: 0x414a4, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a6, value : 32'h0}, //phyinit_io_write: 0x414a5, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a7, value : 32'h0}, //phyinit_io_write: 0x414a6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a8, value : 32'h0}, //phyinit_io_write: 0x414a7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414a9, value : 32'h3b000000}, //phyinit_io_write: 0x414a8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414aa, value : 32'h0}, //phyinit_io_write: 0x414a9, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ab, value : 32'h0}, //phyinit_io_write: 0x414aa, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ac, value : 32'h0}, //phyinit_io_write: 0x414ab, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ad, value : 32'h0}, //phyinit_io_write: 0x414ac, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ae, value : 32'hd058}, //phyinit_io_write: 0x414ad, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414af, value : 32'h100000}, //phyinit_io_write: 0x414ae, 0xd058
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b0, value : 32'hc008}, //phyinit_io_write: 0x414af, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b1, value : 32'h100000}, //phyinit_io_write: 0x414b0, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b2, value : 32'h0}, //phyinit_io_write: 0x414b1, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b3, value : 32'h0}, //phyinit_io_write: 0x414b2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b4, value : 32'h0}, //phyinit_io_write: 0x414b3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b5, value : 32'h3b000000}, //phyinit_io_write: 0x414b4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b6, value : 32'h0}, //phyinit_io_write: 0x414b5, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b7, value : 32'h0}, //phyinit_io_write: 0x414b6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b8, value : 32'h0}, //phyinit_io_write: 0x414b7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414b9, value : 32'h0}, //phyinit_io_write: 0x414b8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ba, value : 32'hd0d8}, //phyinit_io_write: 0x414b9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414bb, value : 32'h100000}, //phyinit_io_write: 0x414ba, 0xd0d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h414bc, value : 32'hc088}, //phyinit_io_write: 0x414bb, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414bd, value : 32'h100000}, //phyinit_io_write: 0x414bc, 0xc088
                          '{ step_type : REG_WRITE, reg_addr : 32'h414be, value : 32'h0}, //phyinit_io_write: 0x414bd, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414bf, value : 32'h0}, //phyinit_io_write: 0x414be, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c0, value : 32'h0}, //phyinit_io_write: 0x414bf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c1, value : 32'h3b000000}, //phyinit_io_write: 0x414c0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c2, value : 32'h0}, //phyinit_io_write: 0x414c1, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c3, value : 32'h0}, //phyinit_io_write: 0x414c2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c4, value : 32'h0}, //phyinit_io_write: 0x414c3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c5, value : 32'h0}, //phyinit_io_write: 0x414c4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c6, value : 32'hd158}, //phyinit_io_write: 0x414c5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c7, value : 32'h100000}, //phyinit_io_write: 0x414c6, 0xd158
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c8, value : 32'hc008}, //phyinit_io_write: 0x414c7, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414c9, value : 32'h100000}, //phyinit_io_write: 0x414c8, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ca, value : 32'h0}, //phyinit_io_write: 0x414c9, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414cb, value : 32'h0}, //phyinit_io_write: 0x414ca, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414cc, value : 32'h0}, //phyinit_io_write: 0x414cb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414cd, value : 32'h6b000000}, //phyinit_io_write: 0x414cc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ce, value : 32'h0}, //phyinit_io_write: 0x414cd, 0x6b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414cf, value : 32'h0}, //phyinit_io_write: 0x414ce, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d0, value : 32'h0}, //phyinit_io_write: 0x414cf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d1, value : 32'h0}, //phyinit_io_write: 0x414d0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d2, value : 32'h0}, //phyinit_io_write: 0x414d1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d3, value : 32'h0}, //phyinit_io_write: 0x414d2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d4, value : 32'hd00402c}, //phyinit_io_write: 0x414d3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d5, value : 32'h4000001}, //phyinit_io_write: 0x414d4, 0xd00402c
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d6, value : 32'h8004050}, //phyinit_io_write: 0x414d5, 0x4000001
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d7, value : 32'h0}, //phyinit_io_write: 0x414d6, 0x8004050
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d8, value : 32'h0}, //phyinit_io_write: 0x414d7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414d9, value : 32'h4000000}, //phyinit_io_write: 0x414d8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414da, value : 32'h0}, //phyinit_io_write: 0x414d9, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414db, value : 32'h0}, //phyinit_io_write: 0x414da, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414dc, value : 32'h0}, //phyinit_io_write: 0x414db, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414dd, value : 32'h4000000}, //phyinit_io_write: 0x414dc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414de, value : 32'h8034050}, //phyinit_io_write: 0x414dd, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414df, value : 32'h0}, //phyinit_io_write: 0x414de, 0x8034050
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e0, value : 32'h0}, //phyinit_io_write: 0x414df, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e1, value : 32'h1f000000}, //phyinit_io_write: 0x414e0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e2, value : 32'h0}, //phyinit_io_write: 0x414e1, 0x1f000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e3, value : 32'h8000000}, //phyinit_io_write: 0x414e2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e4, value : 32'h0}, //phyinit_io_write: 0x414e3, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e5, value : 32'h4000000}, //phyinit_io_write: 0x414e4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e6, value : 32'h407c}, //phyinit_io_write: 0x414e5, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e7, value : 32'h0}, //phyinit_io_write: 0x414e6, 0x407c
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e8, value : 32'h0}, //phyinit_io_write: 0x414e7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414e9, value : 32'h4000000}, //phyinit_io_write: 0x414e8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ea, value : 32'h0}, //phyinit_io_write: 0x414e9, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414eb, value : 32'h0}, //phyinit_io_write: 0x414ea, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ec, value : 32'h0}, //phyinit_io_write: 0x414eb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ed, value : 32'h4000001}, //phyinit_io_write: 0x414ec, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ee, value : 32'h0}, //phyinit_io_write: 0x414ed, 0x4000001
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ef, value : 32'h0}, //phyinit_io_write: 0x414ee, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f0, value : 32'h0}, //phyinit_io_write: 0x414ef, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f1, value : 32'h4000000}, //phyinit_io_write: 0x414f0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f2, value : 32'h0}, //phyinit_io_write: 0x414f1, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f3, value : 32'h0}, //phyinit_io_write: 0x414f2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f4, value : 32'h0}, //phyinit_io_write: 0x414f3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f5, value : 32'h1b000000}, //phyinit_io_write: 0x414f4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f6, value : 32'h0}, //phyinit_io_write: 0x414f5, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f7, value : 32'h0}, //phyinit_io_write: 0x414f6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f8, value : 32'h0}, //phyinit_io_write: 0x414f7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414f9, value : 32'h0}, //phyinit_io_write: 0x414f8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414fa, value : 32'h0}, //phyinit_io_write: 0x414f9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414fb, value : 32'h0}, //phyinit_io_write: 0x414fa, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h414fc, value : 32'hd00802c}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 40
                          '{ step_type : REG_WRITE, reg_addr : 32'h414fd, value : 32'h4100001}, //phyinit_io_write: 0x414fc, 0xd00802c
                          '{ step_type : REG_WRITE, reg_addr : 32'h414fe, value : 32'h8008050}, //phyinit_io_write: 0x414fd, 0x4100001
                          '{ step_type : REG_WRITE, reg_addr : 32'h414ff, value : 32'h100000}, //phyinit_io_write: 0x414fe, 0x8008050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41500, value : 32'h0}, //phyinit_io_write: 0x414ff, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41501, value : 32'h4000000}, //phyinit_io_write: 0x41500, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41502, value : 32'h0}, //phyinit_io_write: 0x41501, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41503, value : 32'h0}, //phyinit_io_write: 0x41502, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41504, value : 32'h0}, //phyinit_io_write: 0x41503, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41505, value : 32'h4000000}, //phyinit_io_write: 0x41504, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41506, value : 32'h8038050}, //phyinit_io_write: 0x41505, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41507, value : 32'h100000}, //phyinit_io_write: 0x41506, 0x8038050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41508, value : 32'h0}, //phyinit_io_write: 0x41507, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41509, value : 32'h1f000000}, //phyinit_io_write: 0x41508, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4150a, value : 32'h0}, //phyinit_io_write: 0x41509, 0x1f000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4150b, value : 32'h8000000}, //phyinit_io_write: 0x4150a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4150c, value : 32'h0}, //phyinit_io_write: 0x4150b, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4150d, value : 32'h4000000}, //phyinit_io_write: 0x4150c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4150e, value : 32'h807c}, //phyinit_io_write: 0x4150d, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4150f, value : 32'h100000}, //phyinit_io_write: 0x4150e, 0x807c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41510, value : 32'h0}, //phyinit_io_write: 0x4150f, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41511, value : 32'h4000000}, //phyinit_io_write: 0x41510, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41512, value : 32'h0}, //phyinit_io_write: 0x41511, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41513, value : 32'h0}, //phyinit_io_write: 0x41512, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41514, value : 32'h0}, //phyinit_io_write: 0x41513, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41515, value : 32'h4000001}, //phyinit_io_write: 0x41514, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41516, value : 32'h0}, //phyinit_io_write: 0x41515, 0x4000001
                          '{ step_type : REG_WRITE, reg_addr : 32'h41517, value : 32'h0}, //phyinit_io_write: 0x41516, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41518, value : 32'h0}, //phyinit_io_write: 0x41517, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41519, value : 32'h4000000}, //phyinit_io_write: 0x41518, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4151a, value : 32'h0}, //phyinit_io_write: 0x41519, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4151b, value : 32'h0}, //phyinit_io_write: 0x4151a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4151c, value : 32'h0}, //phyinit_io_write: 0x4151b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4151d, value : 32'h1b000000}, //phyinit_io_write: 0x4151c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4151e, value : 32'h0}, //phyinit_io_write: 0x4151d, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4151f, value : 32'h0}, //phyinit_io_write: 0x4151e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41520, value : 32'h0}, //phyinit_io_write: 0x4151f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41521, value : 32'h0}, //phyinit_io_write: 0x41520, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41522, value : 32'h0}, //phyinit_io_write: 0x41521, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41523, value : 32'h0}, //phyinit_io_write: 0x41522, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41524, value : 32'hd00402c}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 96
                          '{ step_type : REG_WRITE, reg_addr : 32'h41525, value : 32'h1}, //phyinit_io_write: 0x41524, 0xd00402c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41526, value : 32'h8004050}, //phyinit_io_write: 0x41525, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h41527, value : 32'h0}, //phyinit_io_write: 0x41526, 0x8004050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41528, value : 32'h0}, //phyinit_io_write: 0x41527, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41529, value : 32'h0}, //phyinit_io_write: 0x41528, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4152a, value : 32'h0}, //phyinit_io_write: 0x41529, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4152b, value : 32'h0}, //phyinit_io_write: 0x4152a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4152c, value : 32'h0}, //phyinit_io_write: 0x4152b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4152d, value : 32'h0}, //phyinit_io_write: 0x4152c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4152e, value : 32'h8034050}, //phyinit_io_write: 0x4152d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4152f, value : 32'h0}, //phyinit_io_write: 0x4152e, 0x8034050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41530, value : 32'h0}, //phyinit_io_write: 0x4152f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41531, value : 32'h0}, //phyinit_io_write: 0x41530, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41532, value : 32'h0}, //phyinit_io_write: 0x41531, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41533, value : 32'h0}, //phyinit_io_write: 0x41532, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41534, value : 32'h0}, //phyinit_io_write: 0x41533, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41535, value : 32'h0}, //phyinit_io_write: 0x41534, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41536, value : 32'h8034050}, //phyinit_io_write: 0x41535, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41537, value : 32'h0}, //phyinit_io_write: 0x41536, 0x8034050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41538, value : 32'h0}, //phyinit_io_write: 0x41537, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41539, value : 32'h0}, //phyinit_io_write: 0x41538, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4153a, value : 32'h0}, //phyinit_io_write: 0x41539, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4153b, value : 32'h0}, //phyinit_io_write: 0x4153a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4153c, value : 32'h0}, //phyinit_io_write: 0x4153b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4153d, value : 32'h0}, //phyinit_io_write: 0x4153c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4153e, value : 32'h8004050}, //phyinit_io_write: 0x4153d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4153f, value : 32'h0}, //phyinit_io_write: 0x4153e, 0x8004050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41540, value : 32'h0}, //phyinit_io_write: 0x4153f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41541, value : 32'h1b000000}, //phyinit_io_write: 0x41540, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41542, value : 32'h0}, //phyinit_io_write: 0x41541, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41543, value : 32'h8000000}, //phyinit_io_write: 0x41542, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41544, value : 32'h0}, //phyinit_io_write: 0x41543, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41545, value : 32'h0}, //phyinit_io_write: 0x41544, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41546, value : 32'h407c}, //phyinit_io_write: 0x41545, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41547, value : 32'h0}, //phyinit_io_write: 0x41546, 0x407c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41548, value : 32'h0}, //phyinit_io_write: 0x41547, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41549, value : 32'h0}, //phyinit_io_write: 0x41548, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4154a, value : 32'h0}, //phyinit_io_write: 0x41549, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4154b, value : 32'h0}, //phyinit_io_write: 0x4154a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4154c, value : 32'h0}, //phyinit_io_write: 0x4154b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4154d, value : 32'h1}, //phyinit_io_write: 0x4154c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4154e, value : 32'h0}, //phyinit_io_write: 0x4154d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4154f, value : 32'h0}, //phyinit_io_write: 0x4154e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41550, value : 32'h0}, //phyinit_io_write: 0x4154f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41551, value : 32'h5b000000}, //phyinit_io_write: 0x41550, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41552, value : 32'h0}, //phyinit_io_write: 0x41551, 0x5b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41553, value : 32'h1c000000}, //phyinit_io_write: 0x41552, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41554, value : 32'hd00802c}, //phyinit_io_write: 0x41553, 0x1c000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41555, value : 32'h100001}, //phyinit_io_write: 0x41554, 0xd00802c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41556, value : 32'h8008050}, //phyinit_io_write: 0x41555, 0x100001
                          '{ step_type : REG_WRITE, reg_addr : 32'h41557, value : 32'h100000}, //phyinit_io_write: 0x41556, 0x8008050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41558, value : 32'h0}, //phyinit_io_write: 0x41557, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41559, value : 32'h0}, //phyinit_io_write: 0x41558, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4155a, value : 32'h0}, //phyinit_io_write: 0x41559, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4155b, value : 32'h0}, //phyinit_io_write: 0x4155a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4155c, value : 32'h0}, //phyinit_io_write: 0x4155b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4155d, value : 32'h0}, //phyinit_io_write: 0x4155c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4155e, value : 32'h8038050}, //phyinit_io_write: 0x4155d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4155f, value : 32'h100000}, //phyinit_io_write: 0x4155e, 0x8038050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41560, value : 32'h0}, //phyinit_io_write: 0x4155f, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41561, value : 32'h0}, //phyinit_io_write: 0x41560, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41562, value : 32'h0}, //phyinit_io_write: 0x41561, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41563, value : 32'h0}, //phyinit_io_write: 0x41562, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41564, value : 32'h0}, //phyinit_io_write: 0x41563, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41565, value : 32'h0}, //phyinit_io_write: 0x41564, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41566, value : 32'h8038050}, //phyinit_io_write: 0x41565, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41567, value : 32'h100000}, //phyinit_io_write: 0x41566, 0x8038050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41568, value : 32'h0}, //phyinit_io_write: 0x41567, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41569, value : 32'h0}, //phyinit_io_write: 0x41568, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4156a, value : 32'h0}, //phyinit_io_write: 0x41569, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4156b, value : 32'h0}, //phyinit_io_write: 0x4156a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4156c, value : 32'h0}, //phyinit_io_write: 0x4156b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4156d, value : 32'h0}, //phyinit_io_write: 0x4156c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4156e, value : 32'h8008050}, //phyinit_io_write: 0x4156d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4156f, value : 32'h100000}, //phyinit_io_write: 0x4156e, 0x8008050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41570, value : 32'h0}, //phyinit_io_write: 0x4156f, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41571, value : 32'h1b000000}, //phyinit_io_write: 0x41570, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41572, value : 32'h0}, //phyinit_io_write: 0x41571, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41573, value : 32'h8000000}, //phyinit_io_write: 0x41572, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41574, value : 32'h0}, //phyinit_io_write: 0x41573, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41575, value : 32'h0}, //phyinit_io_write: 0x41574, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41576, value : 32'h807c}, //phyinit_io_write: 0x41575, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41577, value : 32'h100000}, //phyinit_io_write: 0x41576, 0x807c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41578, value : 32'h0}, //phyinit_io_write: 0x41577, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41579, value : 32'h0}, //phyinit_io_write: 0x41578, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4157a, value : 32'h0}, //phyinit_io_write: 0x41579, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4157b, value : 32'h0}, //phyinit_io_write: 0x4157a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4157c, value : 32'h0}, //phyinit_io_write: 0x4157b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4157d, value : 32'h1}, //phyinit_io_write: 0x4157c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4157e, value : 32'h0}, //phyinit_io_write: 0x4157d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4157f, value : 32'h0}, //phyinit_io_write: 0x4157e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41580, value : 32'h0}, //phyinit_io_write: 0x4157f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41581, value : 32'h4b000000}, //phyinit_io_write: 0x41580, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41582, value : 32'h0}, //phyinit_io_write: 0x41581, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41583, value : 32'h28000000}, //phyinit_io_write: 0x41582, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41584, value : 32'hd00402c}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 64
                          '{ step_type : REG_WRITE, reg_addr : 32'h41585, value : 32'h1}, //phyinit_io_write: 0x41584, 0xd00402c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41586, value : 32'h8035198}, //phyinit_io_write: 0x41585, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h41587, value : 32'h0}, //phyinit_io_write: 0x41586, 0x8035198
                          '{ step_type : REG_WRITE, reg_addr : 32'h41588, value : 32'h0}, //phyinit_io_write: 0x41587, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41589, value : 32'h2b000000}, //phyinit_io_write: 0x41588, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4158a, value : 32'h0}, //phyinit_io_write: 0x41589, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4158b, value : 32'h0}, //phyinit_io_write: 0x4158a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4158c, value : 32'h0}, //phyinit_io_write: 0x4158b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4158d, value : 32'h0}, //phyinit_io_write: 0x4158c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4158e, value : 32'h8035218}, //phyinit_io_write: 0x4158d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4158f, value : 32'h0}, //phyinit_io_write: 0x4158e, 0x8035218
                          '{ step_type : REG_WRITE, reg_addr : 32'h41590, value : 32'h0}, //phyinit_io_write: 0x4158f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41591, value : 32'h1b000000}, //phyinit_io_write: 0x41590, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41592, value : 32'h0}, //phyinit_io_write: 0x41591, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41593, value : 32'h8000000}, //phyinit_io_write: 0x41592, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41594, value : 32'h0}, //phyinit_io_write: 0x41593, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41595, value : 32'h0}, //phyinit_io_write: 0x41594, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41596, value : 32'h407c}, //phyinit_io_write: 0x41595, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41597, value : 32'h0}, //phyinit_io_write: 0x41596, 0x407c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41598, value : 32'h0}, //phyinit_io_write: 0x41597, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41599, value : 32'h0}, //phyinit_io_write: 0x41598, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4159a, value : 32'h0}, //phyinit_io_write: 0x41599, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4159b, value : 32'h0}, //phyinit_io_write: 0x4159a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4159c, value : 32'h0}, //phyinit_io_write: 0x4159b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4159d, value : 32'h1}, //phyinit_io_write: 0x4159c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4159e, value : 32'h0}, //phyinit_io_write: 0x4159d, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4159f, value : 32'h0}, //phyinit_io_write: 0x4159e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a0, value : 32'h0}, //phyinit_io_write: 0x4159f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a1, value : 32'h1b000000}, //phyinit_io_write: 0x415a0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a2, value : 32'h0}, //phyinit_io_write: 0x415a1, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a3, value : 32'h0}, //phyinit_io_write: 0x415a2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a4, value : 32'hd00802c}, //phyinit_io_write: 0x415a3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a5, value : 32'h100001}, //phyinit_io_write: 0x415a4, 0xd00802c
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a6, value : 32'h8039198}, //phyinit_io_write: 0x415a5, 0x100001
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a7, value : 32'h100000}, //phyinit_io_write: 0x415a6, 0x8039198
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a8, value : 32'h0}, //phyinit_io_write: 0x415a7, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415a9, value : 32'h2b000000}, //phyinit_io_write: 0x415a8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415aa, value : 32'h0}, //phyinit_io_write: 0x415a9, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ab, value : 32'h0}, //phyinit_io_write: 0x415aa, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ac, value : 32'h0}, //phyinit_io_write: 0x415ab, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ad, value : 32'h0}, //phyinit_io_write: 0x415ac, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ae, value : 32'h8039218}, //phyinit_io_write: 0x415ad, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415af, value : 32'h100000}, //phyinit_io_write: 0x415ae, 0x8039218
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b0, value : 32'h0}, //phyinit_io_write: 0x415af, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b1, value : 32'h1b000000}, //phyinit_io_write: 0x415b0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b2, value : 32'h0}, //phyinit_io_write: 0x415b1, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b3, value : 32'h8000000}, //phyinit_io_write: 0x415b2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b4, value : 32'h0}, //phyinit_io_write: 0x415b3, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b5, value : 32'h0}, //phyinit_io_write: 0x415b4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b6, value : 32'h807c}, //phyinit_io_write: 0x415b5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b7, value : 32'h100000}, //phyinit_io_write: 0x415b6, 0x807c
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b8, value : 32'h0}, //phyinit_io_write: 0x415b7, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415b9, value : 32'h0}, //phyinit_io_write: 0x415b8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ba, value : 32'h0}, //phyinit_io_write: 0x415b9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415bb, value : 32'h0}, //phyinit_io_write: 0x415ba, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415bc, value : 32'h0}, //phyinit_io_write: 0x415bb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415bd, value : 32'h1}, //phyinit_io_write: 0x415bc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415be, value : 32'h0}, //phyinit_io_write: 0x415bd, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h415bf, value : 32'h0}, //phyinit_io_write: 0x415be, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c0, value : 32'h0}, //phyinit_io_write: 0x415bf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c1, value : 32'h3b000000}, //phyinit_io_write: 0x415c0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c2, value : 32'h0}, //phyinit_io_write: 0x415c1, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c3, value : 32'h4000000}, //phyinit_io_write: 0x415c2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c4, value : 32'hd2d8}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 96
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c5, value : 32'h100000}, //phyinit_io_write: 0x415c4, 0xd2d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c6, value : 32'he008}, //phyinit_io_write: 0x415c5, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c7, value : 32'h100000}, //phyinit_io_write: 0x415c6, 0xe008
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c8, value : 32'h0}, //phyinit_io_write: 0x415c7, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415c9, value : 32'h7b000000}, //phyinit_io_write: 0x415c8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ca, value : 32'h0}, //phyinit_io_write: 0x415c9, 0x7b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415cb, value : 32'h0}, //phyinit_io_write: 0x415ca, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415cc, value : 32'hc0f0}, //phyinit_io_write: 0x415cb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415cd, value : 32'h100000}, //phyinit_io_write: 0x415cc, 0xc0f0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ce, value : 32'hcfd8}, //phyinit_io_write: 0x415cd, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415cf, value : 32'h100000}, //phyinit_io_write: 0x415ce, 0xcfd8
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d0, value : 32'hc008}, //phyinit_io_write: 0x415cf, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d1, value : 32'h100000}, //phyinit_io_write: 0x415d0, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d2, value : 32'h0}, //phyinit_io_write: 0x415d1, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d3, value : 32'h0}, //phyinit_io_write: 0x415d2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d4, value : 32'h0}, //phyinit_io_write: 0x415d3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d5, value : 32'h3b000000}, //phyinit_io_write: 0x415d4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d6, value : 32'h0}, //phyinit_io_write: 0x415d5, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d7, value : 32'h0}, //phyinit_io_write: 0x415d6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d8, value : 32'h0}, //phyinit_io_write: 0x415d7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415d9, value : 32'h0}, //phyinit_io_write: 0x415d8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415da, value : 32'hd058}, //phyinit_io_write: 0x415d9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415db, value : 32'h100000}, //phyinit_io_write: 0x415da, 0xd058
                          '{ step_type : REG_WRITE, reg_addr : 32'h415dc, value : 32'hc008}, //phyinit_io_write: 0x415db, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415dd, value : 32'h100000}, //phyinit_io_write: 0x415dc, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h415de, value : 32'h0}, //phyinit_io_write: 0x415dd, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415df, value : 32'h0}, //phyinit_io_write: 0x415de, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e0, value : 32'h0}, //phyinit_io_write: 0x415df, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e1, value : 32'h3b000000}, //phyinit_io_write: 0x415e0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e2, value : 32'h0}, //phyinit_io_write: 0x415e1, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e3, value : 32'h0}, //phyinit_io_write: 0x415e2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e4, value : 32'h0}, //phyinit_io_write: 0x415e3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e5, value : 32'h0}, //phyinit_io_write: 0x415e4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e6, value : 32'hd0d8}, //phyinit_io_write: 0x415e5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e7, value : 32'h100000}, //phyinit_io_write: 0x415e6, 0xd0d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e8, value : 32'hc088}, //phyinit_io_write: 0x415e7, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415e9, value : 32'h100000}, //phyinit_io_write: 0x415e8, 0xc088
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ea, value : 32'h0}, //phyinit_io_write: 0x415e9, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415eb, value : 32'h0}, //phyinit_io_write: 0x415ea, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ec, value : 32'h0}, //phyinit_io_write: 0x415eb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ed, value : 32'h3b000000}, //phyinit_io_write: 0x415ec, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ee, value : 32'h0}, //phyinit_io_write: 0x415ed, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ef, value : 32'h0}, //phyinit_io_write: 0x415ee, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f0, value : 32'h0}, //phyinit_io_write: 0x415ef, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f1, value : 32'h0}, //phyinit_io_write: 0x415f0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f2, value : 32'hd158}, //phyinit_io_write: 0x415f1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f3, value : 32'h100000}, //phyinit_io_write: 0x415f2, 0xd158
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f4, value : 32'hc008}, //phyinit_io_write: 0x415f3, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f5, value : 32'h100000}, //phyinit_io_write: 0x415f4, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f6, value : 32'h0}, //phyinit_io_write: 0x415f5, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f7, value : 32'h0}, //phyinit_io_write: 0x415f6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f8, value : 32'h0}, //phyinit_io_write: 0x415f7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415f9, value : 32'h6b000000}, //phyinit_io_write: 0x415f8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415fa, value : 32'h0}, //phyinit_io_write: 0x415f9, 0x6b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h415fb, value : 32'h0}, //phyinit_io_write: 0x415fa, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415fc, value : 32'h0}, //phyinit_io_write: 0x415fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415fd, value : 32'h0}, //phyinit_io_write: 0x415fc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415fe, value : 32'h0}, //phyinit_io_write: 0x415fd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h415ff, value : 32'h0}, //phyinit_io_write: 0x415fe, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41600, value : 32'hd00402c}, //phyinit_io_write: 0x415ff, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41601, value : 32'h4000001}, //phyinit_io_write: 0x41600, 0xd00402c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41602, value : 32'h8004050}, //phyinit_io_write: 0x41601, 0x4000001
                          '{ step_type : REG_WRITE, reg_addr : 32'h41603, value : 32'h0}, //phyinit_io_write: 0x41602, 0x8004050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41604, value : 32'h0}, //phyinit_io_write: 0x41603, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41605, value : 32'h4000000}, //phyinit_io_write: 0x41604, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41606, value : 32'h8034050}, //phyinit_io_write: 0x41605, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41607, value : 32'h0}, //phyinit_io_write: 0x41606, 0x8034050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41608, value : 32'h0}, //phyinit_io_write: 0x41607, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41609, value : 32'h4f000000}, //phyinit_io_write: 0x41608, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4160a, value : 32'h0}, //phyinit_io_write: 0x41609, 0x4f000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4160b, value : 32'h8000000}, //phyinit_io_write: 0x4160a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4160c, value : 32'h407c}, //phyinit_io_write: 0x4160b, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4160d, value : 32'h4000000}, //phyinit_io_write: 0x4160c, 0x407c
                          '{ step_type : REG_WRITE, reg_addr : 32'h4160e, value : 32'h0}, //phyinit_io_write: 0x4160d, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4160f, value : 32'h0}, //phyinit_io_write: 0x4160e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41610, value : 32'h0}, //phyinit_io_write: 0x4160f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41611, value : 32'h1f000000}, //phyinit_io_write: 0x41610, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41612, value : 32'h0}, //phyinit_io_write: 0x41611, 0x1f000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41613, value : 32'h0}, //phyinit_io_write: 0x41612, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41614, value : 32'h0}, //phyinit_io_write: 0x41613, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41615, value : 32'h4000001}, //phyinit_io_write: 0x41614, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41616, value : 32'h0}, //phyinit_io_write: 0x41615, 0x4000001
                          '{ step_type : REG_WRITE, reg_addr : 32'h41617, value : 32'h0}, //phyinit_io_write: 0x41616, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41618, value : 32'h0}, //phyinit_io_write: 0x41617, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41619, value : 32'h4000000}, //phyinit_io_write: 0x41618, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4161a, value : 32'h0}, //phyinit_io_write: 0x41619, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4161b, value : 32'h0}, //phyinit_io_write: 0x4161a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4161c, value : 32'h0}, //phyinit_io_write: 0x4161b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4161d, value : 32'h1b000000}, //phyinit_io_write: 0x4161c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4161e, value : 32'h0}, //phyinit_io_write: 0x4161d, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4161f, value : 32'h0}, //phyinit_io_write: 0x4161e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41620, value : 32'h0}, //phyinit_io_write: 0x4161f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41621, value : 32'h0}, //phyinit_io_write: 0x41620, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41622, value : 32'h0}, //phyinit_io_write: 0x41621, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41623, value : 32'h0}, //phyinit_io_write: 0x41622, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41624, value : 32'hd00802c}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 36
                          '{ step_type : REG_WRITE, reg_addr : 32'h41625, value : 32'h4100001}, //phyinit_io_write: 0x41624, 0xd00802c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41626, value : 32'h8008050}, //phyinit_io_write: 0x41625, 0x4100001
                          '{ step_type : REG_WRITE, reg_addr : 32'h41627, value : 32'h100000}, //phyinit_io_write: 0x41626, 0x8008050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41628, value : 32'h0}, //phyinit_io_write: 0x41627, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41629, value : 32'h4000000}, //phyinit_io_write: 0x41628, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4162a, value : 32'h8038050}, //phyinit_io_write: 0x41629, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4162b, value : 32'h100000}, //phyinit_io_write: 0x4162a, 0x8038050
                          '{ step_type : REG_WRITE, reg_addr : 32'h4162c, value : 32'h0}, //phyinit_io_write: 0x4162b, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4162d, value : 32'h4f000000}, //phyinit_io_write: 0x4162c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4162e, value : 32'h0}, //phyinit_io_write: 0x4162d, 0x4f000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4162f, value : 32'h8000000}, //phyinit_io_write: 0x4162e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41630, value : 32'h807c}, //phyinit_io_write: 0x4162f, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41631, value : 32'h4100000}, //phyinit_io_write: 0x41630, 0x807c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41632, value : 32'h0}, //phyinit_io_write: 0x41631, 0x4100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41633, value : 32'h0}, //phyinit_io_write: 0x41632, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41634, value : 32'h0}, //phyinit_io_write: 0x41633, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41635, value : 32'h1f000000}, //phyinit_io_write: 0x41634, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41636, value : 32'h0}, //phyinit_io_write: 0x41635, 0x1f000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41637, value : 32'h0}, //phyinit_io_write: 0x41636, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41638, value : 32'h0}, //phyinit_io_write: 0x41637, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41639, value : 32'h4000001}, //phyinit_io_write: 0x41638, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4163a, value : 32'h0}, //phyinit_io_write: 0x41639, 0x4000001
                          '{ step_type : REG_WRITE, reg_addr : 32'h4163b, value : 32'h0}, //phyinit_io_write: 0x4163a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4163c, value : 32'h0}, //phyinit_io_write: 0x4163b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4163d, value : 32'h4000000}, //phyinit_io_write: 0x4163c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4163e, value : 32'h0}, //phyinit_io_write: 0x4163d, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4163f, value : 32'h0}, //phyinit_io_write: 0x4163e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41640, value : 32'h0}, //phyinit_io_write: 0x4163f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41641, value : 32'h1b000000}, //phyinit_io_write: 0x41640, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41642, value : 32'h0}, //phyinit_io_write: 0x41641, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41643, value : 32'h0}, //phyinit_io_write: 0x41642, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41644, value : 32'h0}, //phyinit_io_write: 0x41643, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41645, value : 32'h0}, //phyinit_io_write: 0x41644, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41646, value : 32'h0}, //phyinit_io_write: 0x41645, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41647, value : 32'h0}, //phyinit_io_write: 0x41646, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41648, value : 32'hd00402c}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 72
                          '{ step_type : REG_WRITE, reg_addr : 32'h41649, value : 32'h1}, //phyinit_io_write: 0x41648, 0xd00402c
                          '{ step_type : REG_WRITE, reg_addr : 32'h4164a, value : 32'h8004050}, //phyinit_io_write: 0x41649, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4164b, value : 32'h0}, //phyinit_io_write: 0x4164a, 0x8004050
                          '{ step_type : REG_WRITE, reg_addr : 32'h4164c, value : 32'h0}, //phyinit_io_write: 0x4164b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4164d, value : 32'h0}, //phyinit_io_write: 0x4164c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4164e, value : 32'h8034050}, //phyinit_io_write: 0x4164d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4164f, value : 32'h0}, //phyinit_io_write: 0x4164e, 0x8034050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41650, value : 32'h0}, //phyinit_io_write: 0x4164f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41651, value : 32'h0}, //phyinit_io_write: 0x41650, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41652, value : 32'h8034050}, //phyinit_io_write: 0x41651, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41653, value : 32'h0}, //phyinit_io_write: 0x41652, 0x8034050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41654, value : 32'h0}, //phyinit_io_write: 0x41653, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41655, value : 32'h0}, //phyinit_io_write: 0x41654, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41656, value : 32'h8004050}, //phyinit_io_write: 0x41655, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41657, value : 32'h0}, //phyinit_io_write: 0x41656, 0x8004050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41658, value : 32'h0}, //phyinit_io_write: 0x41657, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41659, value : 32'h4b000000}, //phyinit_io_write: 0x41658, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4165a, value : 32'h0}, //phyinit_io_write: 0x41659, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4165b, value : 32'h8000000}, //phyinit_io_write: 0x4165a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4165c, value : 32'h407c}, //phyinit_io_write: 0x4165b, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4165d, value : 32'h0}, //phyinit_io_write: 0x4165c, 0x407c
                          '{ step_type : REG_WRITE, reg_addr : 32'h4165e, value : 32'h0}, //phyinit_io_write: 0x4165d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4165f, value : 32'h0}, //phyinit_io_write: 0x4165e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41660, value : 32'h0}, //phyinit_io_write: 0x4165f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41661, value : 32'h1b000000}, //phyinit_io_write: 0x41660, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41662, value : 32'h0}, //phyinit_io_write: 0x41661, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41663, value : 32'h0}, //phyinit_io_write: 0x41662, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41664, value : 32'h0}, //phyinit_io_write: 0x41663, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41665, value : 32'h1}, //phyinit_io_write: 0x41664, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41666, value : 32'h0}, //phyinit_io_write: 0x41665, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h41667, value : 32'h0}, //phyinit_io_write: 0x41666, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41668, value : 32'h0}, //phyinit_io_write: 0x41667, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41669, value : 32'h5b000000}, //phyinit_io_write: 0x41668, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4166a, value : 32'h0}, //phyinit_io_write: 0x41669, 0x5b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4166b, value : 32'h1c000000}, //phyinit_io_write: 0x4166a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4166c, value : 32'hd00802c}, //phyinit_io_write: 0x4166b, 0x1c000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4166d, value : 32'h100001}, //phyinit_io_write: 0x4166c, 0xd00802c
                          '{ step_type : REG_WRITE, reg_addr : 32'h4166e, value : 32'h8008050}, //phyinit_io_write: 0x4166d, 0x100001
                          '{ step_type : REG_WRITE, reg_addr : 32'h4166f, value : 32'h100000}, //phyinit_io_write: 0x4166e, 0x8008050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41670, value : 32'h0}, //phyinit_io_write: 0x4166f, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41671, value : 32'h0}, //phyinit_io_write: 0x41670, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41672, value : 32'h8038050}, //phyinit_io_write: 0x41671, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41673, value : 32'h100000}, //phyinit_io_write: 0x41672, 0x8038050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41674, value : 32'h0}, //phyinit_io_write: 0x41673, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41675, value : 32'h0}, //phyinit_io_write: 0x41674, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41676, value : 32'h8038050}, //phyinit_io_write: 0x41675, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41677, value : 32'h100000}, //phyinit_io_write: 0x41676, 0x8038050
                          '{ step_type : REG_WRITE, reg_addr : 32'h41678, value : 32'h0}, //phyinit_io_write: 0x41677, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41679, value : 32'h0}, //phyinit_io_write: 0x41678, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4167a, value : 32'h8008050}, //phyinit_io_write: 0x41679, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4167b, value : 32'h100000}, //phyinit_io_write: 0x4167a, 0x8008050
                          '{ step_type : REG_WRITE, reg_addr : 32'h4167c, value : 32'h0}, //phyinit_io_write: 0x4167b, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4167d, value : 32'h4b000000}, //phyinit_io_write: 0x4167c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4167e, value : 32'h0}, //phyinit_io_write: 0x4167d, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4167f, value : 32'h8000000}, //phyinit_io_write: 0x4167e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41680, value : 32'h807c}, //phyinit_io_write: 0x4167f, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41681, value : 32'h100000}, //phyinit_io_write: 0x41680, 0x807c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41682, value : 32'h0}, //phyinit_io_write: 0x41681, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41683, value : 32'h0}, //phyinit_io_write: 0x41682, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41684, value : 32'h0}, //phyinit_io_write: 0x41683, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41685, value : 32'h1b000000}, //phyinit_io_write: 0x41684, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41686, value : 32'h0}, //phyinit_io_write: 0x41685, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41687, value : 32'h0}, //phyinit_io_write: 0x41686, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41688, value : 32'h0}, //phyinit_io_write: 0x41687, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41689, value : 32'h1}, //phyinit_io_write: 0x41688, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4168a, value : 32'h0}, //phyinit_io_write: 0x41689, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4168b, value : 32'h0}, //phyinit_io_write: 0x4168a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4168c, value : 32'h0}, //phyinit_io_write: 0x4168b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4168d, value : 32'h2b000000}, //phyinit_io_write: 0x4168c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4168e, value : 32'h0}, //phyinit_io_write: 0x4168d, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4168f, value : 32'h28000000}, //phyinit_io_write: 0x4168e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41690, value : 32'hd00402c}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 68
                          '{ step_type : REG_WRITE, reg_addr : 32'h41691, value : 32'h1}, //phyinit_io_write: 0x41690, 0xd00402c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41692, value : 32'h8035198}, //phyinit_io_write: 0x41691, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h41693, value : 32'h0}, //phyinit_io_write: 0x41692, 0x8035198
                          '{ step_type : REG_WRITE, reg_addr : 32'h41694, value : 32'h0}, //phyinit_io_write: 0x41693, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41695, value : 32'h0}, //phyinit_io_write: 0x41694, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41696, value : 32'h0}, //phyinit_io_write: 0x41695, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41697, value : 32'h0}, //phyinit_io_write: 0x41696, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41698, value : 32'h0}, //phyinit_io_write: 0x41697, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41699, value : 32'h0}, //phyinit_io_write: 0x41698, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4169a, value : 32'h8035218}, //phyinit_io_write: 0x41699, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4169b, value : 32'h0}, //phyinit_io_write: 0x4169a, 0x8035218
                          '{ step_type : REG_WRITE, reg_addr : 32'h4169c, value : 32'h0}, //phyinit_io_write: 0x4169b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4169d, value : 32'h4b000000}, //phyinit_io_write: 0x4169c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4169e, value : 32'h0}, //phyinit_io_write: 0x4169d, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4169f, value : 32'h8000000}, //phyinit_io_write: 0x4169e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a0, value : 32'h407c}, //phyinit_io_write: 0x4169f, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a1, value : 32'h0}, //phyinit_io_write: 0x416a0, 0x407c
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a2, value : 32'h0}, //phyinit_io_write: 0x416a1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a3, value : 32'h0}, //phyinit_io_write: 0x416a2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a4, value : 32'h0}, //phyinit_io_write: 0x416a3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a5, value : 32'h1b000000}, //phyinit_io_write: 0x416a4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a6, value : 32'h0}, //phyinit_io_write: 0x416a5, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a7, value : 32'h0}, //phyinit_io_write: 0x416a6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a8, value : 32'h0}, //phyinit_io_write: 0x416a7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416a9, value : 32'h1}, //phyinit_io_write: 0x416a8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416aa, value : 32'h0}, //phyinit_io_write: 0x416a9, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h416ab, value : 32'h0}, //phyinit_io_write: 0x416aa, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416ac, value : 32'h0}, //phyinit_io_write: 0x416ab, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416ad, value : 32'h0}, //phyinit_io_write: 0x416ac, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416ae, value : 32'h0}, //phyinit_io_write: 0x416ad, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416af, value : 32'h0}, //phyinit_io_write: 0x416ae, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b0, value : 32'hd00802c}, //phyinit_io_write: 0x416af, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b1, value : 32'h100001}, //phyinit_io_write: 0x416b0, 0xd00802c
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b2, value : 32'h8039198}, //phyinit_io_write: 0x416b1, 0x100001
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b3, value : 32'h100000}, //phyinit_io_write: 0x416b2, 0x8039198
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b4, value : 32'h0}, //phyinit_io_write: 0x416b3, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b5, value : 32'h0}, //phyinit_io_write: 0x416b4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b6, value : 32'h0}, //phyinit_io_write: 0x416b5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b7, value : 32'h0}, //phyinit_io_write: 0x416b6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b8, value : 32'h0}, //phyinit_io_write: 0x416b7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416b9, value : 32'h0}, //phyinit_io_write: 0x416b8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416ba, value : 32'h8039218}, //phyinit_io_write: 0x416b9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416bb, value : 32'h100000}, //phyinit_io_write: 0x416ba, 0x8039218
                          '{ step_type : REG_WRITE, reg_addr : 32'h416bc, value : 32'h0}, //phyinit_io_write: 0x416bb, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416bd, value : 32'h4b000000}, //phyinit_io_write: 0x416bc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416be, value : 32'h0}, //phyinit_io_write: 0x416bd, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416bf, value : 32'h8000000}, //phyinit_io_write: 0x416be, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c0, value : 32'h807c}, //phyinit_io_write: 0x416bf, 0x8000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c1, value : 32'h100000}, //phyinit_io_write: 0x416c0, 0x807c
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c2, value : 32'h0}, //phyinit_io_write: 0x416c1, 0x100000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c3, value : 32'h0}, //phyinit_io_write: 0x416c2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c4, value : 32'h0}, //phyinit_io_write: 0x416c3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c5, value : 32'h1b000000}, //phyinit_io_write: 0x416c4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c6, value : 32'h0}, //phyinit_io_write: 0x416c5, 0x1b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c7, value : 32'h0}, //phyinit_io_write: 0x416c6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c8, value : 32'h0}, //phyinit_io_write: 0x416c7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416c9, value : 32'h1}, //phyinit_io_write: 0x416c8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416ca, value : 32'h0}, //phyinit_io_write: 0x416c9, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h416cb, value : 32'h0}, //phyinit_io_write: 0x416ca, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416cc, value : 32'h0}, //phyinit_io_write: 0x416cb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416cd, value : 32'h6b000000}, //phyinit_io_write: 0x416cc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416ce, value : 32'h0}, //phyinit_io_write: 0x416cd, 0x6b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h416cf, value : 32'h0}, //phyinit_io_write: 0x416ce, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416d0, value : 32'h0}, //phyinit_io_write: 0x416cf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416d1, value : 32'h0}, //phyinit_io_write: 0x416d0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416d2, value : 32'h0}, //phyinit_io_write: 0x416d1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416d3, value : 32'h0}, //phyinit_io_write: 0x416d2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416d4, value : 32'h0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h416d5, value : 32'h0}, //phyinit_io_write: 0x416d4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416d6, value : 32'h0}, //phyinit_io_write: 0x416d5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h416d7, value : 32'h0}, //phyinit_io_write: 0x416d6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44000, value : 32'h3f7ab480}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44001, value : 32'h16420}, //phyinit_io_write: 0x44000, 0x3f7ab480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44002, value : 32'h400}, //phyinit_io_write: 0x44001, 0x16420
                          '{ step_type : REG_WRITE, reg_addr : 32'h44003, value : 32'h0}, //phyinit_io_write: 0x44002, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44004, value : 32'h80000480}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 12
                          '{ step_type : REG_WRITE, reg_addr : 32'h44005, value : 32'hfc0}, //phyinit_io_write: 0x44004, 0x80000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44006, value : 32'h4000c00}, //phyinit_io_write: 0x44005, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44007, value : 32'h0}, //phyinit_io_write: 0x44006, 0x4000c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h44008, value : 32'h84000480}, //phyinit_io_write: 0x44007, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44009, value : 32'hc00}, //phyinit_io_write: 0x44008, 0x84000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4400a, value : 32'h4000800}, //phyinit_io_write: 0x44009, 0xc00
                          '{ step_type : REG_WRITE, reg_addr : 32'h4400b, value : 32'h0}, //phyinit_io_write: 0x4400a, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4400c, value : 32'h84000080}, //phyinit_io_write: 0x4400b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4400d, value : 32'hc00}, //phyinit_io_write: 0x4400c, 0x84000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4400e, value : 32'h1e0}, //phyinit_io_write: 0x4400d, 0xc00
                          '{ step_type : REG_WRITE, reg_addr : 32'h4400f, value : 32'h0}, //phyinit_io_write: 0x4400e, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44010, value : 32'h80068200}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44011, value : 32'h400f}, //phyinit_io_write: 0x44010, 0x80068200
                          '{ step_type : REG_WRITE, reg_addr : 32'h44012, value : 32'h8940}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 50
                          '{ step_type : REG_WRITE, reg_addr : 32'h44013, value : 32'h0}, //phyinit_io_write: 0x44012, 0x8940
                          '{ step_type : REG_WRITE, reg_addr : 32'h44014, value : 32'ha0000480}, //phyinit_io_write: 0x44013, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44015, value : 32'h2420}, //phyinit_io_write: 0x44014, 0xa0000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44016, value : 32'h4000400}, //phyinit_io_write: 0x44015, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h44017, value : 32'h0}, //phyinit_io_write: 0x44016, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44018, value : 32'h9c001ca0}, //phyinit_io_write: 0x44017, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44019, value : 32'h1c04}, //phyinit_io_write: 0x44018, 0x9c001ca0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4401a, value : 32'ha8000880}, //phyinit_io_write: 0x44019, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4401b, value : 32'h1c06}, //phyinit_io_write: 0x4401a, 0xa8000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4401c, value : 32'h80010080}, //phyinit_io_write: 0x4401b, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h4401d, value : 32'h1c04}, //phyinit_io_write: 0x4401c, 0x80010080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4401e, value : 32'h4000400}, //phyinit_io_write: 0x4401d, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4401f, value : 32'h0}, //phyinit_io_write: 0x4401e, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44020, value : 32'h80010480}, //phyinit_io_write: 0x4401f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44021, value : 32'h1c04}, //phyinit_io_write: 0x44020, 0x80010480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44022, value : 32'h4000800}, //phyinit_io_write: 0x44021, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44023, value : 32'h0}, //phyinit_io_write: 0x44022, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44024, value : 32'h40}, //phyinit_io_write: 0x44023, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44025, value : 32'h6000}, //phyinit_io_write: 0x44024, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h44026, value : 32'ha0000080}, //phyinit_io_write: 0x44025, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44027, value : 32'h2420}, //phyinit_io_write: 0x44026, 0xa0000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44028, value : 32'h1020}, //phyinit_io_write: 0x44027, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h44029, value : 32'h0}, //phyinit_io_write: 0x44028, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h4402a, value : 32'h1020}, //phyinit_io_write: 0x44029, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4402b, value : 32'h0}, //phyinit_io_write: 0x4402a, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h4402c, value : 32'h3020}, //phyinit_io_write: 0x4402b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4402d, value : 32'h0}, //phyinit_io_write: 0x4402c, 0x3020
                          '{ step_type : REG_WRITE, reg_addr : 32'h4402e, value : 32'h80000080}, //phyinit_io_write: 0x4402d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4402f, value : 32'h1c04}, //phyinit_io_write: 0x4402e, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44030, value : 32'ha8000880}, //phyinit_io_write: 0x4402f, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44031, value : 32'h1c06}, //phyinit_io_write: 0x44030, 0xa8000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44032, value : 32'h80010880}, //phyinit_io_write: 0x44031, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h44033, value : 32'h1c04}, //phyinit_io_write: 0x44032, 0x80010880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44034, value : 32'h4000400}, //phyinit_io_write: 0x44033, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44035, value : 32'h0}, //phyinit_io_write: 0x44034, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44036, value : 32'h80010c80}, //phyinit_io_write: 0x44035, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44037, value : 32'h1c04}, //phyinit_io_write: 0x44036, 0x80010c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44038, value : 32'h4000800}, //phyinit_io_write: 0x44037, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44039, value : 32'h0}, //phyinit_io_write: 0x44038, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4403a, value : 32'h1020}, //phyinit_io_write: 0x44039, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4403b, value : 32'h0}, //phyinit_io_write: 0x4403a, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h4403c, value : 32'h2c20}, //phyinit_io_write: 0x4403b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4403d, value : 32'h0}, //phyinit_io_write: 0x4403c, 0x2c20
                          '{ step_type : REG_WRITE, reg_addr : 32'h4403e, value : 32'h2c20}, //phyinit_io_write: 0x4403d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4403f, value : 32'h0}, //phyinit_io_write: 0x4403e, 0x2c20
                          '{ step_type : REG_WRITE, reg_addr : 32'h44040, value : 32'h2c20}, //phyinit_io_write: 0x4403f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44041, value : 32'h0}, //phyinit_io_write: 0x44040, 0x2c20
                          '{ step_type : REG_WRITE, reg_addr : 32'h44042, value : 32'h80000080}, //phyinit_io_write: 0x44041, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44043, value : 32'h1c04}, //phyinit_io_write: 0x44042, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44044, value : 32'h1e0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44045, value : 32'h0}, //phyinit_io_write: 0x44044, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44046, value : 32'ha8000480}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 6
                          '{ step_type : REG_WRITE, reg_addr : 32'h44047, value : 32'h1c04}, //phyinit_io_write: 0x44046, 0xa8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44048, value : 32'h4000400}, //phyinit_io_write: 0x44047, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44049, value : 32'h0}, //phyinit_io_write: 0x44048, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4404a, value : 32'h40004200}, //phyinit_io_write: 0x44049, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4404b, value : 32'h4000}, //phyinit_io_write: 0x4404a, 0x40004200
                          '{ step_type : REG_WRITE, reg_addr : 32'h4404c, value : 32'h10d40}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4404d, value : 32'h0}, //phyinit_io_write: 0x4404c, 0x10d40
                          '{ step_type : REG_WRITE, reg_addr : 32'h4404e, value : 32'hc80038a0}, //phyinit_io_write: 0x4404d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4404f, value : 32'h1c01}, //phyinit_io_write: 0x4404e, 0xc80038a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44050, value : 32'hcc003ca0}, //phyinit_io_write: 0x4404f, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44051, value : 32'h1c01}, //phyinit_io_write: 0x44050, 0xcc003ca0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44052, value : 32'ha40000a0}, //phyinit_io_write: 0x44051, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44053, value : 32'h1c06}, //phyinit_io_write: 0x44052, 0xa40000a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44054, value : 32'ha8001c80}, //phyinit_io_write: 0x44053, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h44055, value : 32'h1c06}, //phyinit_io_write: 0x44054, 0xa8001c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44056, value : 32'h80051080}, //phyinit_io_write: 0x44055, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h44057, value : 32'h1c04}, //phyinit_io_write: 0x44056, 0x80051080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44058, value : 32'h4000400}, //phyinit_io_write: 0x44057, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44059, value : 32'h0}, //phyinit_io_write: 0x44058, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4405a, value : 32'h80051480}, //phyinit_io_write: 0x44059, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4405b, value : 32'h1c04}, //phyinit_io_write: 0x4405a, 0x80051480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4405c, value : 32'h4000800}, //phyinit_io_write: 0x4405b, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4405d, value : 32'h0}, //phyinit_io_write: 0x4405c, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4405e, value : 32'h840}, //phyinit_io_write: 0x4405d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4405f, value : 32'h6000}, //phyinit_io_write: 0x4405e, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h44060, value : 32'h80000080}, //phyinit_io_write: 0x4405f, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44061, value : 32'h1c04}, //phyinit_io_write: 0x44060, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44062, value : 32'hcc000080}, //phyinit_io_write: 0x44061, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44063, value : 32'h1c01}, //phyinit_io_write: 0x44062, 0xcc000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44064, value : 32'ha8001c80}, //phyinit_io_write: 0x44063, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44065, value : 32'h1c06}, //phyinit_io_write: 0x44064, 0xa8001c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44066, value : 32'h80051880}, //phyinit_io_write: 0x44065, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h44067, value : 32'h1c04}, //phyinit_io_write: 0x44066, 0x80051880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44068, value : 32'h4000400}, //phyinit_io_write: 0x44067, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44069, value : 32'h0}, //phyinit_io_write: 0x44068, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4406a, value : 32'h80051c80}, //phyinit_io_write: 0x44069, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4406b, value : 32'h1c04}, //phyinit_io_write: 0x4406a, 0x80051c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h4406c, value : 32'h4000800}, //phyinit_io_write: 0x4406b, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4406d, value : 32'h0}, //phyinit_io_write: 0x4406c, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4406e, value : 32'h840}, //phyinit_io_write: 0x4406d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4406f, value : 32'h6000}, //phyinit_io_write: 0x4406e, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h44070, value : 32'h80000080}, //phyinit_io_write: 0x4406f, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44071, value : 32'h1c04}, //phyinit_io_write: 0x44070, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44072, value : 32'hc8000080}, //phyinit_io_write: 0x44071, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44073, value : 32'h1c01}, //phyinit_io_write: 0x44072, 0xc8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44074, value : 32'hcc003ca0}, //phyinit_io_write: 0x44073, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44075, value : 32'h1c01}, //phyinit_io_write: 0x44074, 0xcc003ca0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44076, value : 32'ha8001c80}, //phyinit_io_write: 0x44075, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44077, value : 32'h1c06}, //phyinit_io_write: 0x44076, 0xa8001c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44078, value : 32'h80052080}, //phyinit_io_write: 0x44077, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h44079, value : 32'h1c04}, //phyinit_io_write: 0x44078, 0x80052080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4407a, value : 32'h4000400}, //phyinit_io_write: 0x44079, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4407b, value : 32'h0}, //phyinit_io_write: 0x4407a, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4407c, value : 32'h80052480}, //phyinit_io_write: 0x4407b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4407d, value : 32'h1c04}, //phyinit_io_write: 0x4407c, 0x80052480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4407e, value : 32'h4000800}, //phyinit_io_write: 0x4407d, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4407f, value : 32'h0}, //phyinit_io_write: 0x4407e, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44080, value : 32'h840}, //phyinit_io_write: 0x4407f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44081, value : 32'h6000}, //phyinit_io_write: 0x44080, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h44082, value : 32'h80000080}, //phyinit_io_write: 0x44081, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44083, value : 32'h1c04}, //phyinit_io_write: 0x44082, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44084, value : 32'hc80038a0}, //phyinit_io_write: 0x44083, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44085, value : 32'h1c01}, //phyinit_io_write: 0x44084, 0xc80038a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44086, value : 32'h54000091}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h44087, value : 32'h18fc0}, //phyinit_io_write: 0x44086, 0x54000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h44088, value : 32'h54000091}, //phyinit_io_write: 0x44087, 0x18fc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44089, value : 32'h14fc0}, //phyinit_io_write: 0x44088, 0x54000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h4408a, value : 32'hf0000091}, //phyinit_io_write: 0x44089, 0x14fc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4408b, value : 32'h187c1}, //phyinit_io_write: 0x4408a, 0xf0000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h4408c, value : 32'hf0000091}, //phyinit_io_write: 0x4408b, 0x187c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4408d, value : 32'h147c1}, //phyinit_io_write: 0x4408c, 0xf0000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h4408e, value : 32'h8000611}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4408f, value : 32'h1800}, //phyinit_io_write: 0x4408e, 0x8000611
                          '{ step_type : REG_WRITE, reg_addr : 32'h44090, value : 32'h13971}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h44091, value : 32'h0}, //phyinit_io_write: 0x44090, 0x13971
                          '{ step_type : REG_WRITE, reg_addr : 32'h44092, value : 32'h4000911}, //phyinit_io_write: 0x44091, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44093, value : 32'h1a420}, //phyinit_io_write: 0x44092, 0x4000911
                          '{ step_type : REG_WRITE, reg_addr : 32'h44094, value : 32'h4001000}, //phyinit_io_write: 0x44093, 0x1a420
                          '{ step_type : REG_WRITE, reg_addr : 32'h44095, value : 32'h0}, //phyinit_io_write: 0x44094, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44096, value : 32'ha11}, //phyinit_io_write: 0x44095, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44097, value : 32'h1800}, //phyinit_io_write: 0x44096, 0xa11
                          '{ step_type : REG_WRITE, reg_addr : 32'h44098, value : 32'h17151}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44099, value : 32'h0}, //phyinit_io_write: 0x44098, 0x17151
                          '{ step_type : REG_WRITE, reg_addr : 32'h4409a, value : 32'h14171}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4409b, value : 32'h0}, //phyinit_io_write: 0x4409a, 0x14171
                          '{ step_type : REG_WRITE, reg_addr : 32'h4409c, value : 32'h611}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4409d, value : 32'h1800}, //phyinit_io_write: 0x4409c, 0x611
                          '{ step_type : REG_WRITE, reg_addr : 32'h4409e, value : 32'h17171}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4409f, value : 32'h0}, //phyinit_io_write: 0x4409e, 0x17171
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a0, value : 32'h24000491}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a1, value : 32'h1e420}, //phyinit_io_write: 0x440a0, 0x24000491
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a2, value : 32'h21d1}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 22
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a3, value : 32'h0}, //phyinit_io_write: 0x440a2, 0x21d1
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a4, value : 32'h1031}, //phyinit_io_write: 0x440a3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a5, value : 32'h0}, //phyinit_io_write: 0x440a4, 0x1031
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a6, value : 32'h1031}, //phyinit_io_write: 0x440a5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a7, value : 32'h0}, //phyinit_io_write: 0x440a6, 0x1031
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a8, value : 32'h2c31}, //phyinit_io_write: 0x440a7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440a9, value : 32'h0}, //phyinit_io_write: 0x440a8, 0x2c31
                          '{ step_type : REG_WRITE, reg_addr : 32'h440aa, value : 32'ha8000091}, //phyinit_io_write: 0x440a9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ab, value : 32'h1c06}, //phyinit_io_write: 0x440aa, 0xa8000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ac, value : 32'h80016891}, //phyinit_io_write: 0x440ab, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ad, value : 32'h1c04}, //phyinit_io_write: 0x440ac, 0x80016891
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ae, value : 32'h4000400}, //phyinit_io_write: 0x440ad, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h440af, value : 32'h0}, //phyinit_io_write: 0x440ae, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b0, value : 32'h80016c91}, //phyinit_io_write: 0x440af, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b1, value : 32'h1c04}, //phyinit_io_write: 0x440b0, 0x80016c91
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b2, value : 32'h4000800}, //phyinit_io_write: 0x440b1, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b3, value : 32'h0}, //phyinit_io_write: 0x440b2, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b4, value : 32'h851}, //phyinit_io_write: 0x440b3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b5, value : 32'h6000}, //phyinit_io_write: 0x440b4, 0x851
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b6, value : 32'h80000091}, //phyinit_io_write: 0x440b5, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b7, value : 32'h1c04}, //phyinit_io_write: 0x440b6, 0x80000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b8, value : 32'ha8000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h440b9, value : 32'h1c04}, //phyinit_io_write: 0x440b8, 0xa8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ba, value : 32'h4000800}, //phyinit_io_write: 0x440b9, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h440bb, value : 32'h0}, //phyinit_io_write: 0x440ba, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h440bc, value : 32'h1e0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h440bd, value : 32'h0}, //phyinit_io_write: 0x440bc, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440be, value : 32'ha8000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 10
                          '{ step_type : REG_WRITE, reg_addr : 32'h440bf, value : 32'h1c06}, //phyinit_io_write: 0x440be, 0xa8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c0, value : 32'h80012880}, //phyinit_io_write: 0x440bf, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c1, value : 32'h1c04}, //phyinit_io_write: 0x440c0, 0x80012880
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c2, value : 32'h4000400}, //phyinit_io_write: 0x440c1, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c3, value : 32'h0}, //phyinit_io_write: 0x440c2, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c4, value : 32'h80012c80}, //phyinit_io_write: 0x440c3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c5, value : 32'h1c04}, //phyinit_io_write: 0x440c4, 0x80012c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c6, value : 32'h4000800}, //phyinit_io_write: 0x440c5, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c7, value : 32'h0}, //phyinit_io_write: 0x440c6, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c8, value : 32'h840}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 6
                          '{ step_type : REG_WRITE, reg_addr : 32'h440c9, value : 32'h6000}, //phyinit_io_write: 0x440c8, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ca, value : 32'h80000080}, //phyinit_io_write: 0x440c9, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h440cb, value : 32'h1c04}, //phyinit_io_write: 0x440ca, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h440cc, value : 32'h1e0}, //phyinit_io_write: 0x440cb, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h440cd, value : 32'h0}, //phyinit_io_write: 0x440cc, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ce, value : 32'h80200}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h440cf, value : 32'h400e}, //phyinit_io_write: 0x440ce, 0x80200
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d0, value : 32'h1b140}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d1, value : 32'h0}, //phyinit_io_write: 0x440d0, 0x1b140
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d2, value : 32'h20200}, //phyinit_io_write: 0x440d1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d3, value : 32'h400e}, //phyinit_io_write: 0x440d2, 0x20200
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d4, value : 32'h1b140}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d5, value : 32'h0}, //phyinit_io_write: 0x440d4, 0x1b140
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d6, value : 32'h80068200}, //phyinit_io_write: 0x440d5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d7, value : 32'h400f}, //phyinit_io_write: 0x440d6, 0x80068200
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d8, value : 32'h30000cc0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h440d9, value : 32'h7c4}, //phyinit_io_write: 0x440d8, 0x30000cc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440da, value : 32'h1e0}, //phyinit_io_write: 0x440d9, 0x7c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h440db, value : 32'h0}, //phyinit_io_write: 0x440da, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440dc, value : 32'h100600}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 116
                          '{ step_type : REG_WRITE, reg_addr : 32'h440dd, value : 32'h10}, //phyinit_io_write: 0x440dc, 0x100600
                          '{ step_type : REG_WRITE, reg_addr : 32'h440de, value : 32'h2c0004c0}, //phyinit_io_write: 0x440dd, 0x10
                          '{ step_type : REG_WRITE, reg_addr : 32'h440df, value : 32'h3c0}, //phyinit_io_write: 0x440de, 0x2c0004c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e0, value : 32'h8c0028a0}, //phyinit_io_write: 0x440df, 0x3c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e1, value : 32'h17bc1}, //phyinit_io_write: 0x440e0, 0x8c0028a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e2, value : 32'ha0000480}, //phyinit_io_write: 0x440e1, 0x17bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e3, value : 32'h2420}, //phyinit_io_write: 0x440e2, 0xa0000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e4, value : 32'h4000400}, //phyinit_io_write: 0x440e3, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e5, value : 32'h0}, //phyinit_io_write: 0x440e4, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e6, value : 32'h8c0014a0}, //phyinit_io_write: 0x440e5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e7, value : 32'h143c1}, //phyinit_io_write: 0x440e6, 0x8c0014a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e8, value : 32'ha0000080}, //phyinit_io_write: 0x440e7, 0x143c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h440e9, value : 32'h2420}, //phyinit_io_write: 0x440e8, 0xa0000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ea, value : 32'h78000480}, //phyinit_io_write: 0x440e9, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h440eb, value : 32'h3d8}, //phyinit_io_write: 0x440ea, 0x78000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ec, value : 32'h7c000480}, //phyinit_io_write: 0x440eb, 0x3d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ed, value : 32'h7f8}, //phyinit_io_write: 0x440ec, 0x7c000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ee, value : 32'h8000080}, //phyinit_io_write: 0x440ed, 0x7f8
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ef, value : 32'hfe0}, //phyinit_io_write: 0x440ee, 0x8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f0, value : 32'h8000080}, //phyinit_io_write: 0x440ef, 0xfe0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f1, value : 32'h7e0}, //phyinit_io_write: 0x440f0, 0x8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f2, value : 32'h80600}, //phyinit_io_write: 0x440f1, 0x7e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f3, value : 32'h8}, //phyinit_io_write: 0x440f2, 0x80600
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f4, value : 32'h4c0}, //phyinit_io_write: 0x440f3, 0x8
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f5, value : 32'h14fc4}, //phyinit_io_write: 0x440f4, 0x4c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f6, value : 32'h4c0}, //phyinit_io_write: 0x440f5, 0x14fc4
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f7, value : 32'h147c4}, //phyinit_io_write: 0x440f6, 0x4c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f8, value : 32'h2420}, //phyinit_io_write: 0x440f7, 0x147c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h440f9, value : 32'h0}, //phyinit_io_write: 0x440f8, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h440fa, value : 32'h8000480}, //phyinit_io_write: 0x440f9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440fb, value : 32'hfe0}, //phyinit_io_write: 0x440fa, 0x8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h440fc, value : 32'h8000480}, //phyinit_io_write: 0x440fb, 0xfe0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440fd, value : 32'h7e0}, //phyinit_io_write: 0x440fc, 0x8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h440fe, value : 32'h80}, //phyinit_io_write: 0x440fd, 0x7e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h440ff, value : 32'h14fc4}, //phyinit_io_write: 0x440fe, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44100, value : 32'h80}, //phyinit_io_write: 0x440ff, 0x14fc4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44101, value : 32'h147c4}, //phyinit_io_write: 0x44100, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44102, value : 32'h78000080}, //phyinit_io_write: 0x44101, 0x147c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44103, value : 32'h3d8}, //phyinit_io_write: 0x44102, 0x78000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44104, value : 32'h7c000080}, //phyinit_io_write: 0x44103, 0x3d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h44105, value : 32'h7f8}, //phyinit_io_write: 0x44104, 0x7c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44106, value : 32'h8c002ca0}, //phyinit_io_write: 0x44105, 0x7f8
                          '{ step_type : REG_WRITE, reg_addr : 32'h44107, value : 32'h17bc1}, //phyinit_io_write: 0x44106, 0x8c002ca0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44108, value : 32'ha0000480}, //phyinit_io_write: 0x44107, 0x17bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44109, value : 32'h2420}, //phyinit_io_write: 0x44108, 0xa0000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4410a, value : 32'h4000400}, //phyinit_io_write: 0x44109, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h4410b, value : 32'h0}, //phyinit_io_write: 0x4410a, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4410c, value : 32'h8c0018a0}, //phyinit_io_write: 0x4410b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4410d, value : 32'h143c1}, //phyinit_io_write: 0x4410c, 0x8c0018a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4410e, value : 32'ha0000080}, //phyinit_io_write: 0x4410d, 0x143c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4410f, value : 32'h2420}, //phyinit_io_write: 0x4410e, 0xa0000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44110, value : 32'h2c000080}, //phyinit_io_write: 0x4410f, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h44111, value : 32'h0}, //phyinit_io_write: 0x44110, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44112, value : 32'h2c000080}, //phyinit_io_write: 0x44111, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44113, value : 32'h40}, //phyinit_io_write: 0x44112, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44114, value : 32'h2c000080}, //phyinit_io_write: 0x44113, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h44115, value : 32'h80}, //phyinit_io_write: 0x44114, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44116, value : 32'h2c000080}, //phyinit_io_write: 0x44115, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44117, value : 32'hc0}, //phyinit_io_write: 0x44116, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44118, value : 32'h2c000080}, //phyinit_io_write: 0x44117, 0xc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44119, value : 32'h100}, //phyinit_io_write: 0x44118, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4411a, value : 32'h2c000080}, //phyinit_io_write: 0x44119, 0x100
                          '{ step_type : REG_WRITE, reg_addr : 32'h4411b, value : 32'h140}, //phyinit_io_write: 0x4411a, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4411c, value : 32'h200600}, //phyinit_io_write: 0x4411b, 0x140
                          '{ step_type : REG_WRITE, reg_addr : 32'h4411d, value : 32'h20}, //phyinit_io_write: 0x4411c, 0x200600
                          '{ step_type : REG_WRITE, reg_addr : 32'h4411e, value : 32'h2c0000c0}, //phyinit_io_write: 0x4411d, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h4411f, value : 32'h1c0}, //phyinit_io_write: 0x4411e, 0x2c0000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44120, value : 32'h2c0000c0}, //phyinit_io_write: 0x4411f, 0x1c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44121, value : 32'h200}, //phyinit_io_write: 0x44120, 0x2c0000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44122, value : 32'h2c0000c0}, //phyinit_io_write: 0x44121, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h44123, value : 32'h240}, //phyinit_io_write: 0x44122, 0x2c0000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44124, value : 32'h2c0000c0}, //phyinit_io_write: 0x44123, 0x240
                          '{ step_type : REG_WRITE, reg_addr : 32'h44125, value : 32'h280}, //phyinit_io_write: 0x44124, 0x2c0000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44126, value : 32'h2c0000c0}, //phyinit_io_write: 0x44125, 0x280
                          '{ step_type : REG_WRITE, reg_addr : 32'h44127, value : 32'h2c0}, //phyinit_io_write: 0x44126, 0x2c0000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44128, value : 32'h2c0000c0}, //phyinit_io_write: 0x44127, 0x2c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44129, value : 32'h300}, //phyinit_io_write: 0x44128, 0x2c0000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4412a, value : 32'hc4000880}, //phyinit_io_write: 0x44129, 0x300
                          '{ step_type : REG_WRITE, reg_addr : 32'h4412b, value : 32'h7c0}, //phyinit_io_write: 0x4412a, 0xc4000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4412c, value : 32'h4000400}, //phyinit_io_write: 0x4412b, 0x7c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4412d, value : 32'h0}, //phyinit_io_write: 0x4412c, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4412e, value : 32'hc000480}, //phyinit_io_write: 0x4412d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4412f, value : 32'hfc4}, //phyinit_io_write: 0x4412e, 0xc000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44130, value : 32'h4002000}, //phyinit_io_write: 0x4412f, 0xfc4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44131, value : 32'h0}, //phyinit_io_write: 0x44130, 0x4002000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44132, value : 32'hc000480}, //phyinit_io_write: 0x44131, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44133, value : 32'h7c4}, //phyinit_io_write: 0x44132, 0xc000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44134, value : 32'h4002000}, //phyinit_io_write: 0x44133, 0x7c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44135, value : 32'h0}, //phyinit_io_write: 0x44134, 0x4002000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44136, value : 32'hc000080}, //phyinit_io_write: 0x44135, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44137, value : 32'hfc4}, //phyinit_io_write: 0x44136, 0xc000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44138, value : 32'hc000080}, //phyinit_io_write: 0x44137, 0xfc4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44139, value : 32'h7c4}, //phyinit_io_write: 0x44138, 0xc000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4413a, value : 32'hc4000080}, //phyinit_io_write: 0x44139, 0x7c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4413b, value : 32'h7c0}, //phyinit_io_write: 0x4413a, 0xc4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4413c, value : 32'h4000400}, //phyinit_io_write: 0x4413b, 0x7c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4413d, value : 32'h0}, //phyinit_io_write: 0x4413c, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4413e, value : 32'he0000480}, //phyinit_io_write: 0x4413d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4413f, value : 32'h803}, //phyinit_io_write: 0x4413e, 0xe0000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44140, value : 32'h4002000}, //phyinit_io_write: 0x4413f, 0x803
                          '{ step_type : REG_WRITE, reg_addr : 32'h44141, value : 32'h0}, //phyinit_io_write: 0x44140, 0x4002000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44142, value : 32'h4000600}, //phyinit_io_write: 0x44141, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44143, value : 32'h400}, //phyinit_io_write: 0x44142, 0x4000600
                          '{ step_type : REG_WRITE, reg_addr : 32'h44144, value : 32'h265a58c0}, //phyinit_io_write: 0x44143, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44145, value : 32'h187c8}, //phyinit_io_write: 0x44144, 0x265a58c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44146, value : 32'h58000080}, //phyinit_io_write: 0x44145, 0x187c8
                          '{ step_type : REG_WRITE, reg_addr : 32'h44147, value : 32'h7c0}, //phyinit_io_write: 0x44146, 0x58000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44148, value : 32'h4000400}, //phyinit_io_write: 0x44147, 0x7c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44149, value : 32'h0}, //phyinit_io_write: 0x44148, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4414a, value : 32'he0000080}, //phyinit_io_write: 0x44149, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4414b, value : 32'h803}, //phyinit_io_write: 0x4414a, 0xe0000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4414c, value : 32'h4002000}, //phyinit_io_write: 0x4414b, 0x803
                          '{ step_type : REG_WRITE, reg_addr : 32'h4414d, value : 32'h0}, //phyinit_io_write: 0x4414c, 0x4002000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4414e, value : 32'h1e0}, //phyinit_io_write: 0x4414d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4414f, value : 32'h0}, //phyinit_io_write: 0x4414e, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44150, value : 32'h50000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 38
                          '{ step_type : REG_WRITE, reg_addr : 32'h44151, value : 32'h1c01}, //phyinit_io_write: 0x44150, 0x50000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44152, value : 32'h40000480}, //phyinit_io_write: 0x44151, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44153, value : 32'h2c0c}, //phyinit_io_write: 0x44152, 0x40000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44154, value : 32'hc4000080}, //phyinit_io_write: 0x44153, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h44155, value : 32'h7c0}, //phyinit_io_write: 0x44154, 0xc4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44156, value : 32'h2c000080}, //phyinit_io_write: 0x44155, 0x7c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44157, value : 32'h7c2}, //phyinit_io_write: 0x44156, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44158, value : 32'h8c200080}, //phyinit_io_write: 0x44157, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44159, value : 32'hfc2}, //phyinit_io_write: 0x44158, 0x8c200080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4415a, value : 32'h200600}, //phyinit_io_write: 0x44159, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4415b, value : 32'h20}, //phyinit_io_write: 0x4415a, 0x200600
                          '{ step_type : REG_WRITE, reg_addr : 32'h4415c, value : 32'h880c0080}, //phyinit_io_write: 0x4415b, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h4415d, value : 32'hc02}, //phyinit_io_write: 0x4415c, 0x880c0080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4415e, value : 32'h880c00c0}, //phyinit_io_write: 0x4415d, 0xc02
                          '{ step_type : REG_WRITE, reg_addr : 32'h4415f, value : 32'hc42}, //phyinit_io_write: 0x4415e, 0x880c00c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44160, value : 32'h247ffc80}, //phyinit_io_write: 0x4415f, 0xc42
                          '{ step_type : REG_WRITE, reg_addr : 32'h44161, value : 32'h7c2}, //phyinit_io_write: 0x44160, 0x247ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44162, value : 32'h281ffc80}, //phyinit_io_write: 0x44161, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44163, value : 32'h7c2}, //phyinit_io_write: 0x44162, 0x281ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44164, value : 32'h4000400}, //phyinit_io_write: 0x44163, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44165, value : 32'h0}, //phyinit_io_write: 0x44164, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44166, value : 32'h800c0080}, //phyinit_io_write: 0x44165, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44167, value : 32'hfc2}, //phyinit_io_write: 0x44166, 0x800c0080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44168, value : 32'h4000800}, //phyinit_io_write: 0x44167, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44169, value : 32'h0}, //phyinit_io_write: 0x44168, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4416a, value : 32'h98000480}, //phyinit_io_write: 0x44169, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4416b, value : 32'hfc2}, //phyinit_io_write: 0x4416a, 0x98000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4416c, value : 32'h28000480}, //phyinit_io_write: 0x4416b, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4416d, value : 32'hfc0}, //phyinit_io_write: 0x4416c, 0x28000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4416e, value : 32'h4001000}, //phyinit_io_write: 0x4416d, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4416f, value : 32'h0}, //phyinit_io_write: 0x4416e, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44170, value : 32'h80fffc80}, //phyinit_io_write: 0x4416f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44171, value : 32'hfc2}, //phyinit_io_write: 0x44170, 0x80fffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44172, value : 32'h30000080}, //phyinit_io_write: 0x44171, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44173, value : 32'h7c4}, //phyinit_io_write: 0x44172, 0x30000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44174, value : 32'h10600}, //phyinit_io_write: 0x44173, 0x7c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44175, value : 32'h1}, //phyinit_io_write: 0x44174, 0x10600
                          '{ step_type : REG_WRITE, reg_addr : 32'h44176, value : 32'h2f940}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44177, value : 32'h0}, //phyinit_io_write: 0x44176, 0x2f940
                          '{ step_type : REG_WRITE, reg_addr : 32'h44178, value : 32'h80068200}, //phyinit_io_write: 0x44177, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44179, value : 32'h400f}, //phyinit_io_write: 0x44178, 0x80068200
                          '{ step_type : REG_WRITE, reg_addr : 32'h4417a, value : 32'h2fd60}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4417b, value : 32'h0}, //phyinit_io_write: 0x4417a, 0x2fd60
                          '{ step_type : REG_WRITE, reg_addr : 32'h4417c, value : 32'h19dc0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4417d, value : 32'h0}, //phyinit_io_write: 0x4417c, 0x19dc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4417e, value : 32'he0000480}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 30
                          '{ step_type : REG_WRITE, reg_addr : 32'h4417f, value : 32'h803}, //phyinit_io_write: 0x4417e, 0xe0000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44180, value : 32'h4001c00}, //phyinit_io_write: 0x4417f, 0x803
                          '{ step_type : REG_WRITE, reg_addr : 32'h44181, value : 32'h0}, //phyinit_io_write: 0x44180, 0x4001c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h44182, value : 32'h28000080}, //phyinit_io_write: 0x44181, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44183, value : 32'hfc0}, //phyinit_io_write: 0x44182, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44184, value : 32'h88000480}, //phyinit_io_write: 0x44183, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44185, value : 32'h802}, //phyinit_io_write: 0x44184, 0x88000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44186, value : 32'h4000400}, //phyinit_io_write: 0x44185, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h44187, value : 32'h0}, //phyinit_io_write: 0x44186, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44188, value : 32'h5c000080}, //phyinit_io_write: 0x44187, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44189, value : 32'h7c2}, //phyinit_io_write: 0x44188, 0x5c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4418a, value : 32'h2000600}, //phyinit_io_write: 0x44189, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4418b, value : 32'h200}, //phyinit_io_write: 0x4418a, 0x2000600
                          '{ step_type : REG_WRITE, reg_addr : 32'h4418c, value : 32'h2c0010c0}, //phyinit_io_write: 0x4418b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h4418d, value : 32'h3bc1}, //phyinit_io_write: 0x4418c, 0x2c0010c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4418e, value : 32'h2c001880}, //phyinit_io_write: 0x4418d, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4418f, value : 32'h3bc1}, //phyinit_io_write: 0x4418e, 0x2c001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44190, value : 32'h18001880}, //phyinit_io_write: 0x4418f, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44191, value : 32'h3bc1}, //phyinit_io_write: 0x44190, 0x18001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44192, value : 32'h1c001880}, //phyinit_io_write: 0x44191, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44193, value : 32'h3bc1}, //phyinit_io_write: 0x44192, 0x1c001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44194, value : 32'h20001880}, //phyinit_io_write: 0x44193, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44195, value : 32'h3bc1}, //phyinit_io_write: 0x44194, 0x20001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44196, value : 32'h24001880}, //phyinit_io_write: 0x44195, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44197, value : 32'h3bc1}, //phyinit_io_write: 0x44196, 0x24001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44198, value : 32'h28001880}, //phyinit_io_write: 0x44197, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44199, value : 32'h3bc1}, //phyinit_io_write: 0x44198, 0x28001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4419a, value : 32'h20200}, //phyinit_io_write: 0x44199, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4419b, value : 32'h400e}, //phyinit_io_write: 0x4419a, 0x20200
                          '{ step_type : REG_WRITE, reg_addr : 32'h4419c, value : 32'h36940}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4419d, value : 32'h0}, //phyinit_io_write: 0x4419c, 0x36940
                          '{ step_type : REG_WRITE, reg_addr : 32'h4419e, value : 32'h40004600}, //phyinit_io_write: 0x4419d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4419f, value : 32'h0}, //phyinit_io_write: 0x4419e, 0x40004600
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a0, value : 32'h35540}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 10
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a1, value : 32'h0}, //phyinit_io_write: 0x441a0, 0x35540
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a2, value : 32'h4000900}, //phyinit_io_write: 0x441a1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a3, value : 32'h1a420}, //phyinit_io_write: 0x441a2, 0x4000900
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a4, value : 32'h4001000}, //phyinit_io_write: 0x441a3, 0x1a420
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a5, value : 32'h0}, //phyinit_io_write: 0x441a4, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a6, value : 32'h40004a00}, //phyinit_io_write: 0x441a5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a7, value : 32'h0}, //phyinit_io_write: 0x441a6, 0x40004a00
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a8, value : 32'hc0010e0}, //phyinit_io_write: 0x441a7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441a9, value : 32'h1800}, //phyinit_io_write: 0x441a8, 0xc0010e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441aa, value : 32'hc0000c0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 10
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ab, value : 32'h1800}, //phyinit_io_write: 0x441aa, 0xc0000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ac, value : 32'h4000480}, //phyinit_io_write: 0x441ab, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ad, value : 32'h1800}, //phyinit_io_write: 0x441ac, 0x4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ae, value : 32'h4000800}, //phyinit_io_write: 0x441ad, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441af, value : 32'h0}, //phyinit_io_write: 0x441ae, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b0, value : 32'h8000480}, //phyinit_io_write: 0x441af, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b1, value : 32'h1800}, //phyinit_io_write: 0x441b0, 0x8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b2, value : 32'h4000800}, //phyinit_io_write: 0x441b1, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b3, value : 32'h0}, //phyinit_io_write: 0x441b2, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b4, value : 32'h1e0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b5, value : 32'h0}, //phyinit_io_write: 0x441b4, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b6, value : 32'h9c000cb1}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b7, value : 32'h1c01}, //phyinit_io_write: 0x441b6, 0x9c000cb1
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b8, value : 32'h9c0010b1}, //phyinit_io_write: 0x441b7, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h441b9, value : 32'h1c03}, //phyinit_io_write: 0x441b8, 0x9c0010b1
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ba, value : 32'h24000091}, //phyinit_io_write: 0x441b9, 0x1c03
                          '{ step_type : REG_WRITE, reg_addr : 32'h441bb, value : 32'h1c01}, //phyinit_io_write: 0x441ba, 0x24000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h441bc, value : 32'h51}, //phyinit_io_write: 0x441bb, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h441bd, value : 32'h4000}, //phyinit_io_write: 0x441bc, 0x51
                          '{ step_type : REG_WRITE, reg_addr : 32'h441be, value : 32'h39131}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h441bf, value : 32'h0}, //phyinit_io_write: 0x441be, 0x39131
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c0, value : 32'h40001a01}, //phyinit_io_write: 0x441bf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c1, value : 32'h0}, //phyinit_io_write: 0x441c0, 0x40001a01
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c2, value : 32'h39161}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 6
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c3, value : 32'h0}, //phyinit_io_write: 0x441c2, 0x39161
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c4, value : 32'h24000081}, //phyinit_io_write: 0x441c3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c5, value : 32'h1c01}, //phyinit_io_write: 0x441c4, 0x24000081
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c6, value : 32'h41}, //phyinit_io_write: 0x441c5, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c7, value : 32'h4000}, //phyinit_io_write: 0x441c6, 0x41
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c8, value : 32'h1e0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h441c9, value : 32'h0}, //phyinit_io_write: 0x441c8, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ca, value : 32'h84000900}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h441cb, value : 32'h241c}, //phyinit_io_write: 0x441ca, 0x84000900
                          '{ step_type : REG_WRITE, reg_addr : 32'h441cc, value : 32'hc0014200}, //phyinit_io_write: 0x441cb, 0x241c
                          '{ step_type : REG_WRITE, reg_addr : 32'h441cd, value : 32'hc001}, //phyinit_io_write: 0x441cc, 0xc0014200
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ce, value : 32'h3a940}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 6
                          '{ step_type : REG_WRITE, reg_addr : 32'h441cf, value : 32'h0}, //phyinit_io_write: 0x441ce, 0x3a940
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d0, value : 32'h4001000}, //phyinit_io_write: 0x441cf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d1, value : 32'h0}, //phyinit_io_write: 0x441d0, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d2, value : 32'h2c0008a0}, //phyinit_io_write: 0x441d1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d3, value : 32'h802}, //phyinit_io_write: 0x441d2, 0x2c0008a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d4, value : 32'h1e0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d5, value : 32'h0}, //phyinit_io_write: 0x441d4, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d6, value : 32'h40000480}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 10
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d7, value : 32'h2c0c}, //phyinit_io_write: 0x441d6, 0x40000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d8, value : 32'h4000400}, //phyinit_io_write: 0x441d7, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h441d9, value : 32'h0}, //phyinit_io_write: 0x441d8, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h441da, value : 32'h4000080}, //phyinit_io_write: 0x441d9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441db, value : 32'h2c00}, //phyinit_io_write: 0x441da, 0x4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h441dc, value : 32'h4000400}, //phyinit_io_write: 0x441db, 0x2c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h441dd, value : 32'h0}, //phyinit_io_write: 0x441dc, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h441de, value : 32'h20200}, //phyinit_io_write: 0x441dd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441df, value : 32'h400e}, //phyinit_io_write: 0x441de, 0x20200
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e0, value : 32'h44140}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e1, value : 32'h0}, //phyinit_io_write: 0x441e0, 0x44140
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e2, value : 32'h40004600}, //phyinit_io_write: 0x441e1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e3, value : 32'h0}, //phyinit_io_write: 0x441e2, 0x40004600
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e4, value : 32'h40004c0}, //phyinit_io_write: 0x441e3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e5, value : 32'h1800}, //phyinit_io_write: 0x441e4, 0x40004c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e6, value : 32'h80004c0}, //phyinit_io_write: 0x441e5, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e7, value : 32'h1800}, //phyinit_io_write: 0x441e6, 0x80004c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e8, value : 32'h44140}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 22
                          '{ step_type : REG_WRITE, reg_addr : 32'h441e9, value : 32'h0}, //phyinit_io_write: 0x441e8, 0x44140
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ea, value : 32'h8000080}, //phyinit_io_write: 0x441e9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441eb, value : 32'h1800}, //phyinit_io_write: 0x441ea, 0x8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ec, value : 32'h4000400}, //phyinit_io_write: 0x441eb, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ed, value : 32'h0}, //phyinit_io_write: 0x441ec, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ee, value : 32'h4000080}, //phyinit_io_write: 0x441ed, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ef, value : 32'h1800}, //phyinit_io_write: 0x441ee, 0x4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f0, value : 32'h81}, //phyinit_io_write: 0x441ef, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f1, value : 32'h1800}, //phyinit_io_write: 0x441f0, 0x81
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f2, value : 32'h4000400}, //phyinit_io_write: 0x441f1, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f3, value : 32'h0}, //phyinit_io_write: 0x441f2, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f4, value : 32'h88000480}, //phyinit_io_write: 0x441f3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f5, value : 32'h802}, //phyinit_io_write: 0x441f4, 0x88000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f6, value : 32'h4000800}, //phyinit_io_write: 0x441f5, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f7, value : 32'h0}, //phyinit_io_write: 0x441f6, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f8, value : 32'hc000900}, //phyinit_io_write: 0x441f7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441f9, value : 32'h1800}, //phyinit_io_write: 0x441f8, 0xc000900
                          '{ step_type : REG_WRITE, reg_addr : 32'h441fa, value : 32'h4001000}, //phyinit_io_write: 0x441f9, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h441fb, value : 32'h0}, //phyinit_io_write: 0x441fa, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h441fc, value : 32'h10a00}, //phyinit_io_write: 0x441fb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h441fd, value : 32'h1}, //phyinit_io_write: 0x441fc, 0x10a00
                          '{ step_type : REG_WRITE, reg_addr : 32'h441fe, value : 32'h41d40}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 14
                          '{ step_type : REG_WRITE, reg_addr : 32'h441ff, value : 32'h0}, //phyinit_io_write: 0x441fe, 0x41d40
                          '{ step_type : REG_WRITE, reg_addr : 32'h44200, value : 32'hc000c80}, //phyinit_io_write: 0x441ff, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44201, value : 32'h1800}, //phyinit_io_write: 0x44200, 0xc000c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44202, value : 32'h20}, //phyinit_io_write: 0x44201, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44203, value : 32'h0}, //phyinit_io_write: 0x44202, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h44204, value : 32'h20}, //phyinit_io_write: 0x44203, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44205, value : 32'h0}, //phyinit_io_write: 0x44204, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h44206, value : 32'hc000880}, //phyinit_io_write: 0x44205, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44207, value : 32'h1800}, //phyinit_io_write: 0x44206, 0xc000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44208, value : 32'h20}, //phyinit_io_write: 0x44207, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44209, value : 32'h0}, //phyinit_io_write: 0x44208, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h4420a, value : 32'hc000080}, //phyinit_io_write: 0x44209, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4420b, value : 32'h1800}, //phyinit_io_write: 0x4420a, 0xc000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4420c, value : 32'h44520}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4420d, value : 32'h0}, //phyinit_io_write: 0x4420c, 0x44520
                          '{ step_type : REG_WRITE, reg_addr : 32'h4420e, value : 32'hc001c80}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 16
                          '{ step_type : REG_WRITE, reg_addr : 32'h4420f, value : 32'h1800}, //phyinit_io_write: 0x4420e, 0xc001c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44210, value : 32'h1020}, //phyinit_io_write: 0x4420f, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44211, value : 32'h0}, //phyinit_io_write: 0x44210, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h44212, value : 32'h1020}, //phyinit_io_write: 0x44211, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44213, value : 32'h0}, //phyinit_io_write: 0x44212, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h44214, value : 32'hc001880}, //phyinit_io_write: 0x44213, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44215, value : 32'h1800}, //phyinit_io_write: 0x44214, 0xc001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44216, value : 32'h1020}, //phyinit_io_write: 0x44215, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44217, value : 32'h0}, //phyinit_io_write: 0x44216, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h44218, value : 32'h1020}, //phyinit_io_write: 0x44217, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44219, value : 32'h0}, //phyinit_io_write: 0x44218, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h4421a, value : 32'h1020}, //phyinit_io_write: 0x44219, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4421b, value : 32'h0}, //phyinit_io_write: 0x4421a, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h4421c, value : 32'hc001080}, //phyinit_io_write: 0x4421b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4421d, value : 32'h1800}, //phyinit_io_write: 0x4421c, 0xc001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4421e, value : 32'h44520}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4421f, value : 32'h0}, //phyinit_io_write: 0x4421e, 0x44520
                          '{ step_type : REG_WRITE, reg_addr : 32'h44220, value : 32'h80}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44221, value : 32'h1800}, //phyinit_io_write: 0x44220, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44222, value : 32'h200600}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44223, value : 32'h20}, //phyinit_io_write: 0x44222, 0x200600
                          '{ step_type : REG_WRITE, reg_addr : 32'h44224, value : 32'h49d60}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 40
                          '{ step_type : REG_WRITE, reg_addr : 32'h44225, value : 32'h0}, //phyinit_io_write: 0x44224, 0x49d60
                          '{ step_type : REG_WRITE, reg_addr : 32'h44226, value : 32'h18000080}, //phyinit_io_write: 0x44225, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44227, value : 32'h3bc1}, //phyinit_io_write: 0x44226, 0x18000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44228, value : 32'h1c000080}, //phyinit_io_write: 0x44227, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44229, value : 32'h3bc1}, //phyinit_io_write: 0x44228, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4422a, value : 32'h20000080}, //phyinit_io_write: 0x44229, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4422b, value : 32'h3bc1}, //phyinit_io_write: 0x4422a, 0x20000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4422c, value : 32'h24000080}, //phyinit_io_write: 0x4422b, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4422d, value : 32'h3bc1}, //phyinit_io_write: 0x4422c, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4422e, value : 32'h28000080}, //phyinit_io_write: 0x4422d, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4422f, value : 32'h3bc1}, //phyinit_io_write: 0x4422e, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44230, value : 32'h2c000880}, //phyinit_io_write: 0x4422f, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44231, value : 32'h3801}, //phyinit_io_write: 0x44230, 0x2c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44232, value : 32'h2c001080}, //phyinit_io_write: 0x44231, 0x3801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44233, value : 32'h3841}, //phyinit_io_write: 0x44232, 0x2c001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44234, value : 32'h2c000880}, //phyinit_io_write: 0x44233, 0x3841
                          '{ step_type : REG_WRITE, reg_addr : 32'h44235, value : 32'h3881}, //phyinit_io_write: 0x44234, 0x2c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44236, value : 32'h2c001080}, //phyinit_io_write: 0x44235, 0x3881
                          '{ step_type : REG_WRITE, reg_addr : 32'h44237, value : 32'h38c1}, //phyinit_io_write: 0x44236, 0x2c001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44238, value : 32'h2c000880}, //phyinit_io_write: 0x44237, 0x38c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44239, value : 32'h3901}, //phyinit_io_write: 0x44238, 0x2c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4423a, value : 32'h2c001080}, //phyinit_io_write: 0x44239, 0x3901
                          '{ step_type : REG_WRITE, reg_addr : 32'h4423b, value : 32'h3941}, //phyinit_io_write: 0x4423a, 0x2c001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4423c, value : 32'h2c000880}, //phyinit_io_write: 0x4423b, 0x3941
                          '{ step_type : REG_WRITE, reg_addr : 32'h4423d, value : 32'h3981}, //phyinit_io_write: 0x4423c, 0x2c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4423e, value : 32'h2c001080}, //phyinit_io_write: 0x4423d, 0x3981
                          '{ step_type : REG_WRITE, reg_addr : 32'h4423f, value : 32'h39c1}, //phyinit_io_write: 0x4423e, 0x2c001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44240, value : 32'h2000600}, //phyinit_io_write: 0x4423f, 0x39c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44241, value : 32'h200}, //phyinit_io_write: 0x44240, 0x2000600
                          '{ step_type : REG_WRITE, reg_addr : 32'h44242, value : 32'h2c0010c0}, //phyinit_io_write: 0x44241, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h44243, value : 32'h3bc1}, //phyinit_io_write: 0x44242, 0x2c0010c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44244, value : 32'h58000080}, //phyinit_io_write: 0x44243, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44245, value : 32'h3cf}, //phyinit_io_write: 0x44244, 0x58000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44246, value : 32'h5c000080}, //phyinit_io_write: 0x44245, 0x3cf
                          '{ step_type : REG_WRITE, reg_addr : 32'h44247, value : 32'h3cf}, //phyinit_io_write: 0x44246, 0x5c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44248, value : 32'h5c000880}, //phyinit_io_write: 0x44247, 0x3cf
                          '{ step_type : REG_WRITE, reg_addr : 32'h44249, value : 32'hcf}, //phyinit_io_write: 0x44248, 0x5c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4424a, value : 32'h5c000880}, //phyinit_io_write: 0x44249, 0xcf
                          '{ step_type : REG_WRITE, reg_addr : 32'h4424b, value : 32'h28f}, //phyinit_io_write: 0x4424a, 0x5c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4424c, value : 32'h52920}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4424d, value : 32'h0}, //phyinit_io_write: 0x4424c, 0x52920
                          '{ step_type : REG_WRITE, reg_addr : 32'h4424e, value : 32'h18000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 70
                          '{ step_type : REG_WRITE, reg_addr : 32'h4424f, value : 32'h3801}, //phyinit_io_write: 0x4424e, 0x18000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44250, value : 32'h18000080}, //phyinit_io_write: 0x4424f, 0x3801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44251, value : 32'h3841}, //phyinit_io_write: 0x44250, 0x18000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44252, value : 32'h18000080}, //phyinit_io_write: 0x44251, 0x3841
                          '{ step_type : REG_WRITE, reg_addr : 32'h44253, value : 32'h3881}, //phyinit_io_write: 0x44252, 0x18000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44254, value : 32'h18000080}, //phyinit_io_write: 0x44253, 0x3881
                          '{ step_type : REG_WRITE, reg_addr : 32'h44255, value : 32'h38c1}, //phyinit_io_write: 0x44254, 0x18000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44256, value : 32'h1c000080}, //phyinit_io_write: 0x44255, 0x38c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44257, value : 32'h3801}, //phyinit_io_write: 0x44256, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44258, value : 32'h1c000080}, //phyinit_io_write: 0x44257, 0x3801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44259, value : 32'h3841}, //phyinit_io_write: 0x44258, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4425a, value : 32'h1c000080}, //phyinit_io_write: 0x44259, 0x3841
                          '{ step_type : REG_WRITE, reg_addr : 32'h4425b, value : 32'h3881}, //phyinit_io_write: 0x4425a, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4425c, value : 32'h1c000080}, //phyinit_io_write: 0x4425b, 0x3881
                          '{ step_type : REG_WRITE, reg_addr : 32'h4425d, value : 32'h38c1}, //phyinit_io_write: 0x4425c, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4425e, value : 32'h20000080}, //phyinit_io_write: 0x4425d, 0x38c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4425f, value : 32'h3801}, //phyinit_io_write: 0x4425e, 0x20000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44260, value : 32'h20000080}, //phyinit_io_write: 0x4425f, 0x3801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44261, value : 32'h3841}, //phyinit_io_write: 0x44260, 0x20000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44262, value : 32'h20000080}, //phyinit_io_write: 0x44261, 0x3841
                          '{ step_type : REG_WRITE, reg_addr : 32'h44263, value : 32'h3881}, //phyinit_io_write: 0x44262, 0x20000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44264, value : 32'h20000080}, //phyinit_io_write: 0x44263, 0x3881
                          '{ step_type : REG_WRITE, reg_addr : 32'h44265, value : 32'h38c1}, //phyinit_io_write: 0x44264, 0x20000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44266, value : 32'h24000080}, //phyinit_io_write: 0x44265, 0x38c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44267, value : 32'h3801}, //phyinit_io_write: 0x44266, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44268, value : 32'h24000080}, //phyinit_io_write: 0x44267, 0x3801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44269, value : 32'h3841}, //phyinit_io_write: 0x44268, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4426a, value : 32'h24000080}, //phyinit_io_write: 0x44269, 0x3841
                          '{ step_type : REG_WRITE, reg_addr : 32'h4426b, value : 32'h3881}, //phyinit_io_write: 0x4426a, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4426c, value : 32'h24000080}, //phyinit_io_write: 0x4426b, 0x3881
                          '{ step_type : REG_WRITE, reg_addr : 32'h4426d, value : 32'h38c1}, //phyinit_io_write: 0x4426c, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4426e, value : 32'h28000080}, //phyinit_io_write: 0x4426d, 0x38c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4426f, value : 32'h3841}, //phyinit_io_write: 0x4426e, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44270, value : 32'h28000080}, //phyinit_io_write: 0x4426f, 0x3841
                          '{ step_type : REG_WRITE, reg_addr : 32'h44271, value : 32'h38c1}, //phyinit_io_write: 0x44270, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44272, value : 32'h2c000880}, //phyinit_io_write: 0x44271, 0x38c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44273, value : 32'h3801}, //phyinit_io_write: 0x44272, 0x2c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44274, value : 32'h2c001080}, //phyinit_io_write: 0x44273, 0x3801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44275, value : 32'h3841}, //phyinit_io_write: 0x44274, 0x2c001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44276, value : 32'h2c000880}, //phyinit_io_write: 0x44275, 0x3841
                          '{ step_type : REG_WRITE, reg_addr : 32'h44277, value : 32'h3881}, //phyinit_io_write: 0x44276, 0x2c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44278, value : 32'h2c001080}, //phyinit_io_write: 0x44277, 0x3881
                          '{ step_type : REG_WRITE, reg_addr : 32'h44279, value : 32'h38c1}, //phyinit_io_write: 0x44278, 0x2c001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4427a, value : 32'h2000600}, //phyinit_io_write: 0x44279, 0x38c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4427b, value : 32'h200}, //phyinit_io_write: 0x4427a, 0x2000600
                          '{ step_type : REG_WRITE, reg_addr : 32'h4427c, value : 32'h2c0010c0}, //phyinit_io_write: 0x4427b, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h4427d, value : 32'h3bc1}, //phyinit_io_write: 0x4427c, 0x2c0010c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4427e, value : 32'h58000080}, //phyinit_io_write: 0x4427d, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4427f, value : 32'hf}, //phyinit_io_write: 0x4427e, 0x58000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44280, value : 32'h5c000080}, //phyinit_io_write: 0x4427f, 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h44281, value : 32'hf}, //phyinit_io_write: 0x44280, 0x5c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44282, value : 32'h58000080}, //phyinit_io_write: 0x44281, 0xf
                          '{ step_type : REG_WRITE, reg_addr : 32'h44283, value : 32'h4f}, //phyinit_io_write: 0x44282, 0x58000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44284, value : 32'h5c000080}, //phyinit_io_write: 0x44283, 0x4f
                          '{ step_type : REG_WRITE, reg_addr : 32'h44285, value : 32'h4f}, //phyinit_io_write: 0x44284, 0x5c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44286, value : 32'h58000080}, //phyinit_io_write: 0x44285, 0x4f
                          '{ step_type : REG_WRITE, reg_addr : 32'h44287, value : 32'h8f}, //phyinit_io_write: 0x44286, 0x58000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44288, value : 32'h5c000080}, //phyinit_io_write: 0x44287, 0x8f
                          '{ step_type : REG_WRITE, reg_addr : 32'h44289, value : 32'h8f}, //phyinit_io_write: 0x44288, 0x5c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4428a, value : 32'h58000080}, //phyinit_io_write: 0x44289, 0x8f
                          '{ step_type : REG_WRITE, reg_addr : 32'h4428b, value : 32'hcf}, //phyinit_io_write: 0x4428a, 0x58000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4428c, value : 32'h58000080}, //phyinit_io_write: 0x4428b, 0xcf
                          '{ step_type : REG_WRITE, reg_addr : 32'h4428d, value : 32'h10f}, //phyinit_io_write: 0x4428c, 0x58000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4428e, value : 32'h5c000080}, //phyinit_io_write: 0x4428d, 0x10f
                          '{ step_type : REG_WRITE, reg_addr : 32'h4428f, value : 32'h10f}, //phyinit_io_write: 0x4428e, 0x5c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44290, value : 32'h58000080}, //phyinit_io_write: 0x4428f, 0x10f
                          '{ step_type : REG_WRITE, reg_addr : 32'h44291, value : 32'h14f}, //phyinit_io_write: 0x44290, 0x58000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44292, value : 32'h5c000080}, //phyinit_io_write: 0x44291, 0x14f
                          '{ step_type : REG_WRITE, reg_addr : 32'h44293, value : 32'h14f}, //phyinit_io_write: 0x44292, 0x5c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44294, value : 32'h20000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44295, value : 32'h2bcc}, //phyinit_io_write: 0x44294, 0x20000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44296, value : 32'h53931}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44297, value : 32'h0}, //phyinit_io_write: 0x44296, 0x53931
                          '{ step_type : REG_WRITE, reg_addr : 32'h44298, value : 32'h40001a00}, //phyinit_io_write: 0x44297, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44299, value : 32'h0}, //phyinit_io_write: 0x44298, 0x40001a00
                          '{ step_type : REG_WRITE, reg_addr : 32'h4429a, value : 32'h53960}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4429b, value : 32'h0}, //phyinit_io_write: 0x4429a, 0x53960
                          '{ step_type : REG_WRITE, reg_addr : 32'h4429c, value : 32'h40030a0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 34
                          '{ step_type : REG_WRITE, reg_addr : 32'h4429d, value : 32'h2c00}, //phyinit_io_write: 0x4429c, 0x40030a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4429e, value : 32'h88000080}, //phyinit_io_write: 0x4429d, 0x2c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h4429f, value : 32'h802}, //phyinit_io_write: 0x4429e, 0x88000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a0, value : 32'h5c1ffc80}, //phyinit_io_write: 0x4429f, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a1, value : 32'h7c2}, //phyinit_io_write: 0x442a0, 0x5c1ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a2, value : 32'h800600}, //phyinit_io_write: 0x442a1, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a3, value : 32'h80}, //phyinit_io_write: 0x442a2, 0x800600
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a4, value : 32'hbc000900}, //phyinit_io_write: 0x442a3, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a5, value : 32'h16c0c}, //phyinit_io_write: 0x442a4, 0xbc000900
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a6, value : 32'h40000c0}, //phyinit_io_write: 0x442a5, 0x16c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a7, value : 32'h2424}, //phyinit_io_write: 0x442a6, 0x40000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a8, value : 32'h40080e0}, //phyinit_io_write: 0x442a7, 0x2424
                          '{ step_type : REG_WRITE, reg_addr : 32'h442a9, value : 32'h2424}, //phyinit_io_write: 0x442a8, 0x40080e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442aa, value : 32'h4000000}, //phyinit_io_write: 0x442a9, 0x2424
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ab, value : 32'h0}, //phyinit_io_write: 0x442aa, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ac, value : 32'h98001cb5}, //phyinit_io_write: 0x442ab, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ad, value : 32'h2c0c}, //phyinit_io_write: 0x442ac, 0x98001cb5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ae, value : 32'h9c0020b5}, //phyinit_io_write: 0x442ad, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442af, value : 32'h2c0c}, //phyinit_io_write: 0x442ae, 0x9c0020b5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b0, value : 32'h98000095}, //phyinit_io_write: 0x442af, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b1, value : 32'h2c0c}, //phyinit_io_write: 0x442b0, 0x98000095
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b2, value : 32'h9c000095}, //phyinit_io_write: 0x442b1, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b3, value : 32'h2c0c}, //phyinit_io_write: 0x442b2, 0x9c000095
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b4, value : 32'h40000095}, //phyinit_io_write: 0x442b3, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b5, value : 32'h2c0c}, //phyinit_io_write: 0x442b4, 0x40000095
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b6, value : 32'h605}, //phyinit_io_write: 0x442b5, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b7, value : 32'h2000}, //phyinit_io_write: 0x442b6, 0x605
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b8, value : 32'h400000c5}, //phyinit_io_write: 0x442b7, 0x2000
                          '{ step_type : REG_WRITE, reg_addr : 32'h442b9, value : 32'h2c0c}, //phyinit_io_write: 0x442b8, 0x400000c5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ba, value : 32'h800004c5}, //phyinit_io_write: 0x442b9, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442bb, value : 32'h2c0c}, //phyinit_io_write: 0x442ba, 0x800004c5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442bc, value : 32'h800000c5}, //phyinit_io_write: 0x442bb, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442bd, value : 32'h2c0c}, //phyinit_io_write: 0x442bc, 0x800000c5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442be, value : 32'h40000e5}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 18
                          '{ step_type : REG_WRITE, reg_addr : 32'h442bf, value : 32'h2c00}, //phyinit_io_write: 0x442be, 0x40000e5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c0, value : 32'hbc0000e5}, //phyinit_io_write: 0x442bf, 0x2c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c1, value : 32'h16c0c}, //phyinit_io_write: 0x442c0, 0xbc0000e5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c2, value : 32'h4000000}, //phyinit_io_write: 0x442c1, 0x16c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c3, value : 32'h0}, //phyinit_io_write: 0x442c2, 0x4000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c4, value : 32'h9bfe04e5}, //phyinit_io_write: 0x442c3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c5, value : 32'h2c0c}, //phyinit_io_write: 0x442c4, 0x9bfe04e5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c6, value : 32'h9ffe04e5}, //phyinit_io_write: 0x442c5, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c7, value : 32'h2c0c}, //phyinit_io_write: 0x442c6, 0x9ffe04e5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c8, value : 32'h9bfe00e5}, //phyinit_io_write: 0x442c7, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442c9, value : 32'h2c0c}, //phyinit_io_write: 0x442c8, 0x9bfe00e5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ca, value : 32'h9ffe00e5}, //phyinit_io_write: 0x442c9, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442cb, value : 32'h2c0c}, //phyinit_io_write: 0x442ca, 0x9ffe00e5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442cc, value : 32'h400004e5}, //phyinit_io_write: 0x442cb, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442cd, value : 32'h2c0c}, //phyinit_io_write: 0x442cc, 0x400004e5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ce, value : 32'h4000400}, //phyinit_io_write: 0x442cd, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442cf, value : 32'h0}, //phyinit_io_write: 0x442ce, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d0, value : 32'hbc0008a5}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d1, value : 32'h16c0c}, //phyinit_io_write: 0x442d0, 0xbc0008a5
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d2, value : 32'h1e0}, //phyinit_io_write: 0x442d1, 0x16c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d3, value : 32'h0}, //phyinit_io_write: 0x442d2, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d4, value : 32'he8030c80}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d5, value : 32'h1c01}, //phyinit_io_write: 0x442d4, 0xe8030c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d6, value : 32'h4000400}, //phyinit_io_write: 0x442d5, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d7, value : 32'h0}, //phyinit_io_write: 0x442d6, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d8, value : 32'he8000080}, //phyinit_io_write: 0x442d7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442d9, value : 32'h1c01}, //phyinit_io_write: 0x442d8, 0xe8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h442da, value : 32'h1e0}, //phyinit_io_write: 0x442d9, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h442db, value : 32'h0}, //phyinit_io_write: 0x442da, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442dc, value : 32'h88000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 40
                          '{ step_type : REG_WRITE, reg_addr : 32'h442dd, value : 32'h802}, //phyinit_io_write: 0x442dc, 0x88000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h442de, value : 32'h4000c00}, //phyinit_io_write: 0x442dd, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h442df, value : 32'h0}, //phyinit_io_write: 0x442de, 0x4000c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e0, value : 32'hcc80}, //phyinit_io_write: 0x442df, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e1, value : 32'h808}, //phyinit_io_write: 0x442e0, 0xcc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e2, value : 32'h1c000480}, //phyinit_io_write: 0x442e1, 0x808
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e3, value : 32'hfc1}, //phyinit_io_write: 0x442e2, 0x1c000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e4, value : 32'h1c000080}, //phyinit_io_write: 0x442e3, 0xfc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e5, value : 32'hfc1}, //phyinit_io_write: 0x442e4, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e6, value : 32'h1c000480}, //phyinit_io_write: 0x442e5, 0xfc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e7, value : 32'h7c1}, //phyinit_io_write: 0x442e6, 0x1c000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e8, value : 32'h1c000080}, //phyinit_io_write: 0x442e7, 0x7c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h442e9, value : 32'h7c1}, //phyinit_io_write: 0x442e8, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ea, value : 32'h80}, //phyinit_io_write: 0x442e9, 0x7c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h442eb, value : 32'h808}, //phyinit_io_write: 0x442ea, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ec, value : 32'h50000080}, //phyinit_io_write: 0x442eb, 0x808
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ed, value : 32'h1c01}, //phyinit_io_write: 0x442ec, 0x50000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ee, value : 32'hb8000480}, //phyinit_io_write: 0x442ed, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ef, value : 32'h801}, //phyinit_io_write: 0x442ee, 0xb8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f0, value : 32'h4000400}, //phyinit_io_write: 0x442ef, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f1, value : 32'h0}, //phyinit_io_write: 0x442f0, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f2, value : 32'h40600}, //phyinit_io_write: 0x442f1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f3, value : 32'h4}, //phyinit_io_write: 0x442f2, 0x40600
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f4, value : 32'h598000e0}, //phyinit_io_write: 0x442f3, 0x4
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f5, value : 32'h7c0}, //phyinit_io_write: 0x442f4, 0x598000e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f6, value : 32'h28000480}, //phyinit_io_write: 0x442f5, 0x7c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f7, value : 32'hfc0}, //phyinit_io_write: 0x442f6, 0x28000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f8, value : 32'h4001000}, //phyinit_io_write: 0x442f7, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442f9, value : 32'h0}, //phyinit_io_write: 0x442f8, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h442fa, value : 32'he0000080}, //phyinit_io_write: 0x442f9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442fb, value : 32'h803}, //phyinit_io_write: 0x442fa, 0xe0000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h442fc, value : 32'h4001400}, //phyinit_io_write: 0x442fb, 0x803
                          '{ step_type : REG_WRITE, reg_addr : 32'h442fd, value : 32'h0}, //phyinit_io_write: 0x442fc, 0x4001400
                          '{ step_type : REG_WRITE, reg_addr : 32'h442fe, value : 32'h88000880}, //phyinit_io_write: 0x442fd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h442ff, value : 32'h802}, //phyinit_io_write: 0x442fe, 0x88000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44300, value : 32'hc20}, //phyinit_io_write: 0x442ff, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h44301, value : 32'h0}, //phyinit_io_write: 0x44300, 0xc20
                          '{ step_type : REG_WRITE, reg_addr : 32'h44302, value : 32'h40004600}, //phyinit_io_write: 0x44301, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44303, value : 32'h0}, //phyinit_io_write: 0x44302, 0x40004600
                          '{ step_type : REG_WRITE, reg_addr : 32'h44304, value : 32'h60d60}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44305, value : 32'h0}, //phyinit_io_write: 0x44304, 0x60d60
                          '{ step_type : REG_WRITE, reg_addr : 32'h44306, value : 32'h1c000880}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 12
                          '{ step_type : REG_WRITE, reg_addr : 32'h44307, value : 32'hfc1}, //phyinit_io_write: 0x44306, 0x1c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44308, value : 32'h1c000080}, //phyinit_io_write: 0x44307, 0xfc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44309, value : 32'hfc1}, //phyinit_io_write: 0x44308, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4430a, value : 32'h1c000880}, //phyinit_io_write: 0x44309, 0xfc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4430b, value : 32'h7c1}, //phyinit_io_write: 0x4430a, 0x1c000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4430c, value : 32'h1c000080}, //phyinit_io_write: 0x4430b, 0x7c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4430d, value : 32'h7c1}, //phyinit_io_write: 0x4430c, 0x1c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4430e, value : 32'h4003c00}, //phyinit_io_write: 0x4430d, 0x7c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4430f, value : 32'h0}, //phyinit_io_write: 0x4430e, 0x4003c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h44310, value : 32'h40600}, //phyinit_io_write: 0x4430f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44311, value : 32'h4}, //phyinit_io_write: 0x44310, 0x40600
                          '{ step_type : REG_WRITE, reg_addr : 32'h44312, value : 32'h62d40}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44313, value : 32'h0}, //phyinit_io_write: 0x44312, 0x62d40
                          '{ step_type : REG_WRITE, reg_addr : 32'h44314, value : 32'h1b9c0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44315, value : 32'h0}, //phyinit_io_write: 0x44314, 0x1b9c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44316, value : 32'h28000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 14
                          '{ step_type : REG_WRITE, reg_addr : 32'h44317, value : 32'hfc0}, //phyinit_io_write: 0x44316, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44318, value : 32'h80000080}, //phyinit_io_write: 0x44317, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44319, value : 32'hfc2}, //phyinit_io_write: 0x44318, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4431a, value : 32'h98000080}, //phyinit_io_write: 0x44319, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4431b, value : 32'hfc2}, //phyinit_io_write: 0x4431a, 0x98000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4431c, value : 32'h24000080}, //phyinit_io_write: 0x4431b, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4431d, value : 32'h7c2}, //phyinit_io_write: 0x4431c, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4431e, value : 32'h28000080}, //phyinit_io_write: 0x4431d, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4431f, value : 32'h7c2}, //phyinit_io_write: 0x4431e, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44320, value : 32'h883c0080}, //phyinit_io_write: 0x4431f, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44321, value : 32'hfc2}, //phyinit_io_write: 0x44320, 0x883c0080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44322, value : 32'h80040200}, //phyinit_io_write: 0x44321, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44323, value : 32'h400f}, //phyinit_io_write: 0x44322, 0x80040200
                          '{ step_type : REG_WRITE, reg_addr : 32'h44324, value : 32'h66540}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44325, value : 32'h0}, //phyinit_io_write: 0x44324, 0x66540
                          '{ step_type : REG_WRITE, reg_addr : 32'h44326, value : 32'h80200}, //phyinit_io_write: 0x44325, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44327, value : 32'h400e}, //phyinit_io_write: 0x44326, 0x80200
                          '{ step_type : REG_WRITE, reg_addr : 32'h44328, value : 32'h66540}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 10
                          '{ step_type : REG_WRITE, reg_addr : 32'h44329, value : 32'h0}, //phyinit_io_write: 0x44328, 0x66540
                          '{ step_type : REG_WRITE, reg_addr : 32'h4432a, value : 32'he4000480}, //phyinit_io_write: 0x44329, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4432b, value : 32'h801}, //phyinit_io_write: 0x4432a, 0xe4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4432c, value : 32'h4000800}, //phyinit_io_write: 0x4432b, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h4432d, value : 32'h0}, //phyinit_io_write: 0x4432c, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4432e, value : 32'he4000080}, //phyinit_io_write: 0x4432d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4432f, value : 32'h801}, //phyinit_io_write: 0x4432e, 0xe4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44330, value : 32'h4000800}, //phyinit_io_write: 0x4432f, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44331, value : 32'h0}, //phyinit_io_write: 0x44330, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44332, value : 32'he8030c81}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 10
                          '{ step_type : REG_WRITE, reg_addr : 32'h44333, value : 32'h1c01}, //phyinit_io_write: 0x44332, 0xe8030c81
                          '{ step_type : REG_WRITE, reg_addr : 32'h44334, value : 32'h4000800}, //phyinit_io_write: 0x44333, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44335, value : 32'h0}, //phyinit_io_write: 0x44334, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44336, value : 32'he8000081}, //phyinit_io_write: 0x44335, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44337, value : 32'h1c01}, //phyinit_io_write: 0x44336, 0xe8000081
                          '{ step_type : REG_WRITE, reg_addr : 32'h44338, value : 32'h4000400}, //phyinit_io_write: 0x44337, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44339, value : 32'h0}, //phyinit_io_write: 0x44338, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4433a, value : 32'h40001a01}, //phyinit_io_write: 0x44339, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4433b, value : 32'h0}, //phyinit_io_write: 0x4433a, 0x40001a01
                          '{ step_type : REG_WRITE, reg_addr : 32'h4433c, value : 32'h69141}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4433d, value : 32'h0}, //phyinit_io_write: 0x4433c, 0x69141
                          '{ step_type : REG_WRITE, reg_addr : 32'h4433e, value : 32'ha0000481}, //phyinit_io_write: 0x4433d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4433f, value : 32'h2420}, //phyinit_io_write: 0x4433e, 0xa0000481
                          '{ step_type : REG_WRITE, reg_addr : 32'h44340, value : 32'h4000400}, //phyinit_io_write: 0x4433f, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h44341, value : 32'h0}, //phyinit_io_write: 0x44340, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44342, value : 32'h40003201}, //phyinit_io_write: 0x44341, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44343, value : 32'h0}, //phyinit_io_write: 0x44342, 0x40003201
                          '{ step_type : REG_WRITE, reg_addr : 32'h44344, value : 32'h6b141}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44345, value : 32'h0}, //phyinit_io_write: 0x44344, 0x6b141
                          '{ step_type : REG_WRITE, reg_addr : 32'h44346, value : 32'h69161}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44347, value : 32'h0}, //phyinit_io_write: 0x44346, 0x69161
                          '{ step_type : REG_WRITE, reg_addr : 32'h44348, value : 32'h1c21}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 16
                          '{ step_type : REG_WRITE, reg_addr : 32'h44349, value : 32'h0}, //phyinit_io_write: 0x44348, 0x1c21
                          '{ step_type : REG_WRITE, reg_addr : 32'h4434a, value : 32'ha0000081}, //phyinit_io_write: 0x44349, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4434b, value : 32'h2420}, //phyinit_io_write: 0x4434a, 0xa0000081
                          '{ step_type : REG_WRITE, reg_addr : 32'h4434c, value : 32'h4000400}, //phyinit_io_write: 0x4434b, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h4434d, value : 32'h0}, //phyinit_io_write: 0x4434c, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4434e, value : 32'h20601}, //phyinit_io_write: 0x4434d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4434f, value : 32'h2}, //phyinit_io_write: 0x4434e, 0x20601
                          '{ step_type : REG_WRITE, reg_addr : 32'h44350, value : 32'he8030cc1}, //phyinit_io_write: 0x4434f, 0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44351, value : 32'h1c01}, //phyinit_io_write: 0x44350, 0xe8030cc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44352, value : 32'h4000800}, //phyinit_io_write: 0x44351, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44353, value : 32'h0}, //phyinit_io_write: 0x44352, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44354, value : 32'he80000c1}, //phyinit_io_write: 0x44353, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44355, value : 32'h1c01}, //phyinit_io_write: 0x44354, 0xe80000c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44356, value : 32'h4000400}, //phyinit_io_write: 0x44355, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44357, value : 32'h0}, //phyinit_io_write: 0x44356, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44358, value : 32'ha0000081}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 16
                          '{ step_type : REG_WRITE, reg_addr : 32'h44359, value : 32'h2420}, //phyinit_io_write: 0x44358, 0xa0000081
                          '{ step_type : REG_WRITE, reg_addr : 32'h4435a, value : 32'h4000400}, //phyinit_io_write: 0x44359, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h4435b, value : 32'h0}, //phyinit_io_write: 0x4435a, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4435c, value : 32'he8030c91}, //phyinit_io_write: 0x4435b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4435d, value : 32'h1c01}, //phyinit_io_write: 0x4435c, 0xe8030c91
                          '{ step_type : REG_WRITE, reg_addr : 32'h4435e, value : 32'h4000800}, //phyinit_io_write: 0x4435d, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h4435f, value : 32'h0}, //phyinit_io_write: 0x4435e, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44360, value : 32'he8000091}, //phyinit_io_write: 0x4435f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44361, value : 32'h1c01}, //phyinit_io_write: 0x44360, 0xe8000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h44362, value : 32'h4000400}, //phyinit_io_write: 0x44361, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44363, value : 32'h0}, //phyinit_io_write: 0x44362, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44364, value : 32'ha8000480}, //phyinit_io_write: 0x44363, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44365, value : 32'h1c04}, //phyinit_io_write: 0x44364, 0xa8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44366, value : 32'h4000400}, //phyinit_io_write: 0x44365, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44367, value : 32'h0}, //phyinit_io_write: 0x44366, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44368, value : 32'h18000081}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44369, value : 32'h1e420}, //phyinit_io_write: 0x44368, 0x18000081
                          '{ step_type : REG_WRITE, reg_addr : 32'h4436a, value : 32'h40006611}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4436b, value : 32'h0}, //phyinit_io_write: 0x4436a, 0x40006611
                          '{ step_type : REG_WRITE, reg_addr : 32'h4436c, value : 32'h6e151}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4436d, value : 32'h0}, //phyinit_io_write: 0x4436c, 0x6e151
                          '{ step_type : REG_WRITE, reg_addr : 32'h4436e, value : 32'h21d1}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4436f, value : 32'h0}, //phyinit_io_write: 0x4436e, 0x21d1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44370, value : 32'ha0000491}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 12
                          '{ step_type : REG_WRITE, reg_addr : 32'h44371, value : 32'h2420}, //phyinit_io_write: 0x44370, 0xa0000491
                          '{ step_type : REG_WRITE, reg_addr : 32'h44372, value : 32'h4000400}, //phyinit_io_write: 0x44371, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h44373, value : 32'h0}, //phyinit_io_write: 0x44372, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44374, value : 32'h540020b1}, //phyinit_io_write: 0x44373, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44375, value : 32'h14fc0}, //phyinit_io_write: 0x44374, 0x540020b1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44376, value : 32'hf00024b1}, //phyinit_io_write: 0x44375, 0x14fc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44377, value : 32'h147c1}, //phyinit_io_write: 0x44376, 0xf00024b1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44378, value : 32'ha0000091}, //phyinit_io_write: 0x44377, 0x147c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44379, value : 32'h2420}, //phyinit_io_write: 0x44378, 0xa0000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h4437a, value : 32'h1e0}, //phyinit_io_write: 0x44379, 0x2420
                          '{ step_type : REG_WRITE, reg_addr : 32'h4437b, value : 32'h0}, //phyinit_io_write: 0x4437a, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4437c, value : 32'ha8000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 30
                          '{ step_type : REG_WRITE, reg_addr : 32'h4437d, value : 32'h1c06}, //phyinit_io_write: 0x4437c, 0xa8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4437e, value : 32'h80013080}, //phyinit_io_write: 0x4437d, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h4437f, value : 32'h1c04}, //phyinit_io_write: 0x4437e, 0x80013080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44380, value : 32'h4000400}, //phyinit_io_write: 0x4437f, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44381, value : 32'h0}, //phyinit_io_write: 0x44380, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44382, value : 32'h80013480}, //phyinit_io_write: 0x44381, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44383, value : 32'h1c04}, //phyinit_io_write: 0x44382, 0x80013480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44384, value : 32'h4000800}, //phyinit_io_write: 0x44383, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44385, value : 32'h0}, //phyinit_io_write: 0x44384, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44386, value : 32'h4001c00}, //phyinit_io_write: 0x44385, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44387, value : 32'h0}, //phyinit_io_write: 0x44386, 0x4001c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h44388, value : 32'h80000080}, //phyinit_io_write: 0x44387, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44389, value : 32'h1c04}, //phyinit_io_write: 0x44388, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4438a, value : 32'h420}, //phyinit_io_write: 0x44389, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4438b, value : 32'h0}, //phyinit_io_write: 0x4438a, 0x420
                          '{ step_type : REG_WRITE, reg_addr : 32'h4438c, value : 32'ha8000080}, //phyinit_io_write: 0x4438b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4438d, value : 32'h1c06}, //phyinit_io_write: 0x4438c, 0xa8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4438e, value : 32'h80013880}, //phyinit_io_write: 0x4438d, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h4438f, value : 32'h1c04}, //phyinit_io_write: 0x4438e, 0x80013880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44390, value : 32'h4000400}, //phyinit_io_write: 0x4438f, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44391, value : 32'h0}, //phyinit_io_write: 0x44390, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44392, value : 32'h80013c80}, //phyinit_io_write: 0x44391, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44393, value : 32'h1c04}, //phyinit_io_write: 0x44392, 0x80013c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44394, value : 32'h4000800}, //phyinit_io_write: 0x44393, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44395, value : 32'h0}, //phyinit_io_write: 0x44394, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44396, value : 32'h4001c00}, //phyinit_io_write: 0x44395, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44397, value : 32'h0}, //phyinit_io_write: 0x44396, 0x4001c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h44398, value : 32'h80000080}, //phyinit_io_write: 0x44397, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44399, value : 32'h1c04}, //phyinit_io_write: 0x44398, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4439a, value : 32'h1e0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4439b, value : 32'h0}, //phyinit_io_write: 0x4439a, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4439c, value : 32'h20000086}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 176
                          '{ step_type : REG_WRITE, reg_addr : 32'h4439d, value : 32'h1c7c4}, //phyinit_io_write: 0x4439c, 0x20000086
                          '{ step_type : REG_WRITE, reg_addr : 32'h4439e, value : 32'h9e000480}, //phyinit_io_write: 0x4439d, 0x1c7c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4439f, value : 32'h7c2}, //phyinit_io_write: 0x4439e, 0x9e000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a0, value : 32'hc4060080}, //phyinit_io_write: 0x4439f, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a1, value : 32'h7c2}, //phyinit_io_write: 0x443a0, 0xc4060080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a2, value : 32'hd4000480}, //phyinit_io_write: 0x443a1, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a3, value : 32'h7c2}, //phyinit_io_write: 0x443a2, 0xd4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a4, value : 32'he4000480}, //phyinit_io_write: 0x443a3, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a5, value : 32'h7c2}, //phyinit_io_write: 0x443a4, 0xe4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a6, value : 32'h9c003080}, //phyinit_io_write: 0x443a5, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a7, value : 32'h1c04}, //phyinit_io_write: 0x443a6, 0x9c003080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a8, value : 32'h7c000080}, //phyinit_io_write: 0x443a7, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h443a9, value : 32'h1c7c1}, //phyinit_io_write: 0x443a8, 0x7c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443aa, value : 32'h88000c80}, //phyinit_io_write: 0x443a9, 0x1c7c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ab, value : 32'h7c2}, //phyinit_io_write: 0x443aa, 0x88000c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ac, value : 32'h64000c80}, //phyinit_io_write: 0x443ab, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ad, value : 32'h801}, //phyinit_io_write: 0x443ac, 0x64000c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ae, value : 32'h90000880}, //phyinit_io_write: 0x443ad, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h443af, value : 32'h7c2}, //phyinit_io_write: 0x443ae, 0x90000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b0, value : 32'hec0ffc80}, //phyinit_io_write: 0x443af, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b1, value : 32'h7c2}, //phyinit_io_write: 0x443b0, 0xec0ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b2, value : 32'hec000080}, //phyinit_io_write: 0x443b1, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b3, value : 32'h7c2}, //phyinit_io_write: 0x443b2, 0xec000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b4, value : 32'hf8000080}, //phyinit_io_write: 0x443b3, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b5, value : 32'h7fe}, //phyinit_io_write: 0x443b4, 0xf8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b6, value : 32'hf8000480}, //phyinit_io_write: 0x443b5, 0x7fe
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b7, value : 32'h7c2}, //phyinit_io_write: 0x443b6, 0xf8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b8, value : 32'hf8000480}, //phyinit_io_write: 0x443b7, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443b9, value : 32'h7d2}, //phyinit_io_write: 0x443b8, 0xf8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ba, value : 32'ha8001080}, //phyinit_io_write: 0x443b9, 0x7d2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443bb, value : 32'h1c06}, //phyinit_io_write: 0x443ba, 0xa8001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443bc, value : 32'h80014880}, //phyinit_io_write: 0x443bb, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h443bd, value : 32'h1c04}, //phyinit_io_write: 0x443bc, 0x80014880
                          '{ step_type : REG_WRITE, reg_addr : 32'h443be, value : 32'h4000400}, //phyinit_io_write: 0x443bd, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h443bf, value : 32'h0}, //phyinit_io_write: 0x443be, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c0, value : 32'h80014c80}, //phyinit_io_write: 0x443bf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c1, value : 32'h1c04}, //phyinit_io_write: 0x443c0, 0x80014c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c2, value : 32'h4000800}, //phyinit_io_write: 0x443c1, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c3, value : 32'h0}, //phyinit_io_write: 0x443c2, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c4, value : 32'h840}, //phyinit_io_write: 0x443c3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c5, value : 32'h6000}, //phyinit_io_write: 0x443c4, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c6, value : 32'h80000080}, //phyinit_io_write: 0x443c5, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c7, value : 32'h1c04}, //phyinit_io_write: 0x443c6, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c8, value : 32'hf8000080}, //phyinit_io_write: 0x443c7, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h443c9, value : 32'h7c2}, //phyinit_io_write: 0x443c8, 0xf8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ca, value : 32'hf8000080}, //phyinit_io_write: 0x443c9, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443cb, value : 32'h7d2}, //phyinit_io_write: 0x443ca, 0xf8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443cc, value : 32'hec0ffc80}, //phyinit_io_write: 0x443cb, 0x7d2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443cd, value : 32'h7c2}, //phyinit_io_write: 0x443cc, 0xec0ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ce, value : 32'hec000080}, //phyinit_io_write: 0x443cd, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443cf, value : 32'h7c2}, //phyinit_io_write: 0x443ce, 0xec000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d0, value : 32'hf8000480}, //phyinit_io_write: 0x443cf, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d1, value : 32'h7c6}, //phyinit_io_write: 0x443d0, 0xf8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d2, value : 32'hf8000480}, //phyinit_io_write: 0x443d1, 0x7c6
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d3, value : 32'h7d6}, //phyinit_io_write: 0x443d2, 0xf8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d4, value : 32'ha8001080}, //phyinit_io_write: 0x443d3, 0x7d6
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d5, value : 32'h1c06}, //phyinit_io_write: 0x443d4, 0xa8001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d6, value : 32'h80015080}, //phyinit_io_write: 0x443d5, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d7, value : 32'h1c04}, //phyinit_io_write: 0x443d6, 0x80015080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d8, value : 32'h4000400}, //phyinit_io_write: 0x443d7, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h443d9, value : 32'h0}, //phyinit_io_write: 0x443d8, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h443da, value : 32'h80015480}, //phyinit_io_write: 0x443d9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443db, value : 32'h1c04}, //phyinit_io_write: 0x443da, 0x80015480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443dc, value : 32'h4000800}, //phyinit_io_write: 0x443db, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h443dd, value : 32'h0}, //phyinit_io_write: 0x443dc, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h443de, value : 32'h840}, //phyinit_io_write: 0x443dd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443df, value : 32'h6000}, //phyinit_io_write: 0x443de, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e0, value : 32'h80000080}, //phyinit_io_write: 0x443df, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e1, value : 32'h1c04}, //phyinit_io_write: 0x443e0, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e2, value : 32'hf8000080}, //phyinit_io_write: 0x443e1, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e3, value : 32'h7c6}, //phyinit_io_write: 0x443e2, 0xf8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e4, value : 32'hf8000080}, //phyinit_io_write: 0x443e3, 0x7c6
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e5, value : 32'h7d6}, //phyinit_io_write: 0x443e4, 0xf8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e6, value : 32'h64000880}, //phyinit_io_write: 0x443e5, 0x7d6
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e7, value : 32'h801}, //phyinit_io_write: 0x443e6, 0x64000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e8, value : 32'h1420}, //phyinit_io_write: 0x443e7, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h443e9, value : 32'h0}, //phyinit_io_write: 0x443e8, 0x1420
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ea, value : 32'hc4000480}, //phyinit_io_write: 0x443e9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443eb, value : 32'h7c0}, //phyinit_io_write: 0x443ea, 0xc4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ec, value : 32'h4001000}, //phyinit_io_write: 0x443eb, 0x7c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ed, value : 32'h0}, //phyinit_io_write: 0x443ec, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ee, value : 32'hc4000080}, //phyinit_io_write: 0x443ed, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ef, value : 32'h7c0}, //phyinit_io_write: 0x443ee, 0xc4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f0, value : 32'h4000600}, //phyinit_io_write: 0x443ef, 0x7c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f1, value : 32'h400}, //phyinit_io_write: 0x443f0, 0x4000600
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f2, value : 32'h24c8c8c0}, //phyinit_io_write: 0x443f1, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f3, value : 32'h147c8}, //phyinit_io_write: 0x443f2, 0x24c8c8c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f4, value : 32'h80000480}, //phyinit_io_write: 0x443f3, 0x147c8
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f5, value : 32'h802}, //phyinit_io_write: 0x443f4, 0x80000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f6, value : 32'h4000400}, //phyinit_io_write: 0x443f5, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f7, value : 32'h0}, //phyinit_io_write: 0x443f6, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f8, value : 32'h80000080}, //phyinit_io_write: 0x443f7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h443f9, value : 32'h802}, //phyinit_io_write: 0x443f8, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443fa, value : 32'h90000080}, //phyinit_io_write: 0x443f9, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h443fb, value : 32'h7c2}, //phyinit_io_write: 0x443fa, 0x90000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h443fc, value : 32'h98000c80}, //phyinit_io_write: 0x443fb, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443fd, value : 32'h7c2}, //phyinit_io_write: 0x443fc, 0x98000c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h443fe, value : 32'ha8001080}, //phyinit_io_write: 0x443fd, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h443ff, value : 32'h1c06}, //phyinit_io_write: 0x443fe, 0xa8001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44400, value : 32'h80015880}, //phyinit_io_write: 0x443ff, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h44401, value : 32'h1c04}, //phyinit_io_write: 0x44400, 0x80015880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44402, value : 32'h4000400}, //phyinit_io_write: 0x44401, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44403, value : 32'h0}, //phyinit_io_write: 0x44402, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44404, value : 32'h80015c80}, //phyinit_io_write: 0x44403, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44405, value : 32'h1c04}, //phyinit_io_write: 0x44404, 0x80015c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44406, value : 32'h4000800}, //phyinit_io_write: 0x44405, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44407, value : 32'h0}, //phyinit_io_write: 0x44406, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44408, value : 32'h840}, //phyinit_io_write: 0x44407, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44409, value : 32'h6000}, //phyinit_io_write: 0x44408, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h4440a, value : 32'h80000080}, //phyinit_io_write: 0x44409, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4440b, value : 32'h1c04}, //phyinit_io_write: 0x4440a, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4440c, value : 32'h4000800}, //phyinit_io_write: 0x4440b, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4440d, value : 32'h0}, //phyinit_io_write: 0x4440c, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4440e, value : 32'h98000080}, //phyinit_io_write: 0x4440d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4440f, value : 32'h7c2}, //phyinit_io_write: 0x4440e, 0x98000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44410, value : 32'h88000080}, //phyinit_io_write: 0x4440f, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44411, value : 32'h7c2}, //phyinit_io_write: 0x44410, 0x88000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44412, value : 32'h64000080}, //phyinit_io_write: 0x44411, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44413, value : 32'h801}, //phyinit_io_write: 0x44412, 0x64000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44414, value : 32'h7c000480}, //phyinit_io_write: 0x44413, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44415, value : 32'h1c7c1}, //phyinit_io_write: 0x44414, 0x7c000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44416, value : 32'he4000480}, //phyinit_io_write: 0x44415, 0x1c7c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h44417, value : 32'h801}, //phyinit_io_write: 0x44416, 0xe4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44418, value : 32'h4000800}, //phyinit_io_write: 0x44417, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44419, value : 32'h0}, //phyinit_io_write: 0x44418, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4441a, value : 32'he4000080}, //phyinit_io_write: 0x44419, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4441b, value : 32'h801}, //phyinit_io_write: 0x4441a, 0xe4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4441c, value : 32'h4000800}, //phyinit_io_write: 0x4441b, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h4441d, value : 32'h0}, //phyinit_io_write: 0x4441c, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4441e, value : 32'h1820}, //phyinit_io_write: 0x4441d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4441f, value : 32'h0}, //phyinit_io_write: 0x4441e, 0x1820
                          '{ step_type : REG_WRITE, reg_addr : 32'h44420, value : 32'h90000480}, //phyinit_io_write: 0x4441f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44421, value : 32'h7c2}, //phyinit_io_write: 0x44420, 0x90000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44422, value : 32'ha8001080}, //phyinit_io_write: 0x44421, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44423, value : 32'h1c06}, //phyinit_io_write: 0x44422, 0xa8001080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44424, value : 32'h80016080}, //phyinit_io_write: 0x44423, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h44425, value : 32'h1c04}, //phyinit_io_write: 0x44424, 0x80016080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44426, value : 32'h4000400}, //phyinit_io_write: 0x44425, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44427, value : 32'h0}, //phyinit_io_write: 0x44426, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44428, value : 32'h80016480}, //phyinit_io_write: 0x44427, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44429, value : 32'h1c04}, //phyinit_io_write: 0x44428, 0x80016480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4442a, value : 32'h4000800}, //phyinit_io_write: 0x44429, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4442b, value : 32'h0}, //phyinit_io_write: 0x4442a, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4442c, value : 32'h840}, //phyinit_io_write: 0x4442b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4442d, value : 32'h6000}, //phyinit_io_write: 0x4442c, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h4442e, value : 32'h80000080}, //phyinit_io_write: 0x4442d, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4442f, value : 32'h1c04}, //phyinit_io_write: 0x4442e, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44430, value : 32'h4000800}, //phyinit_io_write: 0x4442f, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44431, value : 32'h0}, //phyinit_io_write: 0x44430, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44432, value : 32'h80000480}, //phyinit_io_write: 0x44431, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44433, value : 32'h802}, //phyinit_io_write: 0x44432, 0x80000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44434, value : 32'h4000400}, //phyinit_io_write: 0x44433, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h44435, value : 32'h0}, //phyinit_io_write: 0x44434, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44436, value : 32'h80000080}, //phyinit_io_write: 0x44435, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44437, value : 32'h802}, //phyinit_io_write: 0x44436, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44438, value : 32'h90000080}, //phyinit_io_write: 0x44437, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h44439, value : 32'h7c2}, //phyinit_io_write: 0x44438, 0x90000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4443a, value : 32'h4000800}, //phyinit_io_write: 0x44439, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4443b, value : 32'h0}, //phyinit_io_write: 0x4443a, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4443c, value : 32'he4000480}, //phyinit_io_write: 0x4443b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4443d, value : 32'h801}, //phyinit_io_write: 0x4443c, 0xe4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4443e, value : 32'h4000800}, //phyinit_io_write: 0x4443d, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h4443f, value : 32'h0}, //phyinit_io_write: 0x4443e, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44440, value : 32'he4000080}, //phyinit_io_write: 0x4443f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44441, value : 32'h801}, //phyinit_io_write: 0x44440, 0xe4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44442, value : 32'h4000800}, //phyinit_io_write: 0x44441, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44443, value : 32'h0}, //phyinit_io_write: 0x44442, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44444, value : 32'ha8000080}, //phyinit_io_write: 0x44443, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44445, value : 32'h1c04}, //phyinit_io_write: 0x44444, 0xa8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44446, value : 32'h50000480}, //phyinit_io_write: 0x44445, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44447, value : 32'h1c01}, //phyinit_io_write: 0x44446, 0x50000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44448, value : 32'h20000486}, //phyinit_io_write: 0x44447, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44449, value : 32'h1c7c4}, //phyinit_io_write: 0x44448, 0x20000486
                          '{ step_type : REG_WRITE, reg_addr : 32'h4444a, value : 32'h1e0}, //phyinit_io_write: 0x44449, 0x1c7c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4444b, value : 32'h0}, //phyinit_io_write: 0x4444a, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4444c, value : 32'h80008600}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4444d, value : 32'h0}, //phyinit_io_write: 0x4444c, 0x80008600
                          '{ step_type : REG_WRITE, reg_addr : 32'h4444e, value : 32'h8c160}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 18
                          '{ step_type : REG_WRITE, reg_addr : 32'h4444f, value : 32'h0}, //phyinit_io_write: 0x4444e, 0x8c160
                          '{ step_type : REG_WRITE, reg_addr : 32'h44450, value : 32'h80000480}, //phyinit_io_write: 0x4444f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44451, value : 32'h802}, //phyinit_io_write: 0x44450, 0x80000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44452, value : 32'h4000400}, //phyinit_io_write: 0x44451, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h44453, value : 32'h0}, //phyinit_io_write: 0x44452, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44454, value : 32'h80000080}, //phyinit_io_write: 0x44453, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44455, value : 32'h802}, //phyinit_io_write: 0x44454, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44456, value : 32'h4000400}, //phyinit_io_write: 0x44455, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h44457, value : 32'h0}, //phyinit_io_write: 0x44456, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44458, value : 32'he4000480}, //phyinit_io_write: 0x44457, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44459, value : 32'h801}, //phyinit_io_write: 0x44458, 0xe4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4445a, value : 32'h4000800}, //phyinit_io_write: 0x44459, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h4445b, value : 32'h0}, //phyinit_io_write: 0x4445a, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4445c, value : 32'he4000080}, //phyinit_io_write: 0x4445b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4445d, value : 32'h801}, //phyinit_io_write: 0x4445c, 0xe4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4445e, value : 32'ha8000080}, //phyinit_io_write: 0x4445d, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h4445f, value : 32'h1c04}, //phyinit_io_write: 0x4445e, 0xa8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44460, value : 32'hb8000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 12
                          '{ step_type : REG_WRITE, reg_addr : 32'h44461, value : 32'h801}, //phyinit_io_write: 0x44460, 0xb8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44462, value : 32'h4000800}, //phyinit_io_write: 0x44461, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44463, value : 32'h0}, //phyinit_io_write: 0x44462, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44464, value : 32'h1080}, //phyinit_io_write: 0x44463, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44465, value : 32'h33c2}, //phyinit_io_write: 0x44464, 0x1080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44466, value : 32'h50000480}, //phyinit_io_write: 0x44465, 0x33c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44467, value : 32'h1c01}, //phyinit_io_write: 0x44466, 0x50000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44468, value : 32'hb4000080}, //phyinit_io_write: 0x44467, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44469, value : 32'h2400}, //phyinit_io_write: 0x44468, 0xb4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4446a, value : 32'h88000481}, //phyinit_io_write: 0x44469, 0x2400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4446b, value : 32'hc00}, //phyinit_io_write: 0x4446a, 0x88000481
                          '{ step_type : REG_WRITE, reg_addr : 32'h4446c, value : 32'h24000480}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4446d, value : 32'h1c01}, //phyinit_io_write: 0x4446c, 0x24000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4446e, value : 32'h1e0}, //phyinit_io_write: 0x4446d, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h4446f, value : 32'h0}, //phyinit_io_write: 0x4446e, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44470, value : 32'h40000480}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 84
                          '{ step_type : REG_WRITE, reg_addr : 32'h44471, value : 32'h2c0c}, //phyinit_io_write: 0x44470, 0x40000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44472, value : 32'h2c000080}, //phyinit_io_write: 0x44471, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h44473, value : 32'h7c2}, //phyinit_io_write: 0x44472, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44474, value : 32'h8c000080}, //phyinit_io_write: 0x44473, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44475, value : 32'hfc2}, //phyinit_io_write: 0x44474, 0x8c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44476, value : 32'h200600}, //phyinit_io_write: 0x44475, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44477, value : 32'h20}, //phyinit_io_write: 0x44476, 0x200600
                          '{ step_type : REG_WRITE, reg_addr : 32'h44478, value : 32'h880c0080}, //phyinit_io_write: 0x44477, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h44479, value : 32'hc02}, //phyinit_io_write: 0x44478, 0x880c0080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4447a, value : 32'h880c00c0}, //phyinit_io_write: 0x44479, 0xc02
                          '{ step_type : REG_WRITE, reg_addr : 32'h4447b, value : 32'hc42}, //phyinit_io_write: 0x4447a, 0x880c00c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4447c, value : 32'h247ffc80}, //phyinit_io_write: 0x4447b, 0xc42
                          '{ step_type : REG_WRITE, reg_addr : 32'h4447d, value : 32'h7c2}, //phyinit_io_write: 0x4447c, 0x247ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h4447e, value : 32'h281ffc80}, //phyinit_io_write: 0x4447d, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4447f, value : 32'h7c2}, //phyinit_io_write: 0x4447e, 0x281ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44480, value : 32'h4000400}, //phyinit_io_write: 0x4447f, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44481, value : 32'h0}, //phyinit_io_write: 0x44480, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44482, value : 32'h98000480}, //phyinit_io_write: 0x44481, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44483, value : 32'hfc2}, //phyinit_io_write: 0x44482, 0x98000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44484, value : 32'h28000480}, //phyinit_io_write: 0x44483, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44485, value : 32'hfc0}, //phyinit_io_write: 0x44484, 0x28000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44486, value : 32'h4001000}, //phyinit_io_write: 0x44485, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44487, value : 32'h0}, //phyinit_io_write: 0x44486, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44488, value : 32'h80fffc80}, //phyinit_io_write: 0x44487, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44489, value : 32'hfc2}, //phyinit_io_write: 0x44488, 0x80fffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h4448a, value : 32'h4000400}, //phyinit_io_write: 0x44489, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4448b, value : 32'h0}, //phyinit_io_write: 0x4448a, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h4448c, value : 32'he0000480}, //phyinit_io_write: 0x4448b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4448d, value : 32'h803}, //phyinit_io_write: 0x4448c, 0xe0000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h4448e, value : 32'h4002000}, //phyinit_io_write: 0x4448d, 0x803
                          '{ step_type : REG_WRITE, reg_addr : 32'h4448f, value : 32'h0}, //phyinit_io_write: 0x4448e, 0x4002000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44490, value : 32'h28000080}, //phyinit_io_write: 0x4448f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44491, value : 32'hfc0}, //phyinit_io_write: 0x44490, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44492, value : 32'h50000080}, //phyinit_io_write: 0x44491, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44493, value : 32'h1c01}, //phyinit_io_write: 0x44492, 0x50000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44494, value : 32'h480}, //phyinit_io_write: 0x44493, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44495, value : 32'h1800}, //phyinit_io_write: 0x44494, 0x480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44496, value : 32'hc000080}, //phyinit_io_write: 0x44495, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44497, value : 32'h1800}, //phyinit_io_write: 0x44496, 0xc000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44498, value : 32'h5c000080}, //phyinit_io_write: 0x44497, 0x1800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44499, value : 32'h7c2}, //phyinit_io_write: 0x44498, 0x5c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4449a, value : 32'h4000080}, //phyinit_io_write: 0x44499, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4449b, value : 32'h2c00}, //phyinit_io_write: 0x4449a, 0x4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4449c, value : 32'h2000600}, //phyinit_io_write: 0x4449b, 0x2c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h4449d, value : 32'h200}, //phyinit_io_write: 0x4449c, 0x2000600
                          '{ step_type : REG_WRITE, reg_addr : 32'h4449e, value : 32'h2c0010c0}, //phyinit_io_write: 0x4449d, 0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h4449f, value : 32'h3bc1}, //phyinit_io_write: 0x4449e, 0x2c0010c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a0, value : 32'h2c001880}, //phyinit_io_write: 0x4449f, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a1, value : 32'h3bc1}, //phyinit_io_write: 0x444a0, 0x2c001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a2, value : 32'h18001880}, //phyinit_io_write: 0x444a1, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a3, value : 32'h3bc1}, //phyinit_io_write: 0x444a2, 0x18001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a4, value : 32'h1c001880}, //phyinit_io_write: 0x444a3, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a5, value : 32'h3bc1}, //phyinit_io_write: 0x444a4, 0x1c001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a6, value : 32'h20001880}, //phyinit_io_write: 0x444a5, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a7, value : 32'h3bc1}, //phyinit_io_write: 0x444a6, 0x20001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a8, value : 32'h24001880}, //phyinit_io_write: 0x444a7, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h444a9, value : 32'h3bc1}, //phyinit_io_write: 0x444a8, 0x24001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h444aa, value : 32'h28001880}, //phyinit_io_write: 0x444a9, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ab, value : 32'h3bc1}, //phyinit_io_write: 0x444aa, 0x28001880
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ac, value : 32'h20000880}, //phyinit_io_write: 0x444ab, 0x3bc1
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ad, value : 32'h2bcc}, //phyinit_io_write: 0x444ac, 0x20000880
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ae, value : 32'h40030a0}, //phyinit_io_write: 0x444ad, 0x2bcc
                          '{ step_type : REG_WRITE, reg_addr : 32'h444af, value : 32'h2c00}, //phyinit_io_write: 0x444ae, 0x40030a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b0, value : 32'h24000080}, //phyinit_io_write: 0x444af, 0x2c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b1, value : 32'h1c01}, //phyinit_io_write: 0x444b0, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b2, value : 32'hb4000480}, //phyinit_io_write: 0x444b1, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b3, value : 32'h2400}, //phyinit_io_write: 0x444b2, 0xb4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b4, value : 32'h40}, //phyinit_io_write: 0x444b3, 0x2400
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b5, value : 32'h4000}, //phyinit_io_write: 0x444b4, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b6, value : 32'h20}, //phyinit_io_write: 0x444b5, 0x4000
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b7, value : 32'h0}, //phyinit_io_write: 0x444b6, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b8, value : 32'h20}, //phyinit_io_write: 0x444b7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444b9, value : 32'h0}, //phyinit_io_write: 0x444b8, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ba, value : 32'h88000c80}, //phyinit_io_write: 0x444b9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444bb, value : 32'hc00}, //phyinit_io_write: 0x444ba, 0x88000c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h444bc, value : 32'h80000080}, //phyinit_io_write: 0x444bb, 0xc00
                          '{ step_type : REG_WRITE, reg_addr : 32'h444bd, value : 32'hfc0}, //phyinit_io_write: 0x444bc, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h444be, value : 32'h4000c00}, //phyinit_io_write: 0x444bd, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444bf, value : 32'h0}, //phyinit_io_write: 0x444be, 0x4000c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c0, value : 32'h88000480}, //phyinit_io_write: 0x444bf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c1, value : 32'h802}, //phyinit_io_write: 0x444c0, 0x88000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c2, value : 32'h1e0}, //phyinit_io_write: 0x444c1, 0x802
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c3, value : 32'h0}, //phyinit_io_write: 0x444c2, 0x1e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c4, value : 32'h1880}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c5, value : 32'h33c2}, //phyinit_io_write: 0x444c4, 0x1880
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c6, value : 32'h9c1}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 14
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c7, value : 32'h0}, //phyinit_io_write: 0x444c6, 0x9c1
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c8, value : 32'h9c000d11}, //phyinit_io_write: 0x444c7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444c9, value : 32'h1c01}, //phyinit_io_write: 0x444c8, 0x9c000d11
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ca, value : 32'h4001011}, //phyinit_io_write: 0x444c9, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h444cb, value : 32'h0}, //phyinit_io_write: 0x444ca, 0x4001011
                          '{ step_type : REG_WRITE, reg_addr : 32'h444cc, value : 32'h9c001111}, //phyinit_io_write: 0x444cb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444cd, value : 32'h1c03}, //phyinit_io_write: 0x444cc, 0x9c001111
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ce, value : 32'h4001011}, //phyinit_io_write: 0x444cd, 0x1c03
                          '{ step_type : REG_WRITE, reg_addr : 32'h444cf, value : 32'h0}, //phyinit_io_write: 0x444ce, 0x4001011
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d0, value : 32'h9c000091}, //phyinit_io_write: 0x444cf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d1, value : 32'h1c01}, //phyinit_io_write: 0x444d0, 0x9c000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d2, value : 32'h9c000091}, //phyinit_io_write: 0x444d1, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d3, value : 32'h1c03}, //phyinit_io_write: 0x444d2, 0x9c000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d4, value : 32'h9c921}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d5, value : 32'h0}, //phyinit_io_write: 0x444d4, 0x9c921
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d6, value : 32'hb8000480}, //phyinit_io_write: 0x444d5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d7, value : 32'h801}, //phyinit_io_write: 0x444d6, 0xb8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d8, value : 32'h4000800}, //phyinit_io_write: 0x444d7, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h444d9, value : 32'h0}, //phyinit_io_write: 0x444d8, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h444da, value : 32'h80068200}, //phyinit_io_write: 0x444d9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444db, value : 32'h400f}, //phyinit_io_write: 0x444da, 0x80068200
                          '{ step_type : REG_WRITE, reg_addr : 32'h444dc, value : 32'h9c140}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444dd, value : 32'h0}, //phyinit_io_write: 0x444dc, 0x9c140
                          '{ step_type : REG_WRITE, reg_addr : 32'h444de, value : 32'h8dc0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444df, value : 32'h0}, //phyinit_io_write: 0x444de, 0x8dc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e0, value : 32'h17dc0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e1, value : 32'h0}, //phyinit_io_write: 0x444e0, 0x17dc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e2, value : 32'h2a1c0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e3, value : 32'h0}, //phyinit_io_write: 0x444e2, 0x2a1c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e4, value : 32'h36dc0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e5, value : 32'h0}, //phyinit_io_write: 0x444e4, 0x36dc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e6, value : 32'h395c0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e7, value : 32'h0}, //phyinit_io_write: 0x444e6, 0x395c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e8, value : 32'h3adc0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444e9, value : 32'h0}, //phyinit_io_write: 0x444e8, 0x3adc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ea, value : 32'h5b9c0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 6
                          '{ step_type : REG_WRITE, reg_addr : 32'h444eb, value : 32'h0}, //phyinit_io_write: 0x444ea, 0x5b9c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ec, value : 32'h6001c080}, //phyinit_io_write: 0x444eb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ed, value : 32'h2425}, //phyinit_io_write: 0x444ec, 0x6001c080
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ee, value : 32'h80200}, //phyinit_io_write: 0x444ed, 0x2425
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ef, value : 32'h400e}, //phyinit_io_write: 0x444ee, 0x80200
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f0, value : 32'ha0940}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f1, value : 32'h0}, //phyinit_io_write: 0x444f0, 0xa0940
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f2, value : 32'h9ed31}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f3, value : 32'h0}, //phyinit_io_write: 0x444f2, 0x9ed31
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f4, value : 32'h6f9c0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f5, value : 32'h0}, //phyinit_io_write: 0x444f4, 0x6f9c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f6, value : 32'h80008600}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f7, value : 32'h0}, //phyinit_io_write: 0x444f6, 0x80008600
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f8, value : 32'ha0940}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444f9, value : 32'h0}, //phyinit_io_write: 0x444f8, 0xa0940
                          '{ step_type : REG_WRITE, reg_addr : 32'h444fa, value : 32'h739c2}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444fb, value : 32'h0}, //phyinit_io_write: 0x444fa, 0x739c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h444fc, value : 32'h80068200}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h444fd, value : 32'h400f}, //phyinit_io_write: 0x444fc, 0x80068200
                          '{ step_type : REG_WRITE, reg_addr : 32'h444fe, value : 32'hc40004c0}, //phyinit_io_write: 0x444fd, 0x400f
                          '{ step_type : REG_WRITE, reg_addr : 32'h444ff, value : 32'h7c0}, //phyinit_io_write: 0x444fe, 0xc40004c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44500, value : 32'h4001000}, //phyinit_io_write: 0x444ff, 0x7c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44501, value : 32'h0}, //phyinit_io_write: 0x44500, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44502, value : 32'hc40000c0}, //phyinit_io_write: 0x44501, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44503, value : 32'h7c0}, //phyinit_io_write: 0x44502, 0xc40000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44504, value : 32'h40006611}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44505, value : 32'h0}, //phyinit_io_write: 0x44504, 0x40006611
                          '{ step_type : REG_WRITE, reg_addr : 32'h44506, value : 32'ha5151}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h44507, value : 32'h0}, //phyinit_io_write: 0x44506, 0xa5151
                          '{ step_type : REG_WRITE, reg_addr : 32'h44508, value : 32'h80068211}, //phyinit_io_write: 0x44507, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44509, value : 32'h400f}, //phyinit_io_write: 0x44508, 0x80068211
                          '{ step_type : REG_WRITE, reg_addr : 32'h4450a, value : 32'ha5151}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4450b, value : 32'h0}, //phyinit_io_write: 0x4450a, 0xa5151
                          '{ step_type : REG_WRITE, reg_addr : 32'h4450c, value : 32'h80211}, //phyinit_io_write: 0x4450b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4450d, value : 32'h400e}, //phyinit_io_write: 0x4450c, 0x80211
                          '{ step_type : REG_WRITE, reg_addr : 32'h4450e, value : 32'ha2951}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4450f, value : 32'h0}, //phyinit_io_write: 0x4450e, 0xa2951
                          '{ step_type : REG_WRITE, reg_addr : 32'h44510, value : 32'h80008611}, //phyinit_io_write: 0x4450f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44511, value : 32'h0}, //phyinit_io_write: 0x44510, 0x80008611
                          '{ step_type : REG_WRITE, reg_addr : 32'h44512, value : 32'ha3571}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44513, value : 32'h0}, //phyinit_io_write: 0x44512, 0xa3571
                          '{ step_type : REG_WRITE, reg_addr : 32'h44514, value : 32'h1031}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 6
                          '{ step_type : REG_WRITE, reg_addr : 32'h44515, value : 32'h0}, //phyinit_io_write: 0x44514, 0x1031
                          '{ step_type : REG_WRITE, reg_addr : 32'h44516, value : 32'h1031}, //phyinit_io_write: 0x44515, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44517, value : 32'h0}, //phyinit_io_write: 0x44516, 0x1031
                          '{ step_type : REG_WRITE, reg_addr : 32'h44518, value : 32'h2c31}, //phyinit_io_write: 0x44517, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44519, value : 32'h0}, //phyinit_io_write: 0x44518, 0x2c31
                          '{ step_type : REG_WRITE, reg_addr : 32'h4451a, value : 32'ha8000091}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 14
                          '{ step_type : REG_WRITE, reg_addr : 32'h4451b, value : 32'h1c06}, //phyinit_io_write: 0x4451a, 0xa8000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h4451c, value : 32'h80016891}, //phyinit_io_write: 0x4451b, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h4451d, value : 32'h1c04}, //phyinit_io_write: 0x4451c, 0x80016891
                          '{ step_type : REG_WRITE, reg_addr : 32'h4451e, value : 32'h4000400}, //phyinit_io_write: 0x4451d, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4451f, value : 32'h0}, //phyinit_io_write: 0x4451e, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44520, value : 32'h80016c91}, //phyinit_io_write: 0x4451f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44521, value : 32'h1c04}, //phyinit_io_write: 0x44520, 0x80016c91
                          '{ step_type : REG_WRITE, reg_addr : 32'h44522, value : 32'h4000800}, //phyinit_io_write: 0x44521, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44523, value : 32'h0}, //phyinit_io_write: 0x44522, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44524, value : 32'h851}, //phyinit_io_write: 0x44523, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44525, value : 32'h6000}, //phyinit_io_write: 0x44524, 0x851
                          '{ step_type : REG_WRITE, reg_addr : 32'h44526, value : 32'h80000091}, //phyinit_io_write: 0x44525, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44527, value : 32'h1c04}, //phyinit_io_write: 0x44526, 0x80000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h44528, value : 32'h24000091}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44529, value : 32'h1e420}, //phyinit_io_write: 0x44528, 0x24000091
                          '{ step_type : REG_WRITE, reg_addr : 32'h4452a, value : 32'h899c0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4452b, value : 32'h0}, //phyinit_io_write: 0x4452a, 0x899c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4452c, value : 32'h0}, //phyinit_io_write: 0x4452b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4452d, value : 32'h0}, //phyinit_io_write: 0x4452c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4452e, value : 32'h8e1c0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 6
                          '{ step_type : REG_WRITE, reg_addr : 32'h4452f, value : 32'h0}, //phyinit_io_write: 0x4452e, 0x8e1c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44530, value : 32'h24000480}, //phyinit_io_write: 0x4452f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44531, value : 32'h1c01}, //phyinit_io_write: 0x44530, 0x24000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44532, value : 32'h400}, //phyinit_io_write: 0x44531, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44533, value : 32'h0}, //phyinit_io_write: 0x44532, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44534, value : 32'h50000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 22
                          '{ step_type : REG_WRITE, reg_addr : 32'h44535, value : 32'h1c01}, //phyinit_io_write: 0x44534, 0x50000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44536, value : 32'h9c000d00}, //phyinit_io_write: 0x44535, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44537, value : 32'h1c01}, //phyinit_io_write: 0x44536, 0x9c000d00
                          '{ step_type : REG_WRITE, reg_addr : 32'h44538, value : 32'h4001000}, //phyinit_io_write: 0x44537, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44539, value : 32'h0}, //phyinit_io_write: 0x44538, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4453a, value : 32'h9c001100}, //phyinit_io_write: 0x44539, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4453b, value : 32'h1c03}, //phyinit_io_write: 0x4453a, 0x9c001100
                          '{ step_type : REG_WRITE, reg_addr : 32'h4453c, value : 32'h4001000}, //phyinit_io_write: 0x4453b, 0x1c03
                          '{ step_type : REG_WRITE, reg_addr : 32'h4453d, value : 32'h0}, //phyinit_io_write: 0x4453c, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4453e, value : 32'h9c000080}, //phyinit_io_write: 0x4453d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4453f, value : 32'h1c01}, //phyinit_io_write: 0x4453e, 0x9c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44540, value : 32'h9c000080}, //phyinit_io_write: 0x4453f, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44541, value : 32'h1c03}, //phyinit_io_write: 0x44540, 0x9c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44542, value : 32'h1880}, //phyinit_io_write: 0x44541, 0x1c03
                          '{ step_type : REG_WRITE, reg_addr : 32'h44543, value : 32'h33c2}, //phyinit_io_write: 0x44542, 0x1880
                          '{ step_type : REG_WRITE, reg_addr : 32'h44544, value : 32'hb8000480}, //phyinit_io_write: 0x44543, 0x33c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44545, value : 32'h801}, //phyinit_io_write: 0x44544, 0xb8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44546, value : 32'h4000c00}, //phyinit_io_write: 0x44545, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h44547, value : 32'h0}, //phyinit_io_write: 0x44546, 0x4000c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h44548, value : 32'h24000491}, //phyinit_io_write: 0x44547, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44549, value : 32'h1e420}, //phyinit_io_write: 0x44548, 0x24000491
                          '{ step_type : REG_WRITE, reg_addr : 32'h4454a, value : 32'ha8000080}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 10
                          '{ step_type : REG_WRITE, reg_addr : 32'h4454b, value : 32'h1c06}, //phyinit_io_write: 0x4454a, 0xa8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4454c, value : 32'h80012880}, //phyinit_io_write: 0x4454b, 0x1c06
                          '{ step_type : REG_WRITE, reg_addr : 32'h4454d, value : 32'h1c04}, //phyinit_io_write: 0x4454c, 0x80012880
                          '{ step_type : REG_WRITE, reg_addr : 32'h4454e, value : 32'h4000400}, //phyinit_io_write: 0x4454d, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h4454f, value : 32'h0}, //phyinit_io_write: 0x4454e, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44550, value : 32'h80012c80}, //phyinit_io_write: 0x4454f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44551, value : 32'h1c04}, //phyinit_io_write: 0x44550, 0x80012c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44552, value : 32'h4000800}, //phyinit_io_write: 0x44551, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44553, value : 32'h0}, //phyinit_io_write: 0x44552, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44554, value : 32'h840}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 70
                          '{ step_type : REG_WRITE, reg_addr : 32'h44555, value : 32'h6000}, //phyinit_io_write: 0x44554, 0x840
                          '{ step_type : REG_WRITE, reg_addr : 32'h44556, value : 32'h80000080}, //phyinit_io_write: 0x44555, 0x6000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44557, value : 32'h1c04}, //phyinit_io_write: 0x44556, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44558, value : 32'h2c000080}, //phyinit_io_write: 0x44557, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h44559, value : 32'h7c2}, //phyinit_io_write: 0x44558, 0x2c000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4455a, value : 32'h8c200080}, //phyinit_io_write: 0x44559, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4455b, value : 32'hfc2}, //phyinit_io_write: 0x4455a, 0x8c200080
                          '{ step_type : REG_WRITE, reg_addr : 32'h4455c, value : 32'h200600}, //phyinit_io_write: 0x4455b, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4455d, value : 32'h20}, //phyinit_io_write: 0x4455c, 0x200600
                          '{ step_type : REG_WRITE, reg_addr : 32'h4455e, value : 32'h883c0080}, //phyinit_io_write: 0x4455d, 0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h4455f, value : 32'hc02}, //phyinit_io_write: 0x4455e, 0x883c0080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44560, value : 32'h883c00c0}, //phyinit_io_write: 0x4455f, 0xc02
                          '{ step_type : REG_WRITE, reg_addr : 32'h44561, value : 32'hc42}, //phyinit_io_write: 0x44560, 0x883c00c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44562, value : 32'h98000480}, //phyinit_io_write: 0x44561, 0xc42
                          '{ step_type : REG_WRITE, reg_addr : 32'h44563, value : 32'hfc2}, //phyinit_io_write: 0x44562, 0x98000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44564, value : 32'h28000480}, //phyinit_io_write: 0x44563, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44565, value : 32'hfc0}, //phyinit_io_write: 0x44564, 0x28000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44566, value : 32'h4001000}, //phyinit_io_write: 0x44565, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44567, value : 32'h0}, //phyinit_io_write: 0x44566, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44568, value : 32'h80fffc80}, //phyinit_io_write: 0x44567, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44569, value : 32'hfc2}, //phyinit_io_write: 0x44568, 0x80fffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h4456a, value : 32'h247ffc80}, //phyinit_io_write: 0x44569, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4456b, value : 32'h7c2}, //phyinit_io_write: 0x4456a, 0x247ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h4456c, value : 32'h281ffc80}, //phyinit_io_write: 0x4456b, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4456d, value : 32'h7c2}, //phyinit_io_write: 0x4456c, 0x281ffc80
                          '{ step_type : REG_WRITE, reg_addr : 32'h4456e, value : 32'h4000400}, //phyinit_io_write: 0x4456d, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4456f, value : 32'h0}, //phyinit_io_write: 0x4456e, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h44570, value : 32'he0000480}, //phyinit_io_write: 0x4456f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44571, value : 32'h803}, //phyinit_io_write: 0x44570, 0xe0000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h44572, value : 32'h28000080}, //phyinit_io_write: 0x44571, 0x803
                          '{ step_type : REG_WRITE, reg_addr : 32'h44573, value : 32'hfc0}, //phyinit_io_write: 0x44572, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44574, value : 32'h800600}, //phyinit_io_write: 0x44573, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44575, value : 32'h80}, //phyinit_io_write: 0x44574, 0x800600
                          '{ step_type : REG_WRITE, reg_addr : 32'h44576, value : 32'h40000c0}, //phyinit_io_write: 0x44575, 0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h44577, value : 32'h2424}, //phyinit_io_write: 0x44576, 0x40000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44578, value : 32'h40080e0}, //phyinit_io_write: 0x44577, 0x2424
                          '{ step_type : REG_WRITE, reg_addr : 32'h44579, value : 32'h2424}, //phyinit_io_write: 0x44578, 0x40080e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4457a, value : 32'h400004e2}, //phyinit_io_write: 0x44579, 0x2424
                          '{ step_type : REG_WRITE, reg_addr : 32'h4457b, value : 32'h2c0c}, //phyinit_io_write: 0x4457a, 0x400004e2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4457c, value : 32'h4000800}, //phyinit_io_write: 0x4457b, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h4457d, value : 32'h0}, //phyinit_io_write: 0x4457c, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4457e, value : 32'h400000e2}, //phyinit_io_write: 0x4457d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4457f, value : 32'h2c0c}, //phyinit_io_write: 0x4457e, 0x400000e2
                          '{ step_type : REG_WRITE, reg_addr : 32'h44580, value : 32'h4000800}, //phyinit_io_write: 0x4457f, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h44581, value : 32'h0}, //phyinit_io_write: 0x44580, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44582, value : 32'h800004e0}, //phyinit_io_write: 0x44581, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44583, value : 32'h2c0c}, //phyinit_io_write: 0x44582, 0x800004e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44584, value : 32'h800000e0}, //phyinit_io_write: 0x44583, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h44585, value : 32'h2c0c}, //phyinit_io_write: 0x44584, 0x800000e0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44586, value : 32'h605}, //phyinit_io_write: 0x44585, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h44587, value : 32'h2000}, //phyinit_io_write: 0x44586, 0x605
                          '{ step_type : REG_WRITE, reg_addr : 32'h44588, value : 32'h400004c2}, //phyinit_io_write: 0x44587, 0x2000
                          '{ step_type : REG_WRITE, reg_addr : 32'h44589, value : 32'h2c0c}, //phyinit_io_write: 0x44588, 0x400004c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4458a, value : 32'h4000800}, //phyinit_io_write: 0x44589, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h4458b, value : 32'h0}, //phyinit_io_write: 0x4458a, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h4458c, value : 32'h400000c2}, //phyinit_io_write: 0x4458b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4458d, value : 32'h2c0c}, //phyinit_io_write: 0x4458c, 0x400000c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4458e, value : 32'h4000800}, //phyinit_io_write: 0x4458d, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h4458f, value : 32'h0}, //phyinit_io_write: 0x4458e, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h44590, value : 32'h800004c0}, //phyinit_io_write: 0x4458f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44591, value : 32'h2c0c}, //phyinit_io_write: 0x44590, 0x800004c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44592, value : 32'h800000c0}, //phyinit_io_write: 0x44591, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h44593, value : 32'h2c0c}, //phyinit_io_write: 0x44592, 0x800000c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44594, value : 32'h4000c00}, //phyinit_io_write: 0x44593, 0x2c0c
                          '{ step_type : REG_WRITE, reg_addr : 32'h44595, value : 32'h0}, //phyinit_io_write: 0x44594, 0x4000c00
                          '{ step_type : REG_WRITE, reg_addr : 32'h44596, value : 32'h24000080}, //phyinit_io_write: 0x44595, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h44597, value : 32'h1c01}, //phyinit_io_write: 0x44596, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h44598, value : 32'h10000200}, //phyinit_io_write: 0x44597, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h44599, value : 32'h5000}, //phyinit_io_write: 0x44598, 0x10000200
                          '{ step_type : REG_WRITE, reg_addr : 32'h4459a, value : 32'hb3d40}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4459b, value : 32'h0}, //phyinit_io_write: 0x4459a, 0xb3d40
                          '{ step_type : REG_WRITE, reg_addr : 32'h4459c, value : 32'h40}, //phyinit_io_write: 0x4459b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4459d, value : 32'h4000}, //phyinit_io_write: 0x4459c, 0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h4459e, value : 32'h28000480}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 36
                          '{ step_type : REG_WRITE, reg_addr : 32'h4459f, value : 32'hfc0}, //phyinit_io_write: 0x4459e, 0x28000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a0, value : 32'h4001000}, //phyinit_io_write: 0x4459f, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a1, value : 32'h0}, //phyinit_io_write: 0x445a0, 0x4001000
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a2, value : 32'he0000080}, //phyinit_io_write: 0x445a1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a3, value : 32'h803}, //phyinit_io_write: 0x445a2, 0xe0000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a4, value : 32'h4000800}, //phyinit_io_write: 0x445a3, 0x803
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a5, value : 32'h0}, //phyinit_io_write: 0x445a4, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a6, value : 32'h28000080}, //phyinit_io_write: 0x445a5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a7, value : 32'hfc0}, //phyinit_io_write: 0x445a6, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a8, value : 32'h80000080}, //phyinit_io_write: 0x445a7, 0xfc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445a9, value : 32'hfc2}, //phyinit_io_write: 0x445a8, 0x80000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h445aa, value : 32'h98000080}, //phyinit_io_write: 0x445a9, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h445ab, value : 32'hfc2}, //phyinit_io_write: 0x445aa, 0x98000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h445ac, value : 32'h24000080}, //phyinit_io_write: 0x445ab, 0xfc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h445ad, value : 32'h7c2}, //phyinit_io_write: 0x445ac, 0x24000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h445ae, value : 32'h28000080}, //phyinit_io_write: 0x445ad, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h445af, value : 32'h7c2}, //phyinit_io_write: 0x445ae, 0x28000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b0, value : 32'he4000480}, //phyinit_io_write: 0x445af, 0x7c2
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b1, value : 32'h801}, //phyinit_io_write: 0x445b0, 0xe4000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b2, value : 32'h4000800}, //phyinit_io_write: 0x445b1, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b3, value : 32'h0}, //phyinit_io_write: 0x445b2, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b4, value : 32'he4000080}, //phyinit_io_write: 0x445b3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b5, value : 32'h801}, //phyinit_io_write: 0x445b4, 0xe4000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b6, value : 32'h4000800}, //phyinit_io_write: 0x445b5, 0x801
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b7, value : 32'h0}, //phyinit_io_write: 0x445b6, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b8, value : 32'ha8000480}, //phyinit_io_write: 0x445b7, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445b9, value : 32'h1c04}, //phyinit_io_write: 0x445b8, 0xa8000480
                          '{ step_type : REG_WRITE, reg_addr : 32'h445ba, value : 32'h1020}, //phyinit_io_write: 0x445b9, 0x1c04
                          '{ step_type : REG_WRITE, reg_addr : 32'h445bb, value : 32'h0}, //phyinit_io_write: 0x445ba, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h445bc, value : 32'h1020}, //phyinit_io_write: 0x445bb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445bd, value : 32'h0}, //phyinit_io_write: 0x445bc, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h445be, value : 32'h1020}, //phyinit_io_write: 0x445bd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445bf, value : 32'h0}, //phyinit_io_write: 0x445be, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c0, value : 32'h1020}, //phyinit_io_write: 0x445bf, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c1, value : 32'h0}, //phyinit_io_write: 0x445c0, 0x1020
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c2, value : 32'he8030c80}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 8
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c3, value : 32'h1c01}, //phyinit_io_write: 0x445c2, 0xe8030c80
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c4, value : 32'h4000800}, //phyinit_io_write: 0x445c3, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c5, value : 32'h0}, //phyinit_io_write: 0x445c4, 0x4000800
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c6, value : 32'he8000080}, //phyinit_io_write: 0x445c5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c7, value : 32'h1c01}, //phyinit_io_write: 0x445c6, 0xe8000080
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c8, value : 32'h4000400}, //phyinit_io_write: 0x445c7, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h445c9, value : 32'h0}, //phyinit_io_write: 0x445c8, 0x4000400
                          '{ step_type : REG_WRITE, reg_addr : 32'h445ca, value : 32'h9c000ca0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h445cb, value : 32'h1c01}, //phyinit_io_write: 0x445ca, 0x9c000ca0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445cc, value : 32'h9c0010a0}, //phyinit_io_write: 0x445cb, 0x1c01
                          '{ step_type : REG_WRITE, reg_addr : 32'h445cd, value : 32'h1c03}, //phyinit_io_write: 0x445cc, 0x9c0010a0
                          '{ step_type : REG_WRITE, reg_addr : 32'h445ce, value : 32'h9ed20}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h445cf, value : 32'h0}, //phyinit_io_write: 0x445ce, 0x9ed20
                          '{ step_type : REG_WRITE, reg_addr : 32'hd00e7, value : 32'h600}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 1
                          '{ step_type : REG_WRITE, reg_addr : 32'h7018a, value : 32'h0}, //[dwc_ddrphy_phyinit_LoadPIECodeSections] Writing code section size = 1
                          '{ step_type : REG_WRITE, reg_addr : 32'h70324, value : 32'h1}, //// The number of StartAddr is 65.
                          '{ step_type : REG_WRITE, reg_addr : 32'h70325, value : 32'h19}, //phyinit_io_write: 0x70324, 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h70326, value : 32'h2e}, //phyinit_io_write: 0x70325, 0x19
                          '{ step_type : REG_WRITE, reg_addr : 32'h70327, value : 32'h43}, //phyinit_io_write: 0x70326, 0x2e
                          '{ step_type : REG_WRITE, reg_addr : 32'h70328, value : 32'h5b}, //phyinit_io_write: 0x70327, 0x43
                          '{ step_type : REG_WRITE, reg_addr : 32'h70329, value : 32'h70}, //phyinit_io_write: 0x70328, 0x5b
                          '{ step_type : REG_WRITE, reg_addr : 32'h7032a, value : 32'h85}, //phyinit_io_write: 0x70329, 0x70
                          '{ step_type : REG_WRITE, reg_addr : 32'h7032b, value : 32'h9d}, //phyinit_io_write: 0x7032a, 0x85
                          '{ step_type : REG_WRITE, reg_addr : 32'h7032c, value : 32'hb2}, //phyinit_io_write: 0x7032b, 0x9d
                          '{ step_type : REG_WRITE, reg_addr : 32'h7032d, value : 32'hc7}, //phyinit_io_write: 0x7032c, 0xb2
                          '{ step_type : REG_WRITE, reg_addr : 32'h7032e, value : 32'hdf}, //phyinit_io_write: 0x7032d, 0xc7
                          '{ step_type : REG_WRITE, reg_addr : 32'h7032f, value : 32'hf4}, //phyinit_io_write: 0x7032e, 0xdf
                          '{ step_type : REG_WRITE, reg_addr : 32'h70330, value : 32'h109}, //phyinit_io_write: 0x7032f, 0xf4
                          '{ step_type : REG_WRITE, reg_addr : 32'h70331, value : 32'h113}, //phyinit_io_write: 0x70330, 0x109
                          '{ step_type : REG_WRITE, reg_addr : 32'h70332, value : 32'h115}, //phyinit_io_write: 0x70331, 0x113
                          '{ step_type : REG_WRITE, reg_addr : 32'h70333, value : 32'h119}, //phyinit_io_write: 0x70332, 0x115
                          '{ step_type : REG_WRITE, reg_addr : 32'h70334, value : 32'h11b}, //phyinit_io_write: 0x70333, 0x119
                          '{ step_type : REG_WRITE, reg_addr : 32'h70335, value : 32'h11f}, //phyinit_io_write: 0x70334, 0x11b
                          '{ step_type : REG_WRITE, reg_addr : 32'h70336, value : 32'h121}, //phyinit_io_write: 0x70335, 0x11f
                          '{ step_type : REG_WRITE, reg_addr : 32'h70337, value : 32'h122}, //phyinit_io_write: 0x70336, 0x121
                          '{ step_type : REG_WRITE, reg_addr : 32'h70339, value : 32'h123}, //phyinit_io_write: 0x70337, 0x122
                          '{ step_type : REG_WRITE, reg_addr : 32'h7033a, value : 32'h125}, //phyinit_io_write: 0x70339, 0x123
                          '{ step_type : REG_WRITE, reg_addr : 32'h7033c, value : 32'h126}, //phyinit_io_write: 0x7033a, 0x125
                          '{ step_type : REG_WRITE, reg_addr : 32'h7033d, value : 32'h13f}, //phyinit_io_write: 0x7033c, 0x126
                          '{ step_type : REG_WRITE, reg_addr : 32'h7033e, value : 32'h149}, //phyinit_io_write: 0x7033d, 0x13f
                          '{ step_type : REG_WRITE, reg_addr : 32'h7033f, value : 32'h161}, //phyinit_io_write: 0x7033e, 0x149
                          '{ step_type : REG_WRITE, reg_addr : 32'h70350, value : 32'h171}, //phyinit_io_write: 0x7033f, 0x161
                          '{ step_type : REG_WRITE, reg_addr : 32'h70351, value : 32'h189}, //phyinit_io_write: 0x70350, 0x171
                          '{ step_type : REG_WRITE, reg_addr : 32'h70352, value : 32'h192}, //phyinit_io_write: 0x70351, 0x189
                          '{ step_type : REG_WRITE, reg_addr : 32'h70353, value : 32'h1a4}, //phyinit_io_write: 0x70352, 0x192
                          '{ step_type : REG_WRITE, reg_addr : 32'h7038b, value : 32'h18}, //phyinit_io_write: 0x70353, 0x1a4
                          '{ step_type : REG_WRITE, reg_addr : 32'h7038c, value : 32'h2d}, //phyinit_io_write: 0x7038b, 0x18
                          '{ step_type : REG_WRITE, reg_addr : 32'h7038d, value : 32'h42}, //phyinit_io_write: 0x7038c, 0x2d
                          '{ step_type : REG_WRITE, reg_addr : 32'h7038e, value : 32'h5a}, //phyinit_io_write: 0x7038d, 0x42
                          '{ step_type : REG_WRITE, reg_addr : 32'h7038f, value : 32'h6f}, //phyinit_io_write: 0x7038e, 0x5a
                          '{ step_type : REG_WRITE, reg_addr : 32'h70390, value : 32'h84}, //phyinit_io_write: 0x7038f, 0x6f
                          '{ step_type : REG_WRITE, reg_addr : 32'h70391, value : 32'h9c}, //phyinit_io_write: 0x70390, 0x84
                          '{ step_type : REG_WRITE, reg_addr : 32'h70392, value : 32'hb1}, //phyinit_io_write: 0x70391, 0x9c
                          '{ step_type : REG_WRITE, reg_addr : 32'h70393, value : 32'hc6}, //phyinit_io_write: 0x70392, 0xb1
                          '{ step_type : REG_WRITE, reg_addr : 32'h70394, value : 32'hde}, //phyinit_io_write: 0x70393, 0xc6
                          '{ step_type : REG_WRITE, reg_addr : 32'h70395, value : 32'hf3}, //phyinit_io_write: 0x70394, 0xde
                          '{ step_type : REG_WRITE, reg_addr : 32'h70396, value : 32'h108}, //phyinit_io_write: 0x70395, 0xf3
                          '{ step_type : REG_WRITE, reg_addr : 32'h70397, value : 32'h112}, //phyinit_io_write: 0x70396, 0x108
                          '{ step_type : REG_WRITE, reg_addr : 32'h70398, value : 32'h114}, //phyinit_io_write: 0x70397, 0x112
                          '{ step_type : REG_WRITE, reg_addr : 32'h70399, value : 32'h118}, //phyinit_io_write: 0x70398, 0x114
                          '{ step_type : REG_WRITE, reg_addr : 32'h7039a, value : 32'h11a}, //phyinit_io_write: 0x70399, 0x118
                          '{ step_type : REG_WRITE, reg_addr : 32'h7039b, value : 32'h11e}, //phyinit_io_write: 0x7039a, 0x11a
                          '{ step_type : REG_WRITE, reg_addr : 32'h7039c, value : 32'h120}, //phyinit_io_write: 0x7039b, 0x11e
                          '{ step_type : REG_WRITE, reg_addr : 32'h7039d, value : 32'h121}, //phyinit_io_write: 0x7039c, 0x120
                          '{ step_type : REG_WRITE, reg_addr : 32'h7039e, value : 32'h122}, //phyinit_io_write: 0x7039d, 0x121
                          '{ step_type : REG_WRITE, reg_addr : 32'h703a0, value : 32'h124}, //phyinit_io_write: 0x7039e, 0x122
                          '{ step_type : REG_WRITE, reg_addr : 32'h703a1, value : 32'h125}, //phyinit_io_write: 0x703a0, 0x124
                          '{ step_type : REG_WRITE, reg_addr : 32'h703a3, value : 32'h13e}, //phyinit_io_write: 0x703a1, 0x125
                          '{ step_type : REG_WRITE, reg_addr : 32'h703a4, value : 32'h148}, //phyinit_io_write: 0x703a3, 0x13e
                          '{ step_type : REG_WRITE, reg_addr : 32'h703a5, value : 32'h160}, //phyinit_io_write: 0x703a4, 0x148
                          '{ step_type : REG_WRITE, reg_addr : 32'h703a6, value : 32'h170}, //phyinit_io_write: 0x703a5, 0x160
                          '{ step_type : REG_WRITE, reg_addr : 32'h703b7, value : 32'h188}, //phyinit_io_write: 0x703a6, 0x170
                          '{ step_type : REG_WRITE, reg_addr : 32'h703b8, value : 32'h191}, //phyinit_io_write: 0x703b7, 0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h703b9, value : 32'h1a3}, //phyinit_io_write: 0x703b8, 0x191
                          '{ step_type : REG_WRITE, reg_addr : 32'h703ba, value : 32'h1b4}, //phyinit_io_write: 0x703b9, 0x1a3
                          '{ step_type : REG_WRITE, reg_addr : 32'h70200, value : 32'h40e}, //phyinit_io_write: 0x703ba, 0x1b4
                          '{ step_type : REG_WRITE, reg_addr : 32'h70202, value : 32'h44f}, //phyinit_io_write: 0x70200, 0x40e
                          '{ step_type : REG_WRITE, reg_addr : 32'h70204, value : 32'hc0}, //phyinit_io_write: 0x70202, 0x44f
                          '{ step_type : REG_WRITE, reg_addr : 32'h70205, value : 32'h246}, //phyinit_io_write: 0x70204, 0xc0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70206, value : 32'h101}, //phyinit_io_write: 0x70205, 0x246
                          '{ step_type : REG_WRITE, reg_addr : 32'h70207, value : 32'h287}, //phyinit_io_write: 0x70206, 0x101
                          '{ step_type : REG_WRITE, reg_addr : 32'h70208, value : 32'h142}, //phyinit_io_write: 0x70207, 0x287
                          '{ step_type : REG_WRITE, reg_addr : 32'h70209, value : 32'h2c8}, //phyinit_io_write: 0x70208, 0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h7020a, value : 32'h12}, //phyinit_io_write: 0x70209, 0x2c8
                          '{ step_type : REG_WRITE, reg_addr : 32'h7020b, value : 32'h34c}, //phyinit_io_write: 0x7020a, 0x12
                          '{ step_type : REG_WRITE, reg_addr : 32'h7020c, value : 32'h15}, //phyinit_io_write: 0x7020b, 0x34c
                          '{ step_type : REG_WRITE, reg_addr : 32'h7020e, value : 32'h16}, //phyinit_io_write: 0x7020c, 0x15
                          '{ step_type : REG_WRITE, reg_addr : 32'h70212, value : 32'h2c}, //phyinit_io_write: 0x7020e, 0x16
                          '{ step_type : REG_WRITE, reg_addr : 32'h70213, value : 32'h18}, //phyinit_io_write: 0x70212, 0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h70214, value : 32'h2d}, //phyinit_io_write: 0x70213, 0x18
                          '{ step_type : REG_WRITE, reg_addr : 32'h70215, value : 32'h19}, //phyinit_io_write: 0x70214, 0x2d
                          '{ step_type : REG_WRITE, reg_addr : 32'h70216, value : 32'h2e}, //phyinit_io_write: 0x70215, 0x19
                          '{ step_type : REG_WRITE, reg_addr : 32'h70217, value : 32'h1a}, //phyinit_io_write: 0x70216, 0x2e
                          '{ step_type : REG_WRITE, reg_addr : 32'h70218, value : 32'h2f}, //phyinit_io_write: 0x70217, 0x1a
                          '{ step_type : REG_WRITE, reg_addr : 32'h70219, value : 32'h1b}, //phyinit_io_write: 0x70218, 0x2f
                          '{ step_type : REG_WRITE, reg_addr : 32'h7021a, value : 32'h13}, //phyinit_io_write: 0x70219, 0x1b
                          '{ step_type : REG_WRITE, reg_addr : 32'h9001c, value : 32'h262}, //phyinit_io_write: 0x7021a, 0x13
                          '{ step_type : REG_WRITE, reg_addr : 32'h9001d, value : 32'h262}, //phyinit_io_write: 0x9001c, 0x262
                          '{ step_type : REG_WRITE, reg_addr : 32'h9001e, value : 32'h262}, //phyinit_io_write: 0x9001d, 0x262
                          '{ step_type : REG_WRITE, reg_addr : 32'h9001f, value : 32'h262}, //phyinit_io_write: 0x9001e, 0x262
                          '{ step_type : REG_WRITE, reg_addr : 32'h90020, value : 32'h29a}, //phyinit_io_write: 0x9001f, 0x262
                          '{ step_type : REG_WRITE, reg_addr : 32'h90021, value : 32'h262}, //phyinit_io_write: 0x90020, 0x29a
                          '{ step_type : REG_WRITE, reg_addr : 32'h90022, value : 32'h0}, //phyinit_io_write: 0x90021, 0x262
                          '{ step_type : REG_WRITE, reg_addr : 32'h90023, value : 32'h0}, //phyinit_io_write: 0x90022, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90024, value : 32'h0}, //phyinit_io_write: 0x90023, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90025, value : 32'h0}, //phyinit_io_write: 0x90024, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90026, value : 32'h0}, //phyinit_io_write: 0x90025, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90027, value : 32'h0}, //phyinit_io_write: 0x90026, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h9002b, value : 32'h297}, //phyinit_io_write: 0x90027, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70145, value : 32'h2}, //[loadAcsmMRW] Pstate=0, Programming ACSMRptCntOverride to 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41004, value : 32'hc9d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=19 OP=0x0 CS=0xf at row addr=0x2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41005, value : 32'h0}, //phyinit_io_write: 0x41004, 0xc9d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41006, value : 32'hc008}, //phyinit_io_write: 0x41005, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41007, value : 32'h0}, //phyinit_io_write: 0x41006, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41008, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41009, value : 32'h4b000000}, //phyinit_io_write: 0x41008, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4100a, value : 32'h0}, //phyinit_io_write: 0x41009, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4100b, value : 32'h0}, //phyinit_io_write: 0x4100a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4100c, value : 32'hc958}, //[dwc_ddrphy_mr_inst] Storing MRW MA=18 OP=0x0 CS=0xf at row addr=0x6
                          '{ step_type : REG_WRITE, reg_addr : 32'h4100d, value : 32'h0}, //phyinit_io_write: 0x4100c, 0xc958
                          '{ step_type : REG_WRITE, reg_addr : 32'h4100e, value : 32'hc008}, //phyinit_io_write: 0x4100d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4100f, value : 32'h0}, //phyinit_io_write: 0x4100e, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41010, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41011, value : 32'h4b000000}, //phyinit_io_write: 0x41010, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41012, value : 32'h0}, //phyinit_io_write: 0x41011, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41013, value : 32'h0}, //phyinit_io_write: 0x41012, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41014, value : 32'hc0d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=1 OP=0xb0 CS=0xf at row addr=0xa
                          '{ step_type : REG_WRITE, reg_addr : 32'h41015, value : 32'h0}, //phyinit_io_write: 0x41014, 0xc0d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41016, value : 32'hd848}, //phyinit_io_write: 0x41015, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41017, value : 32'h0}, //phyinit_io_write: 0x41016, 0xd848
                          '{ step_type : REG_WRITE, reg_addr : 32'h41018, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41019, value : 32'h4b000000}, //phyinit_io_write: 0x41018, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4101a, value : 32'h0}, //phyinit_io_write: 0x41019, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4101b, value : 32'h0}, //phyinit_io_write: 0x4101a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4101c, value : 32'hc158}, //[dwc_ddrphy_mr_inst] Storing MRW MA=2 OP=0xbb CS=0xf at row addr=0xe
                          '{ step_type : REG_WRITE, reg_addr : 32'h4101d, value : 32'h0}, //phyinit_io_write: 0x4101c, 0xc158
                          '{ step_type : REG_WRITE, reg_addr : 32'h4101e, value : 32'hddc8}, //phyinit_io_write: 0x4101d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4101f, value : 32'h0}, //phyinit_io_write: 0x4101e, 0xddc8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41020, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41021, value : 32'h4b000000}, //phyinit_io_write: 0x41020, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41022, value : 32'h0}, //phyinit_io_write: 0x41021, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41023, value : 32'h0}, //phyinit_io_write: 0x41022, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41024, value : 32'hc1d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=3 OP=0xe CS=0xf at row addr=0x12
                          '{ step_type : REG_WRITE, reg_addr : 32'h41025, value : 32'h0}, //phyinit_io_write: 0x41024, 0xc1d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41026, value : 32'hc708}, //phyinit_io_write: 0x41025, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41027, value : 32'h0}, //phyinit_io_write: 0x41026, 0xc708
                          '{ step_type : REG_WRITE, reg_addr : 32'h41028, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41029, value : 32'h4b000000}, //phyinit_io_write: 0x41028, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4102a, value : 32'h0}, //phyinit_io_write: 0x41029, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4102b, value : 32'h0}, //phyinit_io_write: 0x4102a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4102c, value : 32'hc558}, //[dwc_ddrphy_mr_inst] Storing MRW MA=10 OP=0x54 CS=0xf at row addr=0x16
                          '{ step_type : REG_WRITE, reg_addr : 32'h4102d, value : 32'h0}, //phyinit_io_write: 0x4102c, 0xc558
                          '{ step_type : REG_WRITE, reg_addr : 32'h4102e, value : 32'hea08}, //phyinit_io_write: 0x4102d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4102f, value : 32'h0}, //phyinit_io_write: 0x4102e, 0xea08
                          '{ step_type : REG_WRITE, reg_addr : 32'h41030, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41031, value : 32'h4b000000}, //phyinit_io_write: 0x41030, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41032, value : 32'h0}, //phyinit_io_write: 0x41031, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41033, value : 32'h0}, //phyinit_io_write: 0x41032, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41034, value : 32'hc5d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=11 OP=0x44 CS=0xf at row addr=0x1a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41035, value : 32'h0}, //phyinit_io_write: 0x41034, 0xc5d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41036, value : 32'he208}, //phyinit_io_write: 0x41035, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41037, value : 32'h0}, //phyinit_io_write: 0x41036, 0xe208
                          '{ step_type : REG_WRITE, reg_addr : 32'h41038, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41039, value : 32'h4b000000}, //phyinit_io_write: 0x41038, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4103a, value : 32'h0}, //phyinit_io_write: 0x41039, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4103b, value : 32'h0}, //phyinit_io_write: 0x4103a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4103c, value : 32'h48d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=17 OP=0x84 CS=0x5 at row addr=0x1e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4103d, value : 32'h0}, //phyinit_io_write: 0x4103c, 0x48d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4103e, value : 32'h4248}, //phyinit_io_write: 0x4103d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4103f, value : 32'h0}, //phyinit_io_write: 0x4103e, 0x4248
                          '{ step_type : REG_WRITE, reg_addr : 32'h41040, value : 32'h88d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=17 OP=0xac CS=0xa at row addr=0x20
                          '{ step_type : REG_WRITE, reg_addr : 32'h41041, value : 32'h0}, //phyinit_io_write: 0x41040, 0x88d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41042, value : 32'h9648}, //phyinit_io_write: 0x41041, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41043, value : 32'h0}, //phyinit_io_write: 0x41042, 0x9648
                          '{ step_type : REG_WRITE, reg_addr : 32'h41044, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41045, value : 32'h4b000000}, //phyinit_io_write: 0x41044, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41046, value : 32'h0}, //phyinit_io_write: 0x41045, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41047, value : 32'h0}, //phyinit_io_write: 0x41046, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41048, value : 32'hca58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=20 OP=0x2 CS=0xf at row addr=0x24
                          '{ step_type : REG_WRITE, reg_addr : 32'h41049, value : 32'h0}, //phyinit_io_write: 0x41048, 0xca58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4104a, value : 32'hc108}, //phyinit_io_write: 0x41049, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4104b, value : 32'h0}, //phyinit_io_write: 0x4104a, 0xc108
                          '{ step_type : REG_WRITE, reg_addr : 32'h4104c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4104d, value : 32'h4b000000}, //phyinit_io_write: 0x4104c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4104e, value : 32'h0}, //phyinit_io_write: 0x4104d, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4104f, value : 32'h0}, //phyinit_io_write: 0x4104e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41050, value : 32'hcb58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=22 OP=0x0 CS=0xf at row addr=0x28
                          '{ step_type : REG_WRITE, reg_addr : 32'h41051, value : 32'h0}, //phyinit_io_write: 0x41050, 0xcb58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41052, value : 32'hc008}, //phyinit_io_write: 0x41051, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41053, value : 32'h0}, //phyinit_io_write: 0x41052, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41054, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41055, value : 32'h4b000000}, //phyinit_io_write: 0x41054, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41056, value : 32'h0}, //phyinit_io_write: 0x41055, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41057, value : 32'h0}, //phyinit_io_write: 0x41056, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41058, value : 32'hd4d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=41 OP=0x60 CS=0xf at row addr=0x2c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41059, value : 32'h0}, //phyinit_io_write: 0x41058, 0xd4d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4105a, value : 32'hf008}, //phyinit_io_write: 0x41059, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4105b, value : 32'h0}, //phyinit_io_write: 0x4105a, 0xf008
                          '{ step_type : REG_WRITE, reg_addr : 32'h4105c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4105d, value : 32'h4b000000}, //phyinit_io_write: 0x4105c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4105e, value : 32'h0}, //phyinit_io_write: 0x4105d, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4105f, value : 32'h0}, //phyinit_io_write: 0x4105e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41060, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=58 at row addr=0x30
                          '{ step_type : REG_WRITE, reg_addr : 32'h41061, value : 32'h0}, //phyinit_io_write: 0x41060, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41062, value : 32'h0}, //phyinit_io_write: 0x41061, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41063, value : 32'h0}, //phyinit_io_write: 0x41062, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41064, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x32
                          '{ step_type : REG_WRITE, reg_addr : 32'h41065, value : 32'h0}, //phyinit_io_write: 0x41064, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h41066, value : 32'h6808}, //phyinit_io_write: 0x41065, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41067, value : 32'h0}, //phyinit_io_write: 0x41066, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41068, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x34
                          '{ step_type : REG_WRITE, reg_addr : 32'h41069, value : 32'h0}, //phyinit_io_write: 0x41068, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h4106a, value : 32'ha808}, //phyinit_io_write: 0x41069, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4106b, value : 32'h0}, //phyinit_io_write: 0x4106a, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h4106c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4106d, value : 32'h4b000000}, //phyinit_io_write: 0x4106c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4106e, value : 32'h0}, //phyinit_io_write: 0x4106d, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4106f, value : 32'h0}, //phyinit_io_write: 0x4106e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41070, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x38
                          '{ step_type : REG_WRITE, reg_addr : 32'h41071, value : 32'h0}, //phyinit_io_write: 0x41070, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h41072, value : 32'h6808}, //phyinit_io_write: 0x41071, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41073, value : 32'h0}, //phyinit_io_write: 0x41072, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41074, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x3a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41075, value : 32'h0}, //phyinit_io_write: 0x41074, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h41076, value : 32'ha808}, //phyinit_io_write: 0x41075, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41077, value : 32'h0}, //phyinit_io_write: 0x41076, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41078, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41079, value : 32'h4b000000}, //phyinit_io_write: 0x41078, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4107a, value : 32'h0}, //phyinit_io_write: 0x41079, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4107b, value : 32'h0}, //phyinit_io_write: 0x4107a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4107c, value : 32'h4758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0x5 at row addr=0x3e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4107d, value : 32'h0}, //phyinit_io_write: 0x4107c, 0x4758
                          '{ step_type : REG_WRITE, reg_addr : 32'h4107e, value : 32'h6808}, //phyinit_io_write: 0x4107d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4107f, value : 32'h0}, //phyinit_io_write: 0x4107e, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41080, value : 32'h8758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0xa at row addr=0x40
                          '{ step_type : REG_WRITE, reg_addr : 32'h41081, value : 32'h0}, //phyinit_io_write: 0x41080, 0x8758
                          '{ step_type : REG_WRITE, reg_addr : 32'h41082, value : 32'ha808}, //phyinit_io_write: 0x41081, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41083, value : 32'h0}, //phyinit_io_write: 0x41082, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41084, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41085, value : 32'h4b000000}, //phyinit_io_write: 0x41084, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41086, value : 32'h0}, //phyinit_io_write: 0x41085, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41087, value : 32'h0}, //phyinit_io_write: 0x41086, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41088, value : 32'h47d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0x5 at row addr=0x44
                          '{ step_type : REG_WRITE, reg_addr : 32'h41089, value : 32'h0}, //phyinit_io_write: 0x41088, 0x47d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4108a, value : 32'h6808}, //phyinit_io_write: 0x41089, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4108b, value : 32'h0}, //phyinit_io_write: 0x4108a, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h4108c, value : 32'h87d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0xa at row addr=0x46
                          '{ step_type : REG_WRITE, reg_addr : 32'h4108d, value : 32'h0}, //phyinit_io_write: 0x4108c, 0x87d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4108e, value : 32'ha808}, //phyinit_io_write: 0x4108d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4108f, value : 32'h0}, //phyinit_io_write: 0x4108e, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41090, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41091, value : 32'h4b000000}, //phyinit_io_write: 0x41090, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41092, value : 32'h0}, //phyinit_io_write: 0x41091, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41093, value : 32'h0}, //phyinit_io_write: 0x41092, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41094, value : 32'h4c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0x5 at row addr=0x4a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41095, value : 32'h0}, //phyinit_io_write: 0x41094, 0x4c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41096, value : 32'h4008}, //phyinit_io_write: 0x41095, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41097, value : 32'h0}, //phyinit_io_write: 0x41096, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41098, value : 32'h8c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0xa at row addr=0x4c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41099, value : 32'h0}, //phyinit_io_write: 0x41098, 0x8c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4109a, value : 32'h8008}, //phyinit_io_write: 0x41099, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4109b, value : 32'h0}, //phyinit_io_write: 0x4109a, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h4109c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h4109d, value : 32'h4b000000}, //phyinit_io_write: 0x4109c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4109e, value : 32'h0}, //phyinit_io_write: 0x4109d, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4109f, value : 32'h0}, //phyinit_io_write: 0x4109e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a0, value : 32'h4f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0x5 at row addr=0x50
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a1, value : 32'h0}, //phyinit_io_write: 0x410a0, 0x4f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a2, value : 32'h4008}, //phyinit_io_write: 0x410a1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a3, value : 32'h0}, //phyinit_io_write: 0x410a2, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a4, value : 32'h8f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0xa at row addr=0x52
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a5, value : 32'h0}, //phyinit_io_write: 0x410a4, 0x8f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a6, value : 32'h8008}, //phyinit_io_write: 0x410a5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a7, value : 32'h0}, //phyinit_io_write: 0x410a6, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a8, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h410a9, value : 32'h4b000000}, //phyinit_io_write: 0x410a8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410aa, value : 32'h0}, //phyinit_io_write: 0x410a9, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ab, value : 32'h0}, //phyinit_io_write: 0x410aa, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ac, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x56
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ad, value : 32'h0}, //phyinit_io_write: 0x410ac, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ae, value : 32'h0}, //phyinit_io_write: 0x410ad, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410af, value : 32'h0}, //phyinit_io_write: 0x410ae, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b0, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x58
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b1, value : 32'h0}, //phyinit_io_write: 0x410b0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b2, value : 32'h0}, //phyinit_io_write: 0x410b1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b3, value : 32'h0}, //phyinit_io_write: 0x410b2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b4, value : 32'h0}, //phyinit_io_write: 0x410b3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b5, value : 32'h0}, //phyinit_io_write: 0x410b4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b6, value : 32'h0}, //phyinit_io_write: 0x410b5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b7, value : 32'h0}, //phyinit_io_write: 0x410b6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b8, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x5c
                          '{ step_type : REG_WRITE, reg_addr : 32'h410b9, value : 32'h0}, //phyinit_io_write: 0x410b8, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ba, value : 32'h6808}, //phyinit_io_write: 0x410b9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410bb, value : 32'h0}, //phyinit_io_write: 0x410ba, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h410bc, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x5e
                          '{ step_type : REG_WRITE, reg_addr : 32'h410bd, value : 32'h0}, //phyinit_io_write: 0x410bc, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h410be, value : 32'ha808}, //phyinit_io_write: 0x410bd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410bf, value : 32'h0}, //phyinit_io_write: 0x410be, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c0, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c1, value : 32'h4b000000}, //phyinit_io_write: 0x410c0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c2, value : 32'h0}, //phyinit_io_write: 0x410c1, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c3, value : 32'h0}, //phyinit_io_write: 0x410c2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c4, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x62
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c5, value : 32'h0}, //phyinit_io_write: 0x410c4, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c6, value : 32'h6808}, //phyinit_io_write: 0x410c5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c7, value : 32'h0}, //phyinit_io_write: 0x410c6, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c8, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x64
                          '{ step_type : REG_WRITE, reg_addr : 32'h410c9, value : 32'h0}, //phyinit_io_write: 0x410c8, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ca, value : 32'ha808}, //phyinit_io_write: 0x410c9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410cb, value : 32'h0}, //phyinit_io_write: 0x410ca, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h410cc, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h410cd, value : 32'h4b000000}, //phyinit_io_write: 0x410cc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ce, value : 32'h0}, //phyinit_io_write: 0x410cd, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h410cf, value : 32'h0}, //phyinit_io_write: 0x410ce, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d0, value : 32'h4758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0x5 at row addr=0x68
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d1, value : 32'h0}, //phyinit_io_write: 0x410d0, 0x4758
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d2, value : 32'h6808}, //phyinit_io_write: 0x410d1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d3, value : 32'h0}, //phyinit_io_write: 0x410d2, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d4, value : 32'h8758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0xa at row addr=0x6a
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d5, value : 32'h0}, //phyinit_io_write: 0x410d4, 0x8758
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d6, value : 32'ha808}, //phyinit_io_write: 0x410d5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d7, value : 32'h0}, //phyinit_io_write: 0x410d6, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d8, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h410d9, value : 32'h4b000000}, //phyinit_io_write: 0x410d8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410da, value : 32'h0}, //phyinit_io_write: 0x410d9, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h410db, value : 32'h0}, //phyinit_io_write: 0x410da, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410dc, value : 32'h47d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0x5 at row addr=0x6e
                          '{ step_type : REG_WRITE, reg_addr : 32'h410dd, value : 32'h0}, //phyinit_io_write: 0x410dc, 0x47d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h410de, value : 32'h6808}, //phyinit_io_write: 0x410dd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410df, value : 32'h0}, //phyinit_io_write: 0x410de, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e0, value : 32'h87d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0xa at row addr=0x70
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e1, value : 32'h0}, //phyinit_io_write: 0x410e0, 0x87d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e2, value : 32'ha808}, //phyinit_io_write: 0x410e1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e3, value : 32'h0}, //phyinit_io_write: 0x410e2, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e4, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e5, value : 32'h4b000000}, //phyinit_io_write: 0x410e4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e6, value : 32'h0}, //phyinit_io_write: 0x410e5, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e7, value : 32'h0}, //phyinit_io_write: 0x410e6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e8, value : 32'h4c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0x5 at row addr=0x74
                          '{ step_type : REG_WRITE, reg_addr : 32'h410e9, value : 32'h0}, //phyinit_io_write: 0x410e8, 0x4c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ea, value : 32'h4008}, //phyinit_io_write: 0x410e9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410eb, value : 32'h0}, //phyinit_io_write: 0x410ea, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ec, value : 32'h8c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0xa at row addr=0x76
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ed, value : 32'h0}, //phyinit_io_write: 0x410ec, 0x8c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ee, value : 32'h8008}, //phyinit_io_write: 0x410ed, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ef, value : 32'h0}, //phyinit_io_write: 0x410ee, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f0, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f1, value : 32'h4b000000}, //phyinit_io_write: 0x410f0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f2, value : 32'h0}, //phyinit_io_write: 0x410f1, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f3, value : 32'h0}, //phyinit_io_write: 0x410f2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f4, value : 32'h4f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0x5 at row addr=0x7a
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f5, value : 32'h0}, //phyinit_io_write: 0x410f4, 0x4f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f6, value : 32'h4008}, //phyinit_io_write: 0x410f5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f7, value : 32'h0}, //phyinit_io_write: 0x410f6, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f8, value : 32'h8f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0xa at row addr=0x7c
                          '{ step_type : REG_WRITE, reg_addr : 32'h410f9, value : 32'h0}, //phyinit_io_write: 0x410f8, 0x8f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h410fa, value : 32'h8008}, //phyinit_io_write: 0x410f9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410fb, value : 32'h0}, //phyinit_io_write: 0x410fa, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h410fc, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 8 cnt = 4
                          '{ step_type : REG_WRITE, reg_addr : 32'h410fd, value : 32'h4b000000}, //phyinit_io_write: 0x410fc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h410fe, value : 32'h0}, //phyinit_io_write: 0x410fd, 0x4b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h410ff, value : 32'h0}, //phyinit_io_write: 0x410fe, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41100, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x80
                          '{ step_type : REG_WRITE, reg_addr : 32'h41101, value : 32'h0}, //phyinit_io_write: 0x41100, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41102, value : 32'h0}, //phyinit_io_write: 0x41101, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41103, value : 32'h0}, //phyinit_io_write: 0x41102, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41104, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x82
                          '{ step_type : REG_WRITE, reg_addr : 32'h41105, value : 32'h0}, //phyinit_io_write: 0x41104, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41106, value : 32'h0}, //phyinit_io_write: 0x41105, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41107, value : 32'h0}, //phyinit_io_write: 0x41106, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41108, value : 32'h0}, //phyinit_io_write: 0x41107, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41109, value : 32'h0}, //phyinit_io_write: 0x41108, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4110a, value : 32'h0}, //phyinit_io_write: 0x41109, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4110b, value : 32'h0}, //phyinit_io_write: 0x4110a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h170145, value : 32'h2}, //[loadAcsmMRW] Pstate=1, Programming ACSMRptCntOverride to 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4110c, value : 32'hc9d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=19 OP=0x0 CS=0xf at row addr=0x86
                          '{ step_type : REG_WRITE, reg_addr : 32'h4110d, value : 32'h0}, //phyinit_io_write: 0x4110c, 0xc9d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4110e, value : 32'hc008}, //phyinit_io_write: 0x4110d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4110f, value : 32'h0}, //phyinit_io_write: 0x4110e, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41110, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41111, value : 32'h3b000000}, //phyinit_io_write: 0x41110, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41112, value : 32'h0}, //phyinit_io_write: 0x41111, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41113, value : 32'h0}, //phyinit_io_write: 0x41112, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41114, value : 32'hc958}, //[dwc_ddrphy_mr_inst] Storing MRW MA=18 OP=0x0 CS=0xf at row addr=0x8a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41115, value : 32'h0}, //phyinit_io_write: 0x41114, 0xc958
                          '{ step_type : REG_WRITE, reg_addr : 32'h41116, value : 32'hc008}, //phyinit_io_write: 0x41115, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41117, value : 32'h0}, //phyinit_io_write: 0x41116, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41118, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41119, value : 32'h3b000000}, //phyinit_io_write: 0x41118, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4111a, value : 32'h0}, //phyinit_io_write: 0x41119, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4111b, value : 32'h0}, //phyinit_io_write: 0x4111a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4111c, value : 32'hc0d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=1 OP=0x80 CS=0xf at row addr=0x8e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4111d, value : 32'h0}, //phyinit_io_write: 0x4111c, 0xc0d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4111e, value : 32'hc048}, //phyinit_io_write: 0x4111d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4111f, value : 32'h0}, //phyinit_io_write: 0x4111e, 0xc048
                          '{ step_type : REG_WRITE, reg_addr : 32'h41120, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41121, value : 32'h3b000000}, //phyinit_io_write: 0x41120, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41122, value : 32'h0}, //phyinit_io_write: 0x41121, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41123, value : 32'h0}, //phyinit_io_write: 0x41122, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41124, value : 32'hc158}, //[dwc_ddrphy_mr_inst] Storing MRW MA=2 OP=0x88 CS=0xf at row addr=0x92
                          '{ step_type : REG_WRITE, reg_addr : 32'h41125, value : 32'h0}, //phyinit_io_write: 0x41124, 0xc158
                          '{ step_type : REG_WRITE, reg_addr : 32'h41126, value : 32'hc448}, //phyinit_io_write: 0x41125, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41127, value : 32'h0}, //phyinit_io_write: 0x41126, 0xc448
                          '{ step_type : REG_WRITE, reg_addr : 32'h41128, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41129, value : 32'h3b000000}, //phyinit_io_write: 0x41128, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4112a, value : 32'h0}, //phyinit_io_write: 0x41129, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4112b, value : 32'h0}, //phyinit_io_write: 0x4112a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4112c, value : 32'hc1d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=3 OP=0xe CS=0xf at row addr=0x96
                          '{ step_type : REG_WRITE, reg_addr : 32'h4112d, value : 32'h0}, //phyinit_io_write: 0x4112c, 0xc1d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4112e, value : 32'hc708}, //phyinit_io_write: 0x4112d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4112f, value : 32'h0}, //phyinit_io_write: 0x4112e, 0xc708
                          '{ step_type : REG_WRITE, reg_addr : 32'h41130, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41131, value : 32'h3b000000}, //phyinit_io_write: 0x41130, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41132, value : 32'h0}, //phyinit_io_write: 0x41131, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41133, value : 32'h0}, //phyinit_io_write: 0x41132, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41134, value : 32'hc558}, //[dwc_ddrphy_mr_inst] Storing MRW MA=10 OP=0x54 CS=0xf at row addr=0x9a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41135, value : 32'h0}, //phyinit_io_write: 0x41134, 0xc558
                          '{ step_type : REG_WRITE, reg_addr : 32'h41136, value : 32'hea08}, //phyinit_io_write: 0x41135, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41137, value : 32'h0}, //phyinit_io_write: 0x41136, 0xea08
                          '{ step_type : REG_WRITE, reg_addr : 32'h41138, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41139, value : 32'h3b000000}, //phyinit_io_write: 0x41138, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4113a, value : 32'h0}, //phyinit_io_write: 0x41139, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4113b, value : 32'h0}, //phyinit_io_write: 0x4113a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4113c, value : 32'hc5d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=11 OP=0x44 CS=0xf at row addr=0x9e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4113d, value : 32'h0}, //phyinit_io_write: 0x4113c, 0xc5d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4113e, value : 32'he208}, //phyinit_io_write: 0x4113d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4113f, value : 32'h0}, //phyinit_io_write: 0x4113e, 0xe208
                          '{ step_type : REG_WRITE, reg_addr : 32'h41140, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41141, value : 32'h3b000000}, //phyinit_io_write: 0x41140, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41142, value : 32'h0}, //phyinit_io_write: 0x41141, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41143, value : 32'h0}, //phyinit_io_write: 0x41142, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41144, value : 32'h48d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=17 OP=0x84 CS=0x5 at row addr=0xa2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41145, value : 32'h0}, //phyinit_io_write: 0x41144, 0x48d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41146, value : 32'h4248}, //phyinit_io_write: 0x41145, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41147, value : 32'h0}, //phyinit_io_write: 0x41146, 0x4248
                          '{ step_type : REG_WRITE, reg_addr : 32'h41148, value : 32'h88d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=17 OP=0xac CS=0xa at row addr=0xa4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41149, value : 32'h0}, //phyinit_io_write: 0x41148, 0x88d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4114a, value : 32'h9648}, //phyinit_io_write: 0x41149, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4114b, value : 32'h0}, //phyinit_io_write: 0x4114a, 0x9648
                          '{ step_type : REG_WRITE, reg_addr : 32'h4114c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h4114d, value : 32'h3b000000}, //phyinit_io_write: 0x4114c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4114e, value : 32'h0}, //phyinit_io_write: 0x4114d, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4114f, value : 32'h0}, //phyinit_io_write: 0x4114e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41150, value : 32'hca58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=20 OP=0x2 CS=0xf at row addr=0xa8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41151, value : 32'h0}, //phyinit_io_write: 0x41150, 0xca58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41152, value : 32'hc108}, //phyinit_io_write: 0x41151, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41153, value : 32'h0}, //phyinit_io_write: 0x41152, 0xc108
                          '{ step_type : REG_WRITE, reg_addr : 32'h41154, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41155, value : 32'h3b000000}, //phyinit_io_write: 0x41154, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41156, value : 32'h0}, //phyinit_io_write: 0x41155, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41157, value : 32'h0}, //phyinit_io_write: 0x41156, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41158, value : 32'hcb58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=22 OP=0x0 CS=0xf at row addr=0xac
                          '{ step_type : REG_WRITE, reg_addr : 32'h41159, value : 32'h0}, //phyinit_io_write: 0x41158, 0xcb58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4115a, value : 32'hc008}, //phyinit_io_write: 0x41159, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4115b, value : 32'h0}, //phyinit_io_write: 0x4115a, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h4115c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h4115d, value : 32'h3b000000}, //phyinit_io_write: 0x4115c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4115e, value : 32'h0}, //phyinit_io_write: 0x4115d, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4115f, value : 32'h0}, //phyinit_io_write: 0x4115e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41160, value : 32'hd4d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=41 OP=0x60 CS=0xf at row addr=0xb0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41161, value : 32'h0}, //phyinit_io_write: 0x41160, 0xd4d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41162, value : 32'hf008}, //phyinit_io_write: 0x41161, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41163, value : 32'h0}, //phyinit_io_write: 0x41162, 0xf008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41164, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41165, value : 32'h3b000000}, //phyinit_io_write: 0x41164, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41166, value : 32'h0}, //phyinit_io_write: 0x41165, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41167, value : 32'h0}, //phyinit_io_write: 0x41166, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41168, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=58 at row addr=0xb4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41169, value : 32'h0}, //phyinit_io_write: 0x41168, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4116a, value : 32'h0}, //phyinit_io_write: 0x41169, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4116b, value : 32'h0}, //phyinit_io_write: 0x4116a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4116c, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0xb6
                          '{ step_type : REG_WRITE, reg_addr : 32'h4116d, value : 32'h0}, //phyinit_io_write: 0x4116c, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h4116e, value : 32'h6808}, //phyinit_io_write: 0x4116d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4116f, value : 32'h0}, //phyinit_io_write: 0x4116e, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41170, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0xb8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41171, value : 32'h0}, //phyinit_io_write: 0x41170, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h41172, value : 32'ha808}, //phyinit_io_write: 0x41171, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41173, value : 32'h0}, //phyinit_io_write: 0x41172, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41174, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41175, value : 32'h3b000000}, //phyinit_io_write: 0x41174, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41176, value : 32'h0}, //phyinit_io_write: 0x41175, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41177, value : 32'h0}, //phyinit_io_write: 0x41176, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41178, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0xbc
                          '{ step_type : REG_WRITE, reg_addr : 32'h41179, value : 32'h0}, //phyinit_io_write: 0x41178, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h4117a, value : 32'h6808}, //phyinit_io_write: 0x41179, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4117b, value : 32'h0}, //phyinit_io_write: 0x4117a, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h4117c, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0xbe
                          '{ step_type : REG_WRITE, reg_addr : 32'h4117d, value : 32'h0}, //phyinit_io_write: 0x4117c, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h4117e, value : 32'ha808}, //phyinit_io_write: 0x4117d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4117f, value : 32'h0}, //phyinit_io_write: 0x4117e, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41180, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41181, value : 32'h3b000000}, //phyinit_io_write: 0x41180, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41182, value : 32'h0}, //phyinit_io_write: 0x41181, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41183, value : 32'h0}, //phyinit_io_write: 0x41182, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41184, value : 32'h4758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0x5 at row addr=0xc2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41185, value : 32'h0}, //phyinit_io_write: 0x41184, 0x4758
                          '{ step_type : REG_WRITE, reg_addr : 32'h41186, value : 32'h6808}, //phyinit_io_write: 0x41185, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41187, value : 32'h0}, //phyinit_io_write: 0x41186, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41188, value : 32'h8758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0xa at row addr=0xc4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41189, value : 32'h0}, //phyinit_io_write: 0x41188, 0x8758
                          '{ step_type : REG_WRITE, reg_addr : 32'h4118a, value : 32'ha808}, //phyinit_io_write: 0x41189, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4118b, value : 32'h0}, //phyinit_io_write: 0x4118a, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h4118c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h4118d, value : 32'h3b000000}, //phyinit_io_write: 0x4118c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4118e, value : 32'h0}, //phyinit_io_write: 0x4118d, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4118f, value : 32'h0}, //phyinit_io_write: 0x4118e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41190, value : 32'h47d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0x5 at row addr=0xc8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41191, value : 32'h0}, //phyinit_io_write: 0x41190, 0x47d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41192, value : 32'h6808}, //phyinit_io_write: 0x41191, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41193, value : 32'h0}, //phyinit_io_write: 0x41192, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41194, value : 32'h87d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0xa at row addr=0xca
                          '{ step_type : REG_WRITE, reg_addr : 32'h41195, value : 32'h0}, //phyinit_io_write: 0x41194, 0x87d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41196, value : 32'ha808}, //phyinit_io_write: 0x41195, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41197, value : 32'h0}, //phyinit_io_write: 0x41196, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41198, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41199, value : 32'h3b000000}, //phyinit_io_write: 0x41198, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4119a, value : 32'h0}, //phyinit_io_write: 0x41199, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4119b, value : 32'h0}, //phyinit_io_write: 0x4119a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4119c, value : 32'h4c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0x5 at row addr=0xce
                          '{ step_type : REG_WRITE, reg_addr : 32'h4119d, value : 32'h0}, //phyinit_io_write: 0x4119c, 0x4c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4119e, value : 32'h4008}, //phyinit_io_write: 0x4119d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4119f, value : 32'h0}, //phyinit_io_write: 0x4119e, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a0, value : 32'h8c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0xa at row addr=0xd0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a1, value : 32'h0}, //phyinit_io_write: 0x411a0, 0x8c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a2, value : 32'h8008}, //phyinit_io_write: 0x411a1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a3, value : 32'h0}, //phyinit_io_write: 0x411a2, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a4, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a5, value : 32'h3b000000}, //phyinit_io_write: 0x411a4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a6, value : 32'h0}, //phyinit_io_write: 0x411a5, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a7, value : 32'h0}, //phyinit_io_write: 0x411a6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a8, value : 32'h4f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0x5 at row addr=0xd4
                          '{ step_type : REG_WRITE, reg_addr : 32'h411a9, value : 32'h0}, //phyinit_io_write: 0x411a8, 0x4f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h411aa, value : 32'h4008}, //phyinit_io_write: 0x411a9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ab, value : 32'h0}, //phyinit_io_write: 0x411aa, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ac, value : 32'h8f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0xa at row addr=0xd6
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ad, value : 32'h0}, //phyinit_io_write: 0x411ac, 0x8f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ae, value : 32'h8008}, //phyinit_io_write: 0x411ad, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411af, value : 32'h0}, //phyinit_io_write: 0x411ae, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b0, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b1, value : 32'h3b000000}, //phyinit_io_write: 0x411b0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b2, value : 32'h0}, //phyinit_io_write: 0x411b1, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b3, value : 32'h0}, //phyinit_io_write: 0x411b2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b4, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0xda
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b5, value : 32'h0}, //phyinit_io_write: 0x411b4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b6, value : 32'h0}, //phyinit_io_write: 0x411b5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b7, value : 32'h0}, //phyinit_io_write: 0x411b6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b8, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0xdc
                          '{ step_type : REG_WRITE, reg_addr : 32'h411b9, value : 32'h0}, //phyinit_io_write: 0x411b8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ba, value : 32'h0}, //phyinit_io_write: 0x411b9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411bb, value : 32'h0}, //phyinit_io_write: 0x411ba, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411bc, value : 32'h0}, //phyinit_io_write: 0x411bb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411bd, value : 32'h0}, //phyinit_io_write: 0x411bc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411be, value : 32'h0}, //phyinit_io_write: 0x411bd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411bf, value : 32'h0}, //phyinit_io_write: 0x411be, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c0, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0xe0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c1, value : 32'h0}, //phyinit_io_write: 0x411c0, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c2, value : 32'h6808}, //phyinit_io_write: 0x411c1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c3, value : 32'h0}, //phyinit_io_write: 0x411c2, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c4, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0xe2
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c5, value : 32'h0}, //phyinit_io_write: 0x411c4, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c6, value : 32'ha808}, //phyinit_io_write: 0x411c5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c7, value : 32'h0}, //phyinit_io_write: 0x411c6, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c8, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h411c9, value : 32'h3b000000}, //phyinit_io_write: 0x411c8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ca, value : 32'h0}, //phyinit_io_write: 0x411c9, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h411cb, value : 32'h0}, //phyinit_io_write: 0x411ca, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411cc, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0xe6
                          '{ step_type : REG_WRITE, reg_addr : 32'h411cd, value : 32'h0}, //phyinit_io_write: 0x411cc, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ce, value : 32'h6808}, //phyinit_io_write: 0x411cd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411cf, value : 32'h0}, //phyinit_io_write: 0x411ce, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d0, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0xe8
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d1, value : 32'h0}, //phyinit_io_write: 0x411d0, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d2, value : 32'ha808}, //phyinit_io_write: 0x411d1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d3, value : 32'h0}, //phyinit_io_write: 0x411d2, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d4, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d5, value : 32'h3b000000}, //phyinit_io_write: 0x411d4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d6, value : 32'h0}, //phyinit_io_write: 0x411d5, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d7, value : 32'h0}, //phyinit_io_write: 0x411d6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d8, value : 32'h4758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0x5 at row addr=0xec
                          '{ step_type : REG_WRITE, reg_addr : 32'h411d9, value : 32'h0}, //phyinit_io_write: 0x411d8, 0x4758
                          '{ step_type : REG_WRITE, reg_addr : 32'h411da, value : 32'h6808}, //phyinit_io_write: 0x411d9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411db, value : 32'h0}, //phyinit_io_write: 0x411da, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h411dc, value : 32'h8758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0xa at row addr=0xee
                          '{ step_type : REG_WRITE, reg_addr : 32'h411dd, value : 32'h0}, //phyinit_io_write: 0x411dc, 0x8758
                          '{ step_type : REG_WRITE, reg_addr : 32'h411de, value : 32'ha808}, //phyinit_io_write: 0x411dd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411df, value : 32'h0}, //phyinit_io_write: 0x411de, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e0, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e1, value : 32'h3b000000}, //phyinit_io_write: 0x411e0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e2, value : 32'h0}, //phyinit_io_write: 0x411e1, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e3, value : 32'h0}, //phyinit_io_write: 0x411e2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e4, value : 32'h47d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0x5 at row addr=0xf2
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e5, value : 32'h0}, //phyinit_io_write: 0x411e4, 0x47d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e6, value : 32'h6808}, //phyinit_io_write: 0x411e5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e7, value : 32'h0}, //phyinit_io_write: 0x411e6, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e8, value : 32'h87d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0xa at row addr=0xf4
                          '{ step_type : REG_WRITE, reg_addr : 32'h411e9, value : 32'h0}, //phyinit_io_write: 0x411e8, 0x87d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ea, value : 32'ha808}, //phyinit_io_write: 0x411e9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411eb, value : 32'h0}, //phyinit_io_write: 0x411ea, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ec, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ed, value : 32'h3b000000}, //phyinit_io_write: 0x411ec, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ee, value : 32'h0}, //phyinit_io_write: 0x411ed, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ef, value : 32'h0}, //phyinit_io_write: 0x411ee, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f0, value : 32'h4c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0x5 at row addr=0xf8
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f1, value : 32'h0}, //phyinit_io_write: 0x411f0, 0x4c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f2, value : 32'h4008}, //phyinit_io_write: 0x411f1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f3, value : 32'h0}, //phyinit_io_write: 0x411f2, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f4, value : 32'h8c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0xa at row addr=0xfa
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f5, value : 32'h0}, //phyinit_io_write: 0x411f4, 0x8c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f6, value : 32'h8008}, //phyinit_io_write: 0x411f5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f7, value : 32'h0}, //phyinit_io_write: 0x411f6, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f8, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h411f9, value : 32'h3b000000}, //phyinit_io_write: 0x411f8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411fa, value : 32'h0}, //phyinit_io_write: 0x411f9, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h411fb, value : 32'h0}, //phyinit_io_write: 0x411fa, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411fc, value : 32'h4f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0x5 at row addr=0xfe
                          '{ step_type : REG_WRITE, reg_addr : 32'h411fd, value : 32'h0}, //phyinit_io_write: 0x411fc, 0x4f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h411fe, value : 32'h4008}, //phyinit_io_write: 0x411fd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h411ff, value : 32'h0}, //phyinit_io_write: 0x411fe, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41200, value : 32'h8f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0xa at row addr=0x100
                          '{ step_type : REG_WRITE, reg_addr : 32'h41201, value : 32'h0}, //phyinit_io_write: 0x41200, 0x8f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41202, value : 32'h8008}, //phyinit_io_write: 0x41201, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41203, value : 32'h0}, //phyinit_io_write: 0x41202, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41204, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 7 cnt = 3
                          '{ step_type : REG_WRITE, reg_addr : 32'h41205, value : 32'h3b000000}, //phyinit_io_write: 0x41204, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41206, value : 32'h0}, //phyinit_io_write: 0x41205, 0x3b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41207, value : 32'h0}, //phyinit_io_write: 0x41206, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41208, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x104
                          '{ step_type : REG_WRITE, reg_addr : 32'h41209, value : 32'h0}, //phyinit_io_write: 0x41208, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4120a, value : 32'h0}, //phyinit_io_write: 0x41209, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4120b, value : 32'h0}, //phyinit_io_write: 0x4120a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4120c, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x106
                          '{ step_type : REG_WRITE, reg_addr : 32'h4120d, value : 32'h0}, //phyinit_io_write: 0x4120c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4120e, value : 32'h0}, //phyinit_io_write: 0x4120d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4120f, value : 32'h0}, //phyinit_io_write: 0x4120e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41210, value : 32'h0}, //phyinit_io_write: 0x4120f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41211, value : 32'h0}, //phyinit_io_write: 0x41210, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41212, value : 32'h0}, //phyinit_io_write: 0x41211, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41213, value : 32'h0}, //phyinit_io_write: 0x41212, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h270145, value : 32'h1}, //[loadAcsmMRW] Pstate=2, Programming ACSMRptCntOverride to 1
                          '{ step_type : REG_WRITE, reg_addr : 32'h41214, value : 32'hc9d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=19 OP=0x0 CS=0xf at row addr=0x10a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41215, value : 32'h0}, //phyinit_io_write: 0x41214, 0xc9d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41216, value : 32'hc008}, //phyinit_io_write: 0x41215, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41217, value : 32'h0}, //phyinit_io_write: 0x41216, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41218, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41219, value : 32'h2b000000}, //phyinit_io_write: 0x41218, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4121a, value : 32'h0}, //phyinit_io_write: 0x41219, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4121b, value : 32'h0}, //phyinit_io_write: 0x4121a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4121c, value : 32'hc958}, //[dwc_ddrphy_mr_inst] Storing MRW MA=18 OP=0x0 CS=0xf at row addr=0x10e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4121d, value : 32'h0}, //phyinit_io_write: 0x4121c, 0xc958
                          '{ step_type : REG_WRITE, reg_addr : 32'h4121e, value : 32'hc008}, //phyinit_io_write: 0x4121d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4121f, value : 32'h0}, //phyinit_io_write: 0x4121e, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41220, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41221, value : 32'h2b000000}, //phyinit_io_write: 0x41220, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41222, value : 32'h0}, //phyinit_io_write: 0x41221, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41223, value : 32'h0}, //phyinit_io_write: 0x41222, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41224, value : 32'hc0d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=1 OP=0x50 CS=0xf at row addr=0x112
                          '{ step_type : REG_WRITE, reg_addr : 32'h41225, value : 32'h0}, //phyinit_io_write: 0x41224, 0xc0d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41226, value : 32'he808}, //phyinit_io_write: 0x41225, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41227, value : 32'h0}, //phyinit_io_write: 0x41226, 0xe808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41228, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41229, value : 32'h2b000000}, //phyinit_io_write: 0x41228, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4122a, value : 32'h0}, //phyinit_io_write: 0x41229, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4122b, value : 32'h0}, //phyinit_io_write: 0x4122a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4122c, value : 32'hc158}, //[dwc_ddrphy_mr_inst] Storing MRW MA=2 OP=0x55 CS=0xf at row addr=0x116
                          '{ step_type : REG_WRITE, reg_addr : 32'h4122d, value : 32'h0}, //phyinit_io_write: 0x4122c, 0xc158
                          '{ step_type : REG_WRITE, reg_addr : 32'h4122e, value : 32'hea88}, //phyinit_io_write: 0x4122d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4122f, value : 32'h0}, //phyinit_io_write: 0x4122e, 0xea88
                          '{ step_type : REG_WRITE, reg_addr : 32'h41230, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41231, value : 32'h2b000000}, //phyinit_io_write: 0x41230, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41232, value : 32'h0}, //phyinit_io_write: 0x41231, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41233, value : 32'h0}, //phyinit_io_write: 0x41232, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41234, value : 32'hc1d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=3 OP=0xe CS=0xf at row addr=0x11a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41235, value : 32'h0}, //phyinit_io_write: 0x41234, 0xc1d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41236, value : 32'hc708}, //phyinit_io_write: 0x41235, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41237, value : 32'h0}, //phyinit_io_write: 0x41236, 0xc708
                          '{ step_type : REG_WRITE, reg_addr : 32'h41238, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41239, value : 32'h2b000000}, //phyinit_io_write: 0x41238, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4123a, value : 32'h0}, //phyinit_io_write: 0x41239, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4123b, value : 32'h0}, //phyinit_io_write: 0x4123a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4123c, value : 32'hc558}, //[dwc_ddrphy_mr_inst] Storing MRW MA=10 OP=0x54 CS=0xf at row addr=0x11e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4123d, value : 32'h0}, //phyinit_io_write: 0x4123c, 0xc558
                          '{ step_type : REG_WRITE, reg_addr : 32'h4123e, value : 32'hea08}, //phyinit_io_write: 0x4123d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4123f, value : 32'h0}, //phyinit_io_write: 0x4123e, 0xea08
                          '{ step_type : REG_WRITE, reg_addr : 32'h41240, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41241, value : 32'h2b000000}, //phyinit_io_write: 0x41240, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41242, value : 32'h0}, //phyinit_io_write: 0x41241, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41243, value : 32'h0}, //phyinit_io_write: 0x41242, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41244, value : 32'hc5d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=11 OP=0x44 CS=0xf at row addr=0x122
                          '{ step_type : REG_WRITE, reg_addr : 32'h41245, value : 32'h0}, //phyinit_io_write: 0x41244, 0xc5d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41246, value : 32'he208}, //phyinit_io_write: 0x41245, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41247, value : 32'h0}, //phyinit_io_write: 0x41246, 0xe208
                          '{ step_type : REG_WRITE, reg_addr : 32'h41248, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41249, value : 32'h2b000000}, //phyinit_io_write: 0x41248, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4124a, value : 32'h0}, //phyinit_io_write: 0x41249, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4124b, value : 32'h0}, //phyinit_io_write: 0x4124a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4124c, value : 32'h48d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=17 OP=0x84 CS=0x5 at row addr=0x126
                          '{ step_type : REG_WRITE, reg_addr : 32'h4124d, value : 32'h0}, //phyinit_io_write: 0x4124c, 0x48d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4124e, value : 32'h4248}, //phyinit_io_write: 0x4124d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4124f, value : 32'h0}, //phyinit_io_write: 0x4124e, 0x4248
                          '{ step_type : REG_WRITE, reg_addr : 32'h41250, value : 32'h88d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=17 OP=0xac CS=0xa at row addr=0x128
                          '{ step_type : REG_WRITE, reg_addr : 32'h41251, value : 32'h0}, //phyinit_io_write: 0x41250, 0x88d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41252, value : 32'h9648}, //phyinit_io_write: 0x41251, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41253, value : 32'h0}, //phyinit_io_write: 0x41252, 0x9648
                          '{ step_type : REG_WRITE, reg_addr : 32'h41254, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41255, value : 32'h2b000000}, //phyinit_io_write: 0x41254, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41256, value : 32'h0}, //phyinit_io_write: 0x41255, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41257, value : 32'h0}, //phyinit_io_write: 0x41256, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41258, value : 32'hca58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=20 OP=0x2 CS=0xf at row addr=0x12c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41259, value : 32'h0}, //phyinit_io_write: 0x41258, 0xca58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4125a, value : 32'hc108}, //phyinit_io_write: 0x41259, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4125b, value : 32'h0}, //phyinit_io_write: 0x4125a, 0xc108
                          '{ step_type : REG_WRITE, reg_addr : 32'h4125c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4125d, value : 32'h2b000000}, //phyinit_io_write: 0x4125c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4125e, value : 32'h0}, //phyinit_io_write: 0x4125d, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4125f, value : 32'h0}, //phyinit_io_write: 0x4125e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41260, value : 32'hcb58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=22 OP=0x0 CS=0xf at row addr=0x130
                          '{ step_type : REG_WRITE, reg_addr : 32'h41261, value : 32'h0}, //phyinit_io_write: 0x41260, 0xcb58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41262, value : 32'hc008}, //phyinit_io_write: 0x41261, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41263, value : 32'h0}, //phyinit_io_write: 0x41262, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41264, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41265, value : 32'h2b000000}, //phyinit_io_write: 0x41264, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41266, value : 32'h0}, //phyinit_io_write: 0x41265, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41267, value : 32'h0}, //phyinit_io_write: 0x41266, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41268, value : 32'hd4d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=41 OP=0x60 CS=0xf at row addr=0x134
                          '{ step_type : REG_WRITE, reg_addr : 32'h41269, value : 32'h0}, //phyinit_io_write: 0x41268, 0xd4d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4126a, value : 32'hf008}, //phyinit_io_write: 0x41269, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4126b, value : 32'h0}, //phyinit_io_write: 0x4126a, 0xf008
                          '{ step_type : REG_WRITE, reg_addr : 32'h4126c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4126d, value : 32'h2b000000}, //phyinit_io_write: 0x4126c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4126e, value : 32'h0}, //phyinit_io_write: 0x4126d, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4126f, value : 32'h0}, //phyinit_io_write: 0x4126e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41270, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=58 at row addr=0x138
                          '{ step_type : REG_WRITE, reg_addr : 32'h41271, value : 32'h0}, //phyinit_io_write: 0x41270, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41272, value : 32'h0}, //phyinit_io_write: 0x41271, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41273, value : 32'h0}, //phyinit_io_write: 0x41272, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41274, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x13a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41275, value : 32'h0}, //phyinit_io_write: 0x41274, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h41276, value : 32'h6808}, //phyinit_io_write: 0x41275, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41277, value : 32'h0}, //phyinit_io_write: 0x41276, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41278, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x13c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41279, value : 32'h0}, //phyinit_io_write: 0x41278, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h4127a, value : 32'ha808}, //phyinit_io_write: 0x41279, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4127b, value : 32'h0}, //phyinit_io_write: 0x4127a, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h4127c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4127d, value : 32'h2b000000}, //phyinit_io_write: 0x4127c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4127e, value : 32'h0}, //phyinit_io_write: 0x4127d, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4127f, value : 32'h0}, //phyinit_io_write: 0x4127e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41280, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x140
                          '{ step_type : REG_WRITE, reg_addr : 32'h41281, value : 32'h0}, //phyinit_io_write: 0x41280, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h41282, value : 32'h6808}, //phyinit_io_write: 0x41281, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41283, value : 32'h0}, //phyinit_io_write: 0x41282, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41284, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x142
                          '{ step_type : REG_WRITE, reg_addr : 32'h41285, value : 32'h0}, //phyinit_io_write: 0x41284, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h41286, value : 32'ha808}, //phyinit_io_write: 0x41285, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41287, value : 32'h0}, //phyinit_io_write: 0x41286, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41288, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41289, value : 32'h2b000000}, //phyinit_io_write: 0x41288, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4128a, value : 32'h0}, //phyinit_io_write: 0x41289, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4128b, value : 32'h0}, //phyinit_io_write: 0x4128a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4128c, value : 32'h4758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0x5 at row addr=0x146
                          '{ step_type : REG_WRITE, reg_addr : 32'h4128d, value : 32'h0}, //phyinit_io_write: 0x4128c, 0x4758
                          '{ step_type : REG_WRITE, reg_addr : 32'h4128e, value : 32'h6808}, //phyinit_io_write: 0x4128d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4128f, value : 32'h0}, //phyinit_io_write: 0x4128e, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41290, value : 32'h8758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0xa at row addr=0x148
                          '{ step_type : REG_WRITE, reg_addr : 32'h41291, value : 32'h0}, //phyinit_io_write: 0x41290, 0x8758
                          '{ step_type : REG_WRITE, reg_addr : 32'h41292, value : 32'ha808}, //phyinit_io_write: 0x41291, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41293, value : 32'h0}, //phyinit_io_write: 0x41292, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41294, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41295, value : 32'h2b000000}, //phyinit_io_write: 0x41294, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41296, value : 32'h0}, //phyinit_io_write: 0x41295, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41297, value : 32'h0}, //phyinit_io_write: 0x41296, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41298, value : 32'h47d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0x5 at row addr=0x14c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41299, value : 32'h0}, //phyinit_io_write: 0x41298, 0x47d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4129a, value : 32'h6808}, //phyinit_io_write: 0x41299, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4129b, value : 32'h0}, //phyinit_io_write: 0x4129a, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h4129c, value : 32'h87d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0xa at row addr=0x14e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4129d, value : 32'h0}, //phyinit_io_write: 0x4129c, 0x87d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4129e, value : 32'ha808}, //phyinit_io_write: 0x4129d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4129f, value : 32'h0}, //phyinit_io_write: 0x4129e, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a0, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a1, value : 32'h2b000000}, //phyinit_io_write: 0x412a0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a2, value : 32'h0}, //phyinit_io_write: 0x412a1, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a3, value : 32'h0}, //phyinit_io_write: 0x412a2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a4, value : 32'h4c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0x5 at row addr=0x152
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a5, value : 32'h0}, //phyinit_io_write: 0x412a4, 0x4c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a6, value : 32'h4008}, //phyinit_io_write: 0x412a5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a7, value : 32'h0}, //phyinit_io_write: 0x412a6, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a8, value : 32'h8c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0xa at row addr=0x154
                          '{ step_type : REG_WRITE, reg_addr : 32'h412a9, value : 32'h0}, //phyinit_io_write: 0x412a8, 0x8c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h412aa, value : 32'h8008}, //phyinit_io_write: 0x412a9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ab, value : 32'h0}, //phyinit_io_write: 0x412aa, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ac, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ad, value : 32'h2b000000}, //phyinit_io_write: 0x412ac, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ae, value : 32'h0}, //phyinit_io_write: 0x412ad, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h412af, value : 32'h0}, //phyinit_io_write: 0x412ae, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b0, value : 32'h4f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0x5 at row addr=0x158
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b1, value : 32'h0}, //phyinit_io_write: 0x412b0, 0x4f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b2, value : 32'h4008}, //phyinit_io_write: 0x412b1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b3, value : 32'h0}, //phyinit_io_write: 0x412b2, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b4, value : 32'h8f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0xa at row addr=0x15a
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b5, value : 32'h0}, //phyinit_io_write: 0x412b4, 0x8f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b6, value : 32'h8008}, //phyinit_io_write: 0x412b5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b7, value : 32'h0}, //phyinit_io_write: 0x412b6, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b8, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h412b9, value : 32'h2b000000}, //phyinit_io_write: 0x412b8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ba, value : 32'h0}, //phyinit_io_write: 0x412b9, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h412bb, value : 32'h0}, //phyinit_io_write: 0x412ba, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412bc, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x15e
                          '{ step_type : REG_WRITE, reg_addr : 32'h412bd, value : 32'h0}, //phyinit_io_write: 0x412bc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412be, value : 32'h0}, //phyinit_io_write: 0x412bd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412bf, value : 32'h0}, //phyinit_io_write: 0x412be, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c0, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x160
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c1, value : 32'h0}, //phyinit_io_write: 0x412c0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c2, value : 32'h0}, //phyinit_io_write: 0x412c1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c3, value : 32'h0}, //phyinit_io_write: 0x412c2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c4, value : 32'h0}, //phyinit_io_write: 0x412c3, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c5, value : 32'h0}, //phyinit_io_write: 0x412c4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c6, value : 32'h0}, //phyinit_io_write: 0x412c5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c7, value : 32'h0}, //phyinit_io_write: 0x412c6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c8, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x164
                          '{ step_type : REG_WRITE, reg_addr : 32'h412c9, value : 32'h0}, //phyinit_io_write: 0x412c8, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ca, value : 32'h6808}, //phyinit_io_write: 0x412c9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412cb, value : 32'h0}, //phyinit_io_write: 0x412ca, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412cc, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x166
                          '{ step_type : REG_WRITE, reg_addr : 32'h412cd, value : 32'h0}, //phyinit_io_write: 0x412cc, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ce, value : 32'ha808}, //phyinit_io_write: 0x412cd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412cf, value : 32'h0}, //phyinit_io_write: 0x412ce, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d0, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d1, value : 32'h2b000000}, //phyinit_io_write: 0x412d0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d2, value : 32'h0}, //phyinit_io_write: 0x412d1, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d3, value : 32'h0}, //phyinit_io_write: 0x412d2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d4, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x16a
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d5, value : 32'h0}, //phyinit_io_write: 0x412d4, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d6, value : 32'h6808}, //phyinit_io_write: 0x412d5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d7, value : 32'h0}, //phyinit_io_write: 0x412d6, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d8, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x16c
                          '{ step_type : REG_WRITE, reg_addr : 32'h412d9, value : 32'h0}, //phyinit_io_write: 0x412d8, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h412da, value : 32'ha808}, //phyinit_io_write: 0x412d9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412db, value : 32'h0}, //phyinit_io_write: 0x412da, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412dc, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h412dd, value : 32'h2b000000}, //phyinit_io_write: 0x412dc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412de, value : 32'h0}, //phyinit_io_write: 0x412dd, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h412df, value : 32'h0}, //phyinit_io_write: 0x412de, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e0, value : 32'h4758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0x5 at row addr=0x170
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e1, value : 32'h0}, //phyinit_io_write: 0x412e0, 0x4758
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e2, value : 32'h6808}, //phyinit_io_write: 0x412e1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e3, value : 32'h0}, //phyinit_io_write: 0x412e2, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e4, value : 32'h8758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0xa at row addr=0x172
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e5, value : 32'h0}, //phyinit_io_write: 0x412e4, 0x8758
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e6, value : 32'ha808}, //phyinit_io_write: 0x412e5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e7, value : 32'h0}, //phyinit_io_write: 0x412e6, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e8, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h412e9, value : 32'h2b000000}, //phyinit_io_write: 0x412e8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ea, value : 32'h0}, //phyinit_io_write: 0x412e9, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h412eb, value : 32'h0}, //phyinit_io_write: 0x412ea, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ec, value : 32'h47d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0x5 at row addr=0x176
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ed, value : 32'h0}, //phyinit_io_write: 0x412ec, 0x47d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ee, value : 32'h6808}, //phyinit_io_write: 0x412ed, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ef, value : 32'h0}, //phyinit_io_write: 0x412ee, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f0, value : 32'h87d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0xa at row addr=0x178
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f1, value : 32'h0}, //phyinit_io_write: 0x412f0, 0x87d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f2, value : 32'ha808}, //phyinit_io_write: 0x412f1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f3, value : 32'h0}, //phyinit_io_write: 0x412f2, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f4, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f5, value : 32'h2b000000}, //phyinit_io_write: 0x412f4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f6, value : 32'h0}, //phyinit_io_write: 0x412f5, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f7, value : 32'h0}, //phyinit_io_write: 0x412f6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f8, value : 32'h4c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0x5 at row addr=0x17c
                          '{ step_type : REG_WRITE, reg_addr : 32'h412f9, value : 32'h0}, //phyinit_io_write: 0x412f8, 0x4c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h412fa, value : 32'h4008}, //phyinit_io_write: 0x412f9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412fb, value : 32'h0}, //phyinit_io_write: 0x412fa, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h412fc, value : 32'h8c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0xa at row addr=0x17e
                          '{ step_type : REG_WRITE, reg_addr : 32'h412fd, value : 32'h0}, //phyinit_io_write: 0x412fc, 0x8c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h412fe, value : 32'h8008}, //phyinit_io_write: 0x412fd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h412ff, value : 32'h0}, //phyinit_io_write: 0x412fe, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41300, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41301, value : 32'h2b000000}, //phyinit_io_write: 0x41300, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41302, value : 32'h0}, //phyinit_io_write: 0x41301, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41303, value : 32'h0}, //phyinit_io_write: 0x41302, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41304, value : 32'h4f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0x5 at row addr=0x182
                          '{ step_type : REG_WRITE, reg_addr : 32'h41305, value : 32'h0}, //phyinit_io_write: 0x41304, 0x4f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41306, value : 32'h4008}, //phyinit_io_write: 0x41305, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41307, value : 32'h0}, //phyinit_io_write: 0x41306, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41308, value : 32'h8f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0xa at row addr=0x184
                          '{ step_type : REG_WRITE, reg_addr : 32'h41309, value : 32'h0}, //phyinit_io_write: 0x41308, 0x8f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4130a, value : 32'h8008}, //phyinit_io_write: 0x41309, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4130b, value : 32'h0}, //phyinit_io_write: 0x4130a, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h4130c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4130d, value : 32'h2b000000}, //phyinit_io_write: 0x4130c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4130e, value : 32'h0}, //phyinit_io_write: 0x4130d, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4130f, value : 32'h0}, //phyinit_io_write: 0x4130e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41310, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x188
                          '{ step_type : REG_WRITE, reg_addr : 32'h41311, value : 32'h0}, //phyinit_io_write: 0x41310, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41312, value : 32'h0}, //phyinit_io_write: 0x41311, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41313, value : 32'h0}, //phyinit_io_write: 0x41312, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41314, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x18a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41315, value : 32'h0}, //phyinit_io_write: 0x41314, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41316, value : 32'h0}, //phyinit_io_write: 0x41315, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41317, value : 32'h0}, //phyinit_io_write: 0x41316, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41318, value : 32'h0}, //phyinit_io_write: 0x41317, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41319, value : 32'h0}, //phyinit_io_write: 0x41318, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4131a, value : 32'h0}, //phyinit_io_write: 0x41319, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4131b, value : 32'h0}, //phyinit_io_write: 0x4131a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h370145, value : 32'h1}, //[loadAcsmMRW] Pstate=3, Programming ACSMRptCntOverride to 1
                          '{ step_type : REG_WRITE, reg_addr : 32'h4131c, value : 32'hc9d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=19 OP=0x0 CS=0xf at row addr=0x18e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4131d, value : 32'h0}, //phyinit_io_write: 0x4131c, 0xc9d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4131e, value : 32'hc008}, //phyinit_io_write: 0x4131d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4131f, value : 32'h0}, //phyinit_io_write: 0x4131e, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41320, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41321, value : 32'h2b000000}, //phyinit_io_write: 0x41320, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41322, value : 32'h0}, //phyinit_io_write: 0x41321, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41323, value : 32'h0}, //phyinit_io_write: 0x41322, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41324, value : 32'hc958}, //[dwc_ddrphy_mr_inst] Storing MRW MA=18 OP=0x0 CS=0xf at row addr=0x192
                          '{ step_type : REG_WRITE, reg_addr : 32'h41325, value : 32'h0}, //phyinit_io_write: 0x41324, 0xc958
                          '{ step_type : REG_WRITE, reg_addr : 32'h41326, value : 32'hc008}, //phyinit_io_write: 0x41325, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41327, value : 32'h0}, //phyinit_io_write: 0x41326, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41328, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41329, value : 32'h2b000000}, //phyinit_io_write: 0x41328, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4132a, value : 32'h0}, //phyinit_io_write: 0x41329, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4132b, value : 32'h0}, //phyinit_io_write: 0x4132a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4132c, value : 32'hc0d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=1 OP=0x20 CS=0xf at row addr=0x196
                          '{ step_type : REG_WRITE, reg_addr : 32'h4132d, value : 32'h0}, //phyinit_io_write: 0x4132c, 0xc0d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4132e, value : 32'hd008}, //phyinit_io_write: 0x4132d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4132f, value : 32'h0}, //phyinit_io_write: 0x4132e, 0xd008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41330, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41331, value : 32'h2b000000}, //phyinit_io_write: 0x41330, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41332, value : 32'h0}, //phyinit_io_write: 0x41331, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41333, value : 32'h0}, //phyinit_io_write: 0x41332, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41334, value : 32'hc158}, //[dwc_ddrphy_mr_inst] Storing MRW MA=2 OP=0x22 CS=0xf at row addr=0x19a
                          '{ step_type : REG_WRITE, reg_addr : 32'h41335, value : 32'h0}, //phyinit_io_write: 0x41334, 0xc158
                          '{ step_type : REG_WRITE, reg_addr : 32'h41336, value : 32'hd108}, //phyinit_io_write: 0x41335, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41337, value : 32'h0}, //phyinit_io_write: 0x41336, 0xd108
                          '{ step_type : REG_WRITE, reg_addr : 32'h41338, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41339, value : 32'h2b000000}, //phyinit_io_write: 0x41338, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4133a, value : 32'h0}, //phyinit_io_write: 0x41339, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4133b, value : 32'h0}, //phyinit_io_write: 0x4133a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4133c, value : 32'hc1d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=3 OP=0xe CS=0xf at row addr=0x19e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4133d, value : 32'h0}, //phyinit_io_write: 0x4133c, 0xc1d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4133e, value : 32'hc708}, //phyinit_io_write: 0x4133d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4133f, value : 32'h0}, //phyinit_io_write: 0x4133e, 0xc708
                          '{ step_type : REG_WRITE, reg_addr : 32'h41340, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41341, value : 32'h2b000000}, //phyinit_io_write: 0x41340, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41342, value : 32'h0}, //phyinit_io_write: 0x41341, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41343, value : 32'h0}, //phyinit_io_write: 0x41342, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41344, value : 32'hc558}, //[dwc_ddrphy_mr_inst] Storing MRW MA=10 OP=0x54 CS=0xf at row addr=0x1a2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41345, value : 32'h0}, //phyinit_io_write: 0x41344, 0xc558
                          '{ step_type : REG_WRITE, reg_addr : 32'h41346, value : 32'hea08}, //phyinit_io_write: 0x41345, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41347, value : 32'h0}, //phyinit_io_write: 0x41346, 0xea08
                          '{ step_type : REG_WRITE, reg_addr : 32'h41348, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41349, value : 32'h2b000000}, //phyinit_io_write: 0x41348, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4134a, value : 32'h0}, //phyinit_io_write: 0x41349, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4134b, value : 32'h0}, //phyinit_io_write: 0x4134a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4134c, value : 32'hc5d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=11 OP=0x44 CS=0xf at row addr=0x1a6
                          '{ step_type : REG_WRITE, reg_addr : 32'h4134d, value : 32'h0}, //phyinit_io_write: 0x4134c, 0xc5d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4134e, value : 32'he208}, //phyinit_io_write: 0x4134d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4134f, value : 32'h0}, //phyinit_io_write: 0x4134e, 0xe208
                          '{ step_type : REG_WRITE, reg_addr : 32'h41350, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41351, value : 32'h2b000000}, //phyinit_io_write: 0x41350, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41352, value : 32'h0}, //phyinit_io_write: 0x41351, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41353, value : 32'h0}, //phyinit_io_write: 0x41352, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41354, value : 32'h48d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=17 OP=0x84 CS=0x5 at row addr=0x1aa
                          '{ step_type : REG_WRITE, reg_addr : 32'h41355, value : 32'h0}, //phyinit_io_write: 0x41354, 0x48d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41356, value : 32'h4248}, //phyinit_io_write: 0x41355, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41357, value : 32'h0}, //phyinit_io_write: 0x41356, 0x4248
                          '{ step_type : REG_WRITE, reg_addr : 32'h41358, value : 32'h88d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=17 OP=0xac CS=0xa at row addr=0x1ac
                          '{ step_type : REG_WRITE, reg_addr : 32'h41359, value : 32'h0}, //phyinit_io_write: 0x41358, 0x88d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h4135a, value : 32'h9648}, //phyinit_io_write: 0x41359, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4135b, value : 32'h0}, //phyinit_io_write: 0x4135a, 0x9648
                          '{ step_type : REG_WRITE, reg_addr : 32'h4135c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4135d, value : 32'h2b000000}, //phyinit_io_write: 0x4135c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4135e, value : 32'h0}, //phyinit_io_write: 0x4135d, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4135f, value : 32'h0}, //phyinit_io_write: 0x4135e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41360, value : 32'hca58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=20 OP=0x2 CS=0xf at row addr=0x1b0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41361, value : 32'h0}, //phyinit_io_write: 0x41360, 0xca58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41362, value : 32'hc108}, //phyinit_io_write: 0x41361, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41363, value : 32'h0}, //phyinit_io_write: 0x41362, 0xc108
                          '{ step_type : REG_WRITE, reg_addr : 32'h41364, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41365, value : 32'h2b000000}, //phyinit_io_write: 0x41364, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41366, value : 32'h0}, //phyinit_io_write: 0x41365, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41367, value : 32'h0}, //phyinit_io_write: 0x41366, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41368, value : 32'hcb58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=22 OP=0x0 CS=0xf at row addr=0x1b4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41369, value : 32'h0}, //phyinit_io_write: 0x41368, 0xcb58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4136a, value : 32'hc008}, //phyinit_io_write: 0x41369, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4136b, value : 32'h0}, //phyinit_io_write: 0x4136a, 0xc008
                          '{ step_type : REG_WRITE, reg_addr : 32'h4136c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4136d, value : 32'h2b000000}, //phyinit_io_write: 0x4136c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4136e, value : 32'h0}, //phyinit_io_write: 0x4136d, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4136f, value : 32'h0}, //phyinit_io_write: 0x4136e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41370, value : 32'hd4d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=41 OP=0x60 CS=0xf at row addr=0x1b8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41371, value : 32'h0}, //phyinit_io_write: 0x41370, 0xd4d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h41372, value : 32'hf008}, //phyinit_io_write: 0x41371, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41373, value : 32'h0}, //phyinit_io_write: 0x41372, 0xf008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41374, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41375, value : 32'h2b000000}, //phyinit_io_write: 0x41374, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41376, value : 32'h0}, //phyinit_io_write: 0x41375, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41377, value : 32'h0}, //phyinit_io_write: 0x41376, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41378, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=58 at row addr=0x1bc
                          '{ step_type : REG_WRITE, reg_addr : 32'h41379, value : 32'h0}, //phyinit_io_write: 0x41378, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4137a, value : 32'h0}, //phyinit_io_write: 0x41379, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4137b, value : 32'h0}, //phyinit_io_write: 0x4137a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4137c, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x1be
                          '{ step_type : REG_WRITE, reg_addr : 32'h4137d, value : 32'h0}, //phyinit_io_write: 0x4137c, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h4137e, value : 32'h6808}, //phyinit_io_write: 0x4137d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4137f, value : 32'h0}, //phyinit_io_write: 0x4137e, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41380, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x1c0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41381, value : 32'h0}, //phyinit_io_write: 0x41380, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h41382, value : 32'ha808}, //phyinit_io_write: 0x41381, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41383, value : 32'h0}, //phyinit_io_write: 0x41382, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41384, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41385, value : 32'h2b000000}, //phyinit_io_write: 0x41384, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41386, value : 32'h0}, //phyinit_io_write: 0x41385, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41387, value : 32'h0}, //phyinit_io_write: 0x41386, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41388, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x1c4
                          '{ step_type : REG_WRITE, reg_addr : 32'h41389, value : 32'h0}, //phyinit_io_write: 0x41388, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h4138a, value : 32'h6808}, //phyinit_io_write: 0x41389, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4138b, value : 32'h0}, //phyinit_io_write: 0x4138a, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h4138c, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x1c6
                          '{ step_type : REG_WRITE, reg_addr : 32'h4138d, value : 32'h0}, //phyinit_io_write: 0x4138c, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h4138e, value : 32'ha808}, //phyinit_io_write: 0x4138d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4138f, value : 32'h0}, //phyinit_io_write: 0x4138e, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41390, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41391, value : 32'h2b000000}, //phyinit_io_write: 0x41390, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41392, value : 32'h0}, //phyinit_io_write: 0x41391, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41393, value : 32'h0}, //phyinit_io_write: 0x41392, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41394, value : 32'h4758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0x5 at row addr=0x1ca
                          '{ step_type : REG_WRITE, reg_addr : 32'h41395, value : 32'h0}, //phyinit_io_write: 0x41394, 0x4758
                          '{ step_type : REG_WRITE, reg_addr : 32'h41396, value : 32'h6808}, //phyinit_io_write: 0x41395, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41397, value : 32'h0}, //phyinit_io_write: 0x41396, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h41398, value : 32'h8758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0xa at row addr=0x1cc
                          '{ step_type : REG_WRITE, reg_addr : 32'h41399, value : 32'h0}, //phyinit_io_write: 0x41398, 0x8758
                          '{ step_type : REG_WRITE, reg_addr : 32'h4139a, value : 32'ha808}, //phyinit_io_write: 0x41399, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4139b, value : 32'h0}, //phyinit_io_write: 0x4139a, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h4139c, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h4139d, value : 32'h2b000000}, //phyinit_io_write: 0x4139c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4139e, value : 32'h0}, //phyinit_io_write: 0x4139d, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4139f, value : 32'h0}, //phyinit_io_write: 0x4139e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a0, value : 32'h47d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0x5 at row addr=0x1d0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a1, value : 32'h0}, //phyinit_io_write: 0x413a0, 0x47d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a2, value : 32'h6808}, //phyinit_io_write: 0x413a1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a3, value : 32'h0}, //phyinit_io_write: 0x413a2, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a4, value : 32'h87d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0xa at row addr=0x1d2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a5, value : 32'h0}, //phyinit_io_write: 0x413a4, 0x87d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a6, value : 32'ha808}, //phyinit_io_write: 0x413a5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a7, value : 32'h0}, //phyinit_io_write: 0x413a6, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a8, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413a9, value : 32'h2b000000}, //phyinit_io_write: 0x413a8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413aa, value : 32'h0}, //phyinit_io_write: 0x413a9, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ab, value : 32'h0}, //phyinit_io_write: 0x413aa, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ac, value : 32'h4c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0x5 at row addr=0x1d6
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ad, value : 32'h0}, //phyinit_io_write: 0x413ac, 0x4c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ae, value : 32'h4008}, //phyinit_io_write: 0x413ad, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413af, value : 32'h0}, //phyinit_io_write: 0x413ae, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b0, value : 32'h8c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0xa at row addr=0x1d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b1, value : 32'h0}, //phyinit_io_write: 0x413b0, 0x8c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b2, value : 32'h8008}, //phyinit_io_write: 0x413b1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b3, value : 32'h0}, //phyinit_io_write: 0x413b2, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b4, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b5, value : 32'h2b000000}, //phyinit_io_write: 0x413b4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b6, value : 32'h0}, //phyinit_io_write: 0x413b5, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b7, value : 32'h0}, //phyinit_io_write: 0x413b6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b8, value : 32'h4f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0x5 at row addr=0x1dc
                          '{ step_type : REG_WRITE, reg_addr : 32'h413b9, value : 32'h0}, //phyinit_io_write: 0x413b8, 0x4f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ba, value : 32'h4008}, //phyinit_io_write: 0x413b9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413bb, value : 32'h0}, //phyinit_io_write: 0x413ba, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h413bc, value : 32'h8f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0xa at row addr=0x1de
                          '{ step_type : REG_WRITE, reg_addr : 32'h413bd, value : 32'h0}, //phyinit_io_write: 0x413bc, 0x8f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h413be, value : 32'h8008}, //phyinit_io_write: 0x413bd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413bf, value : 32'h0}, //phyinit_io_write: 0x413be, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c0, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c1, value : 32'h2b000000}, //phyinit_io_write: 0x413c0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c2, value : 32'h0}, //phyinit_io_write: 0x413c1, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c3, value : 32'h0}, //phyinit_io_write: 0x413c2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c4, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x1e2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c5, value : 32'h0}, //phyinit_io_write: 0x413c4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c6, value : 32'h0}, //phyinit_io_write: 0x413c5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c7, value : 32'h0}, //phyinit_io_write: 0x413c6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c8, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x1e4
                          '{ step_type : REG_WRITE, reg_addr : 32'h413c9, value : 32'h0}, //phyinit_io_write: 0x413c8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ca, value : 32'h0}, //phyinit_io_write: 0x413c9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413cb, value : 32'h0}, //phyinit_io_write: 0x413ca, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413cc, value : 32'h0}, //phyinit_io_write: 0x413cb, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413cd, value : 32'h0}, //phyinit_io_write: 0x413cc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ce, value : 32'h0}, //phyinit_io_write: 0x413cd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413cf, value : 32'h0}, //phyinit_io_write: 0x413ce, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d0, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x1e8
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d1, value : 32'h0}, //phyinit_io_write: 0x413d0, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d2, value : 32'h6808}, //phyinit_io_write: 0x413d1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d3, value : 32'h0}, //phyinit_io_write: 0x413d2, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d4, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x1ea
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d5, value : 32'h0}, //phyinit_io_write: 0x413d4, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d6, value : 32'ha808}, //phyinit_io_write: 0x413d5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d7, value : 32'h0}, //phyinit_io_write: 0x413d6, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d8, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413d9, value : 32'h2b000000}, //phyinit_io_write: 0x413d8, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413da, value : 32'h0}, //phyinit_io_write: 0x413d9, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h413db, value : 32'h0}, //phyinit_io_write: 0x413da, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413dc, value : 32'h4658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0x5 at row addr=0x1ee
                          '{ step_type : REG_WRITE, reg_addr : 32'h413dd, value : 32'h0}, //phyinit_io_write: 0x413dc, 0x4658
                          '{ step_type : REG_WRITE, reg_addr : 32'h413de, value : 32'h6808}, //phyinit_io_write: 0x413dd, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413df, value : 32'h0}, //phyinit_io_write: 0x413de, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e0, value : 32'h8658}, //[dwc_ddrphy_mr_inst] Storing MRW MA=12 OP=0x50 CS=0xa at row addr=0x1f0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e1, value : 32'h0}, //phyinit_io_write: 0x413e0, 0x8658
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e2, value : 32'ha808}, //phyinit_io_write: 0x413e1, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e3, value : 32'h0}, //phyinit_io_write: 0x413e2, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e4, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e5, value : 32'h2b000000}, //phyinit_io_write: 0x413e4, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e6, value : 32'h0}, //phyinit_io_write: 0x413e5, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e7, value : 32'h0}, //phyinit_io_write: 0x413e6, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e8, value : 32'h4758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0x5 at row addr=0x1f4
                          '{ step_type : REG_WRITE, reg_addr : 32'h413e9, value : 32'h0}, //phyinit_io_write: 0x413e8, 0x4758
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ea, value : 32'h6808}, //phyinit_io_write: 0x413e9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413eb, value : 32'h0}, //phyinit_io_write: 0x413ea, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ec, value : 32'h8758}, //[dwc_ddrphy_mr_inst] Storing MRW MA=14 OP=0x50 CS=0xa at row addr=0x1f6
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ed, value : 32'h0}, //phyinit_io_write: 0x413ec, 0x8758
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ee, value : 32'ha808}, //phyinit_io_write: 0x413ed, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ef, value : 32'h0}, //phyinit_io_write: 0x413ee, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f0, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f1, value : 32'h2b000000}, //phyinit_io_write: 0x413f0, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f2, value : 32'h0}, //phyinit_io_write: 0x413f1, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f3, value : 32'h0}, //phyinit_io_write: 0x413f2, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f4, value : 32'h47d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0x5 at row addr=0x1fa
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f5, value : 32'h0}, //phyinit_io_write: 0x413f4, 0x47d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f6, value : 32'h6808}, //phyinit_io_write: 0x413f5, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f7, value : 32'h0}, //phyinit_io_write: 0x413f6, 0x6808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f8, value : 32'h87d8}, //[dwc_ddrphy_mr_inst] Storing MRW MA=15 OP=0x50 CS=0xa at row addr=0x1fc
                          '{ step_type : REG_WRITE, reg_addr : 32'h413f9, value : 32'h0}, //phyinit_io_write: 0x413f8, 0x87d8
                          '{ step_type : REG_WRITE, reg_addr : 32'h413fa, value : 32'ha808}, //phyinit_io_write: 0x413f9, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413fb, value : 32'h0}, //phyinit_io_write: 0x413fa, 0xa808
                          '{ step_type : REG_WRITE, reg_addr : 32'h413fc, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h413fd, value : 32'h2b000000}, //phyinit_io_write: 0x413fc, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h413fe, value : 32'h0}, //phyinit_io_write: 0x413fd, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h413ff, value : 32'h0}, //phyinit_io_write: 0x413fe, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41400, value : 32'h4c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0x5 at row addr=0x200
                          '{ step_type : REG_WRITE, reg_addr : 32'h41401, value : 32'h0}, //phyinit_io_write: 0x41400, 0x4c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41402, value : 32'h4008}, //phyinit_io_write: 0x41401, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41403, value : 32'h0}, //phyinit_io_write: 0x41402, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41404, value : 32'h8c58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=24 OP=0x0 CS=0xa at row addr=0x202
                          '{ step_type : REG_WRITE, reg_addr : 32'h41405, value : 32'h0}, //phyinit_io_write: 0x41404, 0x8c58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41406, value : 32'h8008}, //phyinit_io_write: 0x41405, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41407, value : 32'h0}, //phyinit_io_write: 0x41406, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41408, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41409, value : 32'h2b000000}, //phyinit_io_write: 0x41408, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4140a, value : 32'h0}, //phyinit_io_write: 0x41409, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h4140b, value : 32'h0}, //phyinit_io_write: 0x4140a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4140c, value : 32'h4f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0x5 at row addr=0x206
                          '{ step_type : REG_WRITE, reg_addr : 32'h4140d, value : 32'h0}, //phyinit_io_write: 0x4140c, 0x4f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h4140e, value : 32'h4008}, //phyinit_io_write: 0x4140d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4140f, value : 32'h0}, //phyinit_io_write: 0x4140e, 0x4008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41410, value : 32'h8f58}, //[dwc_ddrphy_mr_inst] Storing MRW MA=30 OP=0x0 CS=0xa at row addr=0x208
                          '{ step_type : REG_WRITE, reg_addr : 32'h41411, value : 32'h0}, //phyinit_io_write: 0x41410, 0x8f58
                          '{ step_type : REG_WRITE, reg_addr : 32'h41412, value : 32'h8008}, //phyinit_io_write: 0x41411, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41413, value : 32'h0}, //phyinit_io_write: 0x41412, 0x8008
                          '{ step_type : REG_WRITE, reg_addr : 32'h41414, value : 32'h0}, //[dwc_ddrphy_mr_inst] dly = 5 cnt = 2
                          '{ step_type : REG_WRITE, reg_addr : 32'h41415, value : 32'h2b000000}, //phyinit_io_write: 0x41414, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41416, value : 32'h0}, //phyinit_io_write: 0x41415, 0x2b000000
                          '{ step_type : REG_WRITE, reg_addr : 32'h41417, value : 32'h0}, //phyinit_io_write: 0x41416, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41418, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x20c
                          '{ step_type : REG_WRITE, reg_addr : 32'h41419, value : 32'h0}, //phyinit_io_write: 0x41418, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4141a, value : 32'h0}, //phyinit_io_write: 0x41419, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4141b, value : 32'h0}, //phyinit_io_write: 0x4141a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4141c, value : 32'h0}, //[dwc_ddrphy_mr_clear] Reserving space for MRW MA=69 at row addr=0x20e
                          '{ step_type : REG_WRITE, reg_addr : 32'h4141d, value : 32'h0}, //phyinit_io_write: 0x4141c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4141e, value : 32'h0}, //phyinit_io_write: 0x4141d, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h4141f, value : 32'h0}, //phyinit_io_write: 0x4141e, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41420, value : 32'h0}, //phyinit_io_write: 0x4141f, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41421, value : 32'h0}, //phyinit_io_write: 0x41420, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41422, value : 32'h0}, //phyinit_io_write: 0x41421, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h41423, value : 32'h0}, //phyinit_io_write: 0x41422, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hd00e7, value : 32'h400}, //[loadAcsmMRW] End of loadAcsmMRW() inPsLoop=0
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0001, value : 32'h5821}, //phyinit_io_write: 0xd00e7, 0x400
                          '{ step_type : REG_WRITE, reg_addr : 32'h9070c, value : 32'h0}, //phyinit_io_write: 0xc0001, 0x5821
                          '{ step_type : REG_WRITE, reg_addr : 32'h9070d, value : 32'hfe}, //phyinit_io_write: 0x9070c, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h9070e, value : 32'hffff}, //phyinit_io_write: 0x9070d, 0xfe
                          '{ step_type : REG_WRITE, reg_addr : 32'h9070f, value : 32'hf040}, //phyinit_io_write: 0x9070e, 0xffff
                          '{ step_type : REG_WRITE, reg_addr : 32'h90710, value : 32'hf040}, //phyinit_io_write: 0x9070f, 0xf040
                          '{ step_type : REG_WRITE, reg_addr : 32'h90711, value : 32'h0}, //phyinit_io_write: 0x90710, 0xf040
                          '{ step_type : REG_WRITE, reg_addr : 32'h90712, value : 32'hffff}, //phyinit_io_write: 0x90711, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90713, value : 32'h0}, //phyinit_io_write: 0x90712, 0xffff
                          '{ step_type : REG_WRITE, reg_addr : 32'h90714, value : 32'h0}, //phyinit_io_write: 0x90713, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90715, value : 32'h0}, //phyinit_io_write: 0x90714, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90716, value : 32'h0}, //phyinit_io_write: 0x90715, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90717, value : 32'h0}, //phyinit_io_write: 0x90716, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90718, value : 32'h0}, //phyinit_io_write: 0x90717, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h90719, value : 32'h0}, //phyinit_io_write: 0x90718, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h9071a, value : 32'h0}, //phyinit_io_write: 0x90719, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h9071b, value : 32'h0}, //phyinit_io_write: 0x9071a, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h700f0, value : 32'hb6d}, //phyinit_io_write: 0x9071b, 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h7007e, value : 32'hc3}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programing Training Hardware Registers for mission mode retraining
                          '{ step_type : REG_WRITE, reg_addr : 32'h701ef, value : 32'h7fff}, //phyinit_io_write: 0x7007e, 0xc3
                          '{ step_type : REG_WRITE, reg_addr : 32'h300a6, value : 32'h1}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming AC0 ForceClkDisable to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h310a6, value : 32'h1}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming AC1 ForceClkDisable to 0x1
                          '{ step_type : REG_WRITE, reg_addr : 32'h701a8, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming PPGC ACSMParityInvert = 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70128, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming PPGC ACSMCkeControl = 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70131, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming PPGC ACSMInfiniteOLRC = 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70132, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming PPGC ACSMDefaultAddr = 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70133, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming PPGC ACSMDefaultCs = 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70134, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming PPGC ACSMStaticCtrl = 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70142, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming PPGC ACSMLowSpeedClockEnable = 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'h70144, value : 32'h0}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Programming PPGC ACSMLowSpeedClockDelay = 0x0
                          '{ step_type : REG_WRITE, reg_addr : 32'hc0080, value : 32'h6}, //[dwc_ddrphy_phyinit_I_loadPIEImage] Disabling Ucclk (PMU)
                          '{ step_type : REG_WRITE, reg_addr : 32'hd0000, value : 32'h1} //[dwc_ddrphy_phyinit_I_loadPIEImage] Isolate the APB access from the internal CSRs by setting the MicroContMuxSel CSR to 1.
//[dwc_ddrphy_phyinit_MicroContMuxSel_write32] phyinit_io_write to csr MicroContMuxSel: 0xd0000, 0x1
//[dwc_ddrphy_phyinit_I_loadPIEImage] End of dwc_ddrphy_phyinit_I_loadPIEImage()
//[dwc_ddrphy_phyinit_userCustom_customPostTrain] End of dwc_ddrphy_phyinit_userCustom_customPostTrain()
   }
                  
// [dwc_ddrphy_phyinit_userCustom_J_enterMissionMode] Start of dwc_ddrphy_phyinit_userCustom_J_enterMissionMode()
// [dwc_ddrphy_phyinit_userCustom_J_enterMissionMode] End of dwc_ddrphy_phyinit_userCustom_J_enterMissionMode()
 
};
