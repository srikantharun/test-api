// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description:
// UVM Incrementors
// Pre-configured incrementors for testbench construction
// Owner: abond

// Package: axe_uvm_incrementor_pkg 
package axe_uvm_incrementor_pkg;
  
    `include "uvm_macros.svh"
  
    import uvm_pkg::*;
  
    `include "axe_uvm_incrementor.svh"
    `include "axe_uvm_bitwise_incrementor.svh"

endpackage : axe_uvm_incrementor_pkg
