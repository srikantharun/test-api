// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024



`ifndef GUARD__TREK_UVM_EVENTS__SV
`define GUARD__TREK_UVM_EVENTS__SV

// This class is used within UVM simulations.
//
// It contains a single class that is simply a wrapper around a uvm_event_pool.
// The unique "key" string for each event corresponds to a "testbench port".
// Each "testbench port" has a string "name" that's called its "tb_path".
//
// TrekSoc indicates that it has data for a particular port ready to be pulled
//   across by firing the associated event.
//
// User-defined sequences will typically call "ev = TrekUvmEvents::get( myPath );"
//   to get the event that they should block and wait for.
//
// The methods here are static and should only be accessed with the "::" syntax
//   as above.
//

class trek_uvm_events;

  static protected bit  m_end_of_test = 0;  // Flag, set to one at end of test
  static protected uvm_event_pool  m_event_pool;  // Singleton instance

  function new();
    uvm_report_fatal("trek_uvm_events",
      "This class should never be instanced. Access it via static methods.",
      /* UVM_NONE */, `__FILE__, `__LINE__);
  endfunction: new

  // Provide information about each event in the managed pool
  static function string info();
    string          key;
    uvm_event_pool  pool;

    pool = get_pool();

    $sformat(info, "%0d events in pool...\n", pool.num());
    if (pool.first(key)) begin: e1
      do begin: e2
        uvm_event e;
        e = pool.get(key);
        $sformat(info, {info, "   %03s %019s (%0d waiters)\n"},
          e.is_on() ? " ON" : "OFF", key,
          e.get_num_waiters());
      end while (pool.next(key));
    end
  endfunction

  // Indicate that values written into memory won't be destroyed due
  //   to other initialization activities.
  static function void do_backdoor_init();
    uvm_event e;
    e = get("_trek_backdoor_init");
    e.trigger();
  endfunction: do_backdoor_init

  // Trek calls this method to indicate that the test is done. No more
  //   data will be sent, and it's time to gracefully shut down.
  static function void set_end_of_test();
    string          key;
    uvm_event_pool  pool;

    pool = get_pool();

    m_end_of_test = 1;

    if (pool.first(key)) begin: e1
      do begin: e2     // Loop through all known
        uvm_event e;   //   events and trigger them.
        e = pool.get(key);
        e.trigger();
      end while (pool.next(key));
    end
  endfunction: set_end_of_test

  // Query if the test is done.
  static function bit end_of_test();
    return m_end_of_test;
  endfunction: end_of_test

  // Return a handle to the singleton instance of the pool. If the
  //   pool doesn't exist yet, then build it.
  static function uvm_event_pool get_pool();
    if (m_event_pool == null) begin: new_pool
      m_event_pool = new("TrekUvmEventPool");
    end
    return m_event_pool;
  endfunction: get_pool

  // Return a handle to the event that manages a specific tb_path.
  static function uvm_event get( string tb_path );
    uvm_event_pool pool;
    pool = get_pool();
    return pool.get( tb_path );
  endfunction: get

  // Reset the pool 
  static function void clear();
    string          key;
    uvm_event_pool  pool;

    pool = get_pool();

    if (pool.first(key)) begin: e1
      do begin: e2     // Loop through all known
        pool.delete(key);
      end while (pool.next(key));
    end
     
    m_end_of_test = 0;
  endfunction: clear
   
endclass: trek_uvm_events

`endif // GUARD__TREK_UVM_EVENTS__SV
