// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_h_south
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_h_south (
    input  wire                                    i_aic_0_aon_clk,
    input  wire                                    i_aic_0_aon_rst_n,
    input  wire                                    i_aic_0_clk,
    input  wire                                    i_aic_0_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_0_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_0_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_0_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_0_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_0_init_ht_axi_s_arlen,
    input  logic                                   i_aic_0_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_0_init_ht_axi_s_arprot,
    output logic                                   o_aic_0_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_0_init_ht_axi_s_arsize,
    input  logic                                   i_aic_0_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_0_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_0_init_ht_axi_s_rid,
    output logic                                   o_aic_0_init_ht_axi_s_rlast,
    input  logic                                   i_aic_0_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_0_init_ht_axi_s_rresp,
    output logic                                   o_aic_0_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_0_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_0_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_0_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_0_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_0_init_ht_axi_s_awlen,
    input  logic                                   i_aic_0_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_0_init_ht_axi_s_awprot,
    output logic                                   o_aic_0_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_0_init_ht_axi_s_awsize,
    input  logic                                   i_aic_0_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_0_init_ht_axi_s_bid,
    input  logic                                   i_aic_0_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_0_init_ht_axi_s_bresp,
    output logic                                   o_aic_0_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_0_init_ht_axi_s_wdata,
    input  logic                                   i_aic_0_init_ht_axi_s_wlast,
    output logic                                   o_aic_0_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_0_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_0_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_0_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_0_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_0_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_0_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_0_init_lt_axi_s_arlen,
    input  logic                                   i_aic_0_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_0_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_0_init_lt_axi_s_arqos,
    output logic                                   o_aic_0_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_0_init_lt_axi_s_arsize,
    input  logic                                   i_aic_0_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_0_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_0_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_0_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_0_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_0_init_lt_axi_s_awlen,
    input  logic                                   i_aic_0_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_0_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_0_init_lt_axi_s_awqos,
    output logic                                   o_aic_0_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_0_init_lt_axi_s_awsize,
    input  logic                                   i_aic_0_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_0_init_lt_axi_s_bid,
    input  logic                                   i_aic_0_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_0_init_lt_axi_s_bresp,
    output logic                                   o_aic_0_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_0_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_0_init_lt_axi_s_rid,
    output logic                                   o_aic_0_init_lt_axi_s_rlast,
    input  logic                                   i_aic_0_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_0_init_lt_axi_s_rresp,
    output logic                                   o_aic_0_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_0_init_lt_axi_s_wdata,
    input  logic                                   i_aic_0_init_lt_axi_s_wlast,
    output logic                                   o_aic_0_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_0_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_0_init_lt_axi_s_wvalid,
    output logic                                   o_aic_0_pwr_idle_val,
    output logic                                   o_aic_0_pwr_idle_ack,
    input  logic                                   i_aic_0_pwr_idle_req,
    input  wire                                    i_aic_0_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_0_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_0_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_0_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_0_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_0_targ_lt_axi_m_arlen,
    output logic                                   o_aic_0_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_0_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_0_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_0_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_0_targ_lt_axi_m_arsize,
    output logic                                   o_aic_0_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_0_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_0_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_0_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_0_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_0_targ_lt_axi_m_awlen,
    output logic                                   o_aic_0_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_0_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_0_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_0_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_0_targ_lt_axi_m_awsize,
    output logic                                   o_aic_0_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_0_targ_lt_axi_m_bid,
    output logic                                   o_aic_0_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_0_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_0_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_0_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_0_targ_lt_axi_m_rid,
    input  logic                                   i_aic_0_targ_lt_axi_m_rlast,
    output logic                                   o_aic_0_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_0_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_0_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_0_targ_lt_axi_m_wdata,
    output logic                                   o_aic_0_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_0_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_0_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_0_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_0_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_0_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_0_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_0_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_0_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_0_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_1_aon_clk,
    input  wire                                    i_aic_1_aon_rst_n,
    input  wire                                    i_aic_1_clk,
    input  wire                                    i_aic_1_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_1_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_1_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_1_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_1_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_1_init_ht_axi_s_arlen,
    input  logic                                   i_aic_1_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_1_init_ht_axi_s_arprot,
    output logic                                   o_aic_1_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_1_init_ht_axi_s_arsize,
    input  logic                                   i_aic_1_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_1_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_1_init_ht_axi_s_rid,
    output logic                                   o_aic_1_init_ht_axi_s_rlast,
    input  logic                                   i_aic_1_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_1_init_ht_axi_s_rresp,
    output logic                                   o_aic_1_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_1_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_1_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_1_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_1_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_1_init_ht_axi_s_awlen,
    input  logic                                   i_aic_1_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_1_init_ht_axi_s_awprot,
    output logic                                   o_aic_1_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_1_init_ht_axi_s_awsize,
    input  logic                                   i_aic_1_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_1_init_ht_axi_s_bid,
    input  logic                                   i_aic_1_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_1_init_ht_axi_s_bresp,
    output logic                                   o_aic_1_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_1_init_ht_axi_s_wdata,
    input  logic                                   i_aic_1_init_ht_axi_s_wlast,
    output logic                                   o_aic_1_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_1_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_1_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_1_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_1_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_1_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_1_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_1_init_lt_axi_s_arlen,
    input  logic                                   i_aic_1_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_1_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_1_init_lt_axi_s_arqos,
    output logic                                   o_aic_1_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_1_init_lt_axi_s_arsize,
    input  logic                                   i_aic_1_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_1_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_1_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_1_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_1_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_1_init_lt_axi_s_awlen,
    input  logic                                   i_aic_1_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_1_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_1_init_lt_axi_s_awqos,
    output logic                                   o_aic_1_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_1_init_lt_axi_s_awsize,
    input  logic                                   i_aic_1_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_1_init_lt_axi_s_bid,
    input  logic                                   i_aic_1_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_1_init_lt_axi_s_bresp,
    output logic                                   o_aic_1_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_1_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_1_init_lt_axi_s_rid,
    output logic                                   o_aic_1_init_lt_axi_s_rlast,
    input  logic                                   i_aic_1_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_1_init_lt_axi_s_rresp,
    output logic                                   o_aic_1_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_1_init_lt_axi_s_wdata,
    input  logic                                   i_aic_1_init_lt_axi_s_wlast,
    output logic                                   o_aic_1_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_1_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_1_init_lt_axi_s_wvalid,
    output logic                                   o_aic_1_pwr_idle_val,
    output logic                                   o_aic_1_pwr_idle_ack,
    input  logic                                   i_aic_1_pwr_idle_req,
    input  wire                                    i_aic_1_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_1_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_1_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_1_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_1_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_1_targ_lt_axi_m_arlen,
    output logic                                   o_aic_1_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_1_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_1_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_1_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_1_targ_lt_axi_m_arsize,
    output logic                                   o_aic_1_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_1_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_1_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_1_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_1_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_1_targ_lt_axi_m_awlen,
    output logic                                   o_aic_1_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_1_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_1_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_1_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_1_targ_lt_axi_m_awsize,
    output logic                                   o_aic_1_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_1_targ_lt_axi_m_bid,
    output logic                                   o_aic_1_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_1_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_1_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_1_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_1_targ_lt_axi_m_rid,
    input  logic                                   i_aic_1_targ_lt_axi_m_rlast,
    output logic                                   o_aic_1_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_1_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_1_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_1_targ_lt_axi_m_wdata,
    output logic                                   o_aic_1_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_1_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_1_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_1_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_1_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_1_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_1_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_1_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_1_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_1_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_2_aon_clk,
    input  wire                                    i_aic_2_aon_rst_n,
    input  wire                                    i_aic_2_clk,
    input  wire                                    i_aic_2_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_2_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_2_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_2_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_2_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_2_init_ht_axi_s_arlen,
    input  logic                                   i_aic_2_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_2_init_ht_axi_s_arprot,
    output logic                                   o_aic_2_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_2_init_ht_axi_s_arsize,
    input  logic                                   i_aic_2_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_2_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_2_init_ht_axi_s_rid,
    output logic                                   o_aic_2_init_ht_axi_s_rlast,
    input  logic                                   i_aic_2_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_2_init_ht_axi_s_rresp,
    output logic                                   o_aic_2_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_2_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_2_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_2_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_2_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_2_init_ht_axi_s_awlen,
    input  logic                                   i_aic_2_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_2_init_ht_axi_s_awprot,
    output logic                                   o_aic_2_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_2_init_ht_axi_s_awsize,
    input  logic                                   i_aic_2_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_2_init_ht_axi_s_bid,
    input  logic                                   i_aic_2_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_2_init_ht_axi_s_bresp,
    output logic                                   o_aic_2_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_2_init_ht_axi_s_wdata,
    input  logic                                   i_aic_2_init_ht_axi_s_wlast,
    output logic                                   o_aic_2_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_2_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_2_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_2_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_2_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_2_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_2_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_2_init_lt_axi_s_arlen,
    input  logic                                   i_aic_2_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_2_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_2_init_lt_axi_s_arqos,
    output logic                                   o_aic_2_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_2_init_lt_axi_s_arsize,
    input  logic                                   i_aic_2_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_2_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_2_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_2_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_2_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_2_init_lt_axi_s_awlen,
    input  logic                                   i_aic_2_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_2_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_2_init_lt_axi_s_awqos,
    output logic                                   o_aic_2_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_2_init_lt_axi_s_awsize,
    input  logic                                   i_aic_2_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_2_init_lt_axi_s_bid,
    input  logic                                   i_aic_2_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_2_init_lt_axi_s_bresp,
    output logic                                   o_aic_2_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_2_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_2_init_lt_axi_s_rid,
    output logic                                   o_aic_2_init_lt_axi_s_rlast,
    input  logic                                   i_aic_2_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_2_init_lt_axi_s_rresp,
    output logic                                   o_aic_2_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_2_init_lt_axi_s_wdata,
    input  logic                                   i_aic_2_init_lt_axi_s_wlast,
    output logic                                   o_aic_2_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_2_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_2_init_lt_axi_s_wvalid,
    output logic                                   o_aic_2_pwr_idle_val,
    output logic                                   o_aic_2_pwr_idle_ack,
    input  logic                                   i_aic_2_pwr_idle_req,
    input  wire                                    i_aic_2_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_2_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_2_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_2_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_2_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_2_targ_lt_axi_m_arlen,
    output logic                                   o_aic_2_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_2_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_2_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_2_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_2_targ_lt_axi_m_arsize,
    output logic                                   o_aic_2_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_2_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_2_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_2_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_2_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_2_targ_lt_axi_m_awlen,
    output logic                                   o_aic_2_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_2_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_2_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_2_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_2_targ_lt_axi_m_awsize,
    output logic                                   o_aic_2_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_2_targ_lt_axi_m_bid,
    output logic                                   o_aic_2_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_2_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_2_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_2_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_2_targ_lt_axi_m_rid,
    input  logic                                   i_aic_2_targ_lt_axi_m_rlast,
    output logic                                   o_aic_2_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_2_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_2_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_2_targ_lt_axi_m_wdata,
    output logic                                   o_aic_2_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_2_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_2_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_2_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_2_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_2_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_2_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_2_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_2_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_2_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_3_aon_clk,
    input  wire                                    i_aic_3_aon_rst_n,
    input  wire                                    i_aic_3_clk,
    input  wire                                    i_aic_3_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_3_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_3_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_3_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_3_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_3_init_ht_axi_s_arlen,
    input  logic                                   i_aic_3_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_3_init_ht_axi_s_arprot,
    output logic                                   o_aic_3_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_3_init_ht_axi_s_arsize,
    input  logic                                   i_aic_3_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_3_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_3_init_ht_axi_s_rid,
    output logic                                   o_aic_3_init_ht_axi_s_rlast,
    input  logic                                   i_aic_3_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_3_init_ht_axi_s_rresp,
    output logic                                   o_aic_3_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_3_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_3_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_3_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_3_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_3_init_ht_axi_s_awlen,
    input  logic                                   i_aic_3_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_3_init_ht_axi_s_awprot,
    output logic                                   o_aic_3_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_3_init_ht_axi_s_awsize,
    input  logic                                   i_aic_3_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_3_init_ht_axi_s_bid,
    input  logic                                   i_aic_3_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_3_init_ht_axi_s_bresp,
    output logic                                   o_aic_3_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_3_init_ht_axi_s_wdata,
    input  logic                                   i_aic_3_init_ht_axi_s_wlast,
    output logic                                   o_aic_3_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_3_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_3_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_3_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_3_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_3_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_3_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_3_init_lt_axi_s_arlen,
    input  logic                                   i_aic_3_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_3_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_3_init_lt_axi_s_arqos,
    output logic                                   o_aic_3_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_3_init_lt_axi_s_arsize,
    input  logic                                   i_aic_3_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_3_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_3_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_3_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_3_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_3_init_lt_axi_s_awlen,
    input  logic                                   i_aic_3_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_3_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_3_init_lt_axi_s_awqos,
    output logic                                   o_aic_3_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_3_init_lt_axi_s_awsize,
    input  logic                                   i_aic_3_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_3_init_lt_axi_s_bid,
    input  logic                                   i_aic_3_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_3_init_lt_axi_s_bresp,
    output logic                                   o_aic_3_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_3_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_3_init_lt_axi_s_rid,
    output logic                                   o_aic_3_init_lt_axi_s_rlast,
    input  logic                                   i_aic_3_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_3_init_lt_axi_s_rresp,
    output logic                                   o_aic_3_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_3_init_lt_axi_s_wdata,
    input  logic                                   i_aic_3_init_lt_axi_s_wlast,
    output logic                                   o_aic_3_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_3_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_3_init_lt_axi_s_wvalid,
    output logic                                   o_aic_3_pwr_idle_val,
    output logic                                   o_aic_3_pwr_idle_ack,
    input  logic                                   i_aic_3_pwr_idle_req,
    input  wire                                    i_aic_3_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_3_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_3_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_3_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_3_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_3_targ_lt_axi_m_arlen,
    output logic                                   o_aic_3_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_3_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_3_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_3_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_3_targ_lt_axi_m_arsize,
    output logic                                   o_aic_3_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_3_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_3_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_3_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_3_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_3_targ_lt_axi_m_awlen,
    output logic                                   o_aic_3_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_3_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_3_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_3_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_3_targ_lt_axi_m_awsize,
    output logic                                   o_aic_3_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_3_targ_lt_axi_m_bid,
    output logic                                   o_aic_3_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_3_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_3_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_3_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_3_targ_lt_axi_m_rid,
    input  logic                                   i_aic_3_targ_lt_axi_m_rlast,
    output logic                                   o_aic_3_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_3_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_3_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_3_targ_lt_axi_m_wdata,
    output logic                                   o_aic_3_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_3_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_3_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_3_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_3_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_3_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_3_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_3_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_3_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_3_targ_syscfg_apb_m_pwrite,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld,
    input  logic [182:0]                           i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld,
    output logic [182:0]                           o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld,
    output logic [182:0]                           o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data,
    output logic                                   o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head,
    input  logic                                   i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy,
    output logic                                   o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail,
    output logic                                   o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld,
    input  logic [182:0]                           i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head,
    output logic                                   o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld,
    input  wire                                    i_l2_0_aon_clk,
    input  wire                                    i_l2_0_aon_rst_n,
    input  wire                                    i_l2_0_clk,
    input  wire                                    i_l2_0_clken,
    output logic                                   o_l2_0_pwr_idle_val,
    output logic                                   o_l2_0_pwr_idle_ack,
    input  logic                                   i_l2_0_pwr_idle_req,
    input  wire                                    i_l2_0_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_0_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_0_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_0_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_0_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_0_targ_ht_axi_m_arlen,
    output logic                                   o_l2_0_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_0_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_0_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_0_targ_ht_axi_m_arsize,
    output logic                                   o_l2_0_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_0_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_0_targ_ht_axi_m_rid,
    input  logic                                   i_l2_0_targ_ht_axi_m_rlast,
    output logic                                   o_l2_0_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_0_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_0_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_0_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_0_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_0_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_0_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_0_targ_ht_axi_m_awlen,
    output logic                                   o_l2_0_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_0_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_0_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_0_targ_ht_axi_m_awsize,
    output logic                                   o_l2_0_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_0_targ_ht_axi_m_bid,
    output logic                                   o_l2_0_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_0_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_0_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_0_targ_ht_axi_m_wdata,
    output logic                                   o_l2_0_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_0_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_0_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_0_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_0_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_0_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_0_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_0_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_0_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_0_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_1_aon_clk,
    input  wire                                    i_l2_1_aon_rst_n,
    input  wire                                    i_l2_1_clk,
    input  wire                                    i_l2_1_clken,
    output logic                                   o_l2_1_pwr_idle_val,
    output logic                                   o_l2_1_pwr_idle_ack,
    input  logic                                   i_l2_1_pwr_idle_req,
    input  wire                                    i_l2_1_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_1_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_1_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_1_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_1_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_1_targ_ht_axi_m_arlen,
    output logic                                   o_l2_1_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_1_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_1_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_1_targ_ht_axi_m_arsize,
    output logic                                   o_l2_1_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_1_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_1_targ_ht_axi_m_rid,
    input  logic                                   i_l2_1_targ_ht_axi_m_rlast,
    output logic                                   o_l2_1_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_1_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_1_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_1_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_1_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_1_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_1_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_1_targ_ht_axi_m_awlen,
    output logic                                   o_l2_1_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_1_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_1_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_1_targ_ht_axi_m_awsize,
    output logic                                   o_l2_1_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_1_targ_ht_axi_m_bid,
    output logic                                   o_l2_1_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_1_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_1_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_1_targ_ht_axi_m_wdata,
    output logic                                   o_l2_1_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_1_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_1_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_1_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_1_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_1_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_1_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_1_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_1_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_1_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_2_aon_clk,
    input  wire                                    i_l2_2_aon_rst_n,
    input  wire                                    i_l2_2_clk,
    input  wire                                    i_l2_2_clken,
    output logic                                   o_l2_2_pwr_idle_val,
    output logic                                   o_l2_2_pwr_idle_ack,
    input  logic                                   i_l2_2_pwr_idle_req,
    input  wire                                    i_l2_2_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_2_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_2_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_2_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_2_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_2_targ_ht_axi_m_arlen,
    output logic                                   o_l2_2_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_2_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_2_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_2_targ_ht_axi_m_arsize,
    output logic                                   o_l2_2_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_2_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_2_targ_ht_axi_m_rid,
    input  logic                                   i_l2_2_targ_ht_axi_m_rlast,
    output logic                                   o_l2_2_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_2_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_2_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_2_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_2_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_2_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_2_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_2_targ_ht_axi_m_awlen,
    output logic                                   o_l2_2_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_2_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_2_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_2_targ_ht_axi_m_awsize,
    output logic                                   o_l2_2_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_2_targ_ht_axi_m_bid,
    output logic                                   o_l2_2_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_2_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_2_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_2_targ_ht_axi_m_wdata,
    output logic                                   o_l2_2_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_2_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_2_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_2_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_2_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_2_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_2_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_2_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_2_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_2_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_3_aon_clk,
    input  wire                                    i_l2_3_aon_rst_n,
    input  wire                                    i_l2_3_clk,
    input  wire                                    i_l2_3_clken,
    output logic                                   o_l2_3_pwr_idle_val,
    output logic                                   o_l2_3_pwr_idle_ack,
    input  logic                                   i_l2_3_pwr_idle_req,
    input  wire                                    i_l2_3_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_3_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_3_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_3_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_3_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_3_targ_ht_axi_m_arlen,
    output logic                                   o_l2_3_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_3_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_3_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_3_targ_ht_axi_m_arsize,
    output logic                                   o_l2_3_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_3_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_3_targ_ht_axi_m_rid,
    input  logic                                   i_l2_3_targ_ht_axi_m_rlast,
    output logic                                   o_l2_3_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_3_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_3_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_3_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_3_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_3_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_3_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_3_targ_ht_axi_m_awlen,
    output logic                                   o_l2_3_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_3_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_3_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_3_targ_ht_axi_m_awsize,
    output logic                                   o_l2_3_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_3_targ_ht_axi_m_bid,
    output logic                                   o_l2_3_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_3_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_3_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_3_targ_ht_axi_m_wdata,
    output logic                                   o_l2_3_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_3_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_3_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_3_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_3_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_3_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_3_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_3_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_3_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_3_targ_syscfg_apb_m_pwrite,
    input  logic                                   i_l2_addr_mode_port_b0,
    input  logic                                   i_l2_addr_mode_port_b1,
    input  logic                                   i_l2_intr_mode_port_b0,
    input  logic                                   i_l2_intr_mode_port_b1,
    input  logic                                   i_lpddr_graph_addr_mode_port_b0,
    input  logic                                   i_lpddr_graph_addr_mode_port_b1,
    input  logic                                   i_lpddr_graph_intr_mode_port_b0,
    input  logic                                   i_lpddr_graph_intr_mode_port_b1,
    input  logic                                   i_lpddr_ppp_addr_mode_port_b0,
    input  logic                                   i_lpddr_ppp_addr_mode_port_b1,
    input  logic                                   i_lpddr_ppp_intr_mode_port_b0,
    input  logic                                   i_lpddr_ppp_intr_mode_port_b1,
    input  wire                                    i_noc_clk,
    input  wire                                    i_noc_rst_n,
    input  logic                                   scan_en
);

    // Automated Address MSB fix: extra nets declaration
    logic[40:0] aic_0_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] aic_0_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_0_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] aic_0_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_0_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] aic_0_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] aic_1_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] aic_1_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_1_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] aic_1_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_1_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] aic_1_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] aic_2_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] aic_2_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_2_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] aic_2_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_2_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] aic_2_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] aic_3_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] aic_3_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_3_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] aic_3_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_3_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] aic_3_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] l2_0_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] l2_0_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] l2_1_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] l2_1_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] l2_2_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] l2_2_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] l2_3_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] l2_3_targ_ht_axi_m_awaddr_msb_fixed;

    // Automated Address MSB fix: Initiator-side assignments to extend addresses by 1 bit
    noc_common_addr_msb_setter u_addr_msb_fix_aic_0_init_ht (
        .i_axi_araddr_40b (i_aic_0_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (aic_0_init_ht_axi_s_araddr_msb_fixed)
    );
    assign aic_0_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_aic_0_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_0_init_lt (
        .i_axi_araddr_40b (i_aic_0_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (aic_0_init_lt_axi_s_araddr_msb_fixed)
    );
    assign aic_0_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_aic_0_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_1_init_ht (
        .i_axi_araddr_40b (i_aic_1_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (aic_1_init_ht_axi_s_araddr_msb_fixed)
    );
    assign aic_1_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_aic_1_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_1_init_lt (
        .i_axi_araddr_40b (i_aic_1_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (aic_1_init_lt_axi_s_araddr_msb_fixed)
    );
    assign aic_1_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_aic_1_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_2_init_ht (
        .i_axi_araddr_40b (i_aic_2_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (aic_2_init_ht_axi_s_araddr_msb_fixed)
    );
    assign aic_2_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_aic_2_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_2_init_lt (
        .i_axi_araddr_40b (i_aic_2_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (aic_2_init_lt_axi_s_araddr_msb_fixed)
    );
    assign aic_2_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_aic_2_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_3_init_ht (
        .i_axi_araddr_40b (i_aic_3_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (aic_3_init_ht_axi_s_araddr_msb_fixed)
    );
    assign aic_3_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_aic_3_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_3_init_lt (
        .i_axi_araddr_40b (i_aic_3_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (aic_3_init_lt_axi_s_araddr_msb_fixed)
    );
    assign aic_3_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_aic_3_init_lt_axi_s_awaddr};

    // Automated Address MSB fix: Target-side assignments to drop unused MSB
    assign o_aic_0_targ_lt_axi_m_araddr = aic_0_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_aic_0_targ_lt_axi_m_awaddr = aic_0_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_aic_1_targ_lt_axi_m_araddr = aic_1_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_aic_1_targ_lt_axi_m_awaddr = aic_1_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_aic_2_targ_lt_axi_m_araddr = aic_2_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_aic_2_targ_lt_axi_m_awaddr = aic_2_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_aic_3_targ_lt_axi_m_araddr = aic_3_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_aic_3_targ_lt_axi_m_awaddr = aic_3_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_l2_0_targ_ht_axi_m_araddr = l2_0_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_l2_0_targ_ht_axi_m_awaddr = l2_0_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_l2_1_targ_ht_axi_m_araddr = l2_1_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_l2_1_targ_ht_axi_m_awaddr = l2_1_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_l2_2_targ_ht_axi_m_araddr = l2_2_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_l2_2_targ_ht_axi_m_awaddr = l2_2_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_l2_3_targ_ht_axi_m_araddr = l2_3_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_l2_3_targ_ht_axi_m_awaddr = l2_3_targ_ht_axi_m_awaddr_msb_fixed[39:0];


    noc_art_h_south u_noc_art_h_south (
    .aic_0_aon_clk(i_aic_0_aon_clk),
    .aic_0_aon_rst_n(i_aic_0_aon_rst_n),
    .aic_0_clk(i_aic_0_clk),
    .aic_0_clken(i_aic_0_clken),
    .aic_0_init_ht_rd_Ar_Addr(aic_0_init_ht_axi_s_araddr_msb_fixed),
    .aic_0_init_ht_rd_Ar_Burst(i_aic_0_init_ht_axi_s_arburst),
    .aic_0_init_ht_rd_Ar_Cache(i_aic_0_init_ht_axi_s_arcache),
    .aic_0_init_ht_rd_Ar_Id(i_aic_0_init_ht_axi_s_arid),
    .aic_0_init_ht_rd_Ar_Len(i_aic_0_init_ht_axi_s_arlen),
    .aic_0_init_ht_rd_Ar_Lock(i_aic_0_init_ht_axi_s_arlock),
    .aic_0_init_ht_rd_Ar_Prot(i_aic_0_init_ht_axi_s_arprot),
    .aic_0_init_ht_rd_Ar_Ready(o_aic_0_init_ht_axi_s_arready),
    .aic_0_init_ht_rd_Ar_Size(i_aic_0_init_ht_axi_s_arsize),
    .aic_0_init_ht_rd_Ar_Valid(i_aic_0_init_ht_axi_s_arvalid),
    .aic_0_init_ht_rd_R_Data(o_aic_0_init_ht_axi_s_rdata),
    .aic_0_init_ht_rd_R_Id(o_aic_0_init_ht_axi_s_rid),
    .aic_0_init_ht_rd_R_Last(o_aic_0_init_ht_axi_s_rlast),
    .aic_0_init_ht_rd_R_Ready(i_aic_0_init_ht_axi_s_rready),
    .aic_0_init_ht_rd_R_Resp(o_aic_0_init_ht_axi_s_rresp),
    .aic_0_init_ht_rd_R_Valid(o_aic_0_init_ht_axi_s_rvalid),
    .aic_0_init_ht_wr_Aw_Addr(aic_0_init_ht_axi_s_awaddr_msb_fixed),
    .aic_0_init_ht_wr_Aw_Burst(i_aic_0_init_ht_axi_s_awburst),
    .aic_0_init_ht_wr_Aw_Cache(i_aic_0_init_ht_axi_s_awcache),
    .aic_0_init_ht_wr_Aw_Id(i_aic_0_init_ht_axi_s_awid),
    .aic_0_init_ht_wr_Aw_Len(i_aic_0_init_ht_axi_s_awlen),
    .aic_0_init_ht_wr_Aw_Lock(i_aic_0_init_ht_axi_s_awlock),
    .aic_0_init_ht_wr_Aw_Prot(i_aic_0_init_ht_axi_s_awprot),
    .aic_0_init_ht_wr_Aw_Ready(o_aic_0_init_ht_axi_s_awready),
    .aic_0_init_ht_wr_Aw_Size(i_aic_0_init_ht_axi_s_awsize),
    .aic_0_init_ht_wr_Aw_Valid(i_aic_0_init_ht_axi_s_awvalid),
    .aic_0_init_ht_wr_B_Id(o_aic_0_init_ht_axi_s_bid),
    .aic_0_init_ht_wr_B_Ready(i_aic_0_init_ht_axi_s_bready),
    .aic_0_init_ht_wr_B_Resp(o_aic_0_init_ht_axi_s_bresp),
    .aic_0_init_ht_wr_B_Valid(o_aic_0_init_ht_axi_s_bvalid),
    .aic_0_init_ht_wr_W_Data(i_aic_0_init_ht_axi_s_wdata),
    .aic_0_init_ht_wr_W_Last(i_aic_0_init_ht_axi_s_wlast),
    .aic_0_init_ht_wr_W_Ready(o_aic_0_init_ht_axi_s_wready),
    .aic_0_init_ht_wr_W_Strb(i_aic_0_init_ht_axi_s_wstrb),
    .aic_0_init_ht_wr_W_Valid(i_aic_0_init_ht_axi_s_wvalid),
    .aic_0_init_lt_Ar_Addr(aic_0_init_lt_axi_s_araddr_msb_fixed),
    .aic_0_init_lt_Ar_Burst(i_aic_0_init_lt_axi_s_arburst),
    .aic_0_init_lt_Ar_Cache(i_aic_0_init_lt_axi_s_arcache),
    .aic_0_init_lt_Ar_Id(i_aic_0_init_lt_axi_s_arid),
    .aic_0_init_lt_Ar_Len(i_aic_0_init_lt_axi_s_arlen),
    .aic_0_init_lt_Ar_Lock(i_aic_0_init_lt_axi_s_arlock),
    .aic_0_init_lt_Ar_Prot(i_aic_0_init_lt_axi_s_arprot),
    .aic_0_init_lt_Ar_Qos(i_aic_0_init_lt_axi_s_arqos),
    .aic_0_init_lt_Ar_Ready(o_aic_0_init_lt_axi_s_arready),
    .aic_0_init_lt_Ar_Size(i_aic_0_init_lt_axi_s_arsize),
    .aic_0_init_lt_Ar_Valid(i_aic_0_init_lt_axi_s_arvalid),
    .aic_0_init_lt_Aw_Addr(aic_0_init_lt_axi_s_awaddr_msb_fixed),
    .aic_0_init_lt_Aw_Burst(i_aic_0_init_lt_axi_s_awburst),
    .aic_0_init_lt_Aw_Cache(i_aic_0_init_lt_axi_s_awcache),
    .aic_0_init_lt_Aw_Id(i_aic_0_init_lt_axi_s_awid),
    .aic_0_init_lt_Aw_Len(i_aic_0_init_lt_axi_s_awlen),
    .aic_0_init_lt_Aw_Lock(i_aic_0_init_lt_axi_s_awlock),
    .aic_0_init_lt_Aw_Prot(i_aic_0_init_lt_axi_s_awprot),
    .aic_0_init_lt_Aw_Qos(i_aic_0_init_lt_axi_s_awqos),
    .aic_0_init_lt_Aw_Ready(o_aic_0_init_lt_axi_s_awready),
    .aic_0_init_lt_Aw_Size(i_aic_0_init_lt_axi_s_awsize),
    .aic_0_init_lt_Aw_Valid(i_aic_0_init_lt_axi_s_awvalid),
    .aic_0_init_lt_B_Id(o_aic_0_init_lt_axi_s_bid),
    .aic_0_init_lt_B_Ready(i_aic_0_init_lt_axi_s_bready),
    .aic_0_init_lt_B_Resp(o_aic_0_init_lt_axi_s_bresp),
    .aic_0_init_lt_B_Valid(o_aic_0_init_lt_axi_s_bvalid),
    .aic_0_init_lt_R_Data(o_aic_0_init_lt_axi_s_rdata),
    .aic_0_init_lt_R_Id(o_aic_0_init_lt_axi_s_rid),
    .aic_0_init_lt_R_Last(o_aic_0_init_lt_axi_s_rlast),
    .aic_0_init_lt_R_Ready(i_aic_0_init_lt_axi_s_rready),
    .aic_0_init_lt_R_Resp(o_aic_0_init_lt_axi_s_rresp),
    .aic_0_init_lt_R_Valid(o_aic_0_init_lt_axi_s_rvalid),
    .aic_0_init_lt_W_Data(i_aic_0_init_lt_axi_s_wdata),
    .aic_0_init_lt_W_Last(i_aic_0_init_lt_axi_s_wlast),
    .aic_0_init_lt_W_Ready(o_aic_0_init_lt_axi_s_wready),
    .aic_0_init_lt_W_Strb(i_aic_0_init_lt_axi_s_wstrb),
    .aic_0_init_lt_W_Valid(i_aic_0_init_lt_axi_s_wvalid),
    .aic_0_pwr_Idle(o_aic_0_pwr_idle_val),
    .aic_0_pwr_IdleAck(o_aic_0_pwr_idle_ack),
    .aic_0_pwr_IdleReq(i_aic_0_pwr_idle_req),
    .aic_0_rst_n(i_aic_0_rst_n),
    .aic_0_targ_lt_Ar_Addr(aic_0_targ_lt_axi_m_araddr_msb_fixed),
    .aic_0_targ_lt_Ar_Burst(o_aic_0_targ_lt_axi_m_arburst),
    .aic_0_targ_lt_Ar_Cache(o_aic_0_targ_lt_axi_m_arcache),
    .aic_0_targ_lt_Ar_Id(o_aic_0_targ_lt_axi_m_arid),
    .aic_0_targ_lt_Ar_Len(o_aic_0_targ_lt_axi_m_arlen),
    .aic_0_targ_lt_Ar_Lock(o_aic_0_targ_lt_axi_m_arlock),
    .aic_0_targ_lt_Ar_Prot(o_aic_0_targ_lt_axi_m_arprot),
    .aic_0_targ_lt_Ar_Qos(o_aic_0_targ_lt_axi_m_arqos),
    .aic_0_targ_lt_Ar_Ready(i_aic_0_targ_lt_axi_m_arready),
    .aic_0_targ_lt_Ar_Size(o_aic_0_targ_lt_axi_m_arsize),
    .aic_0_targ_lt_Ar_Valid(o_aic_0_targ_lt_axi_m_arvalid),
    .aic_0_targ_lt_Aw_Addr(aic_0_targ_lt_axi_m_awaddr_msb_fixed),
    .aic_0_targ_lt_Aw_Burst(o_aic_0_targ_lt_axi_m_awburst),
    .aic_0_targ_lt_Aw_Cache(o_aic_0_targ_lt_axi_m_awcache),
    .aic_0_targ_lt_Aw_Id(o_aic_0_targ_lt_axi_m_awid),
    .aic_0_targ_lt_Aw_Len(o_aic_0_targ_lt_axi_m_awlen),
    .aic_0_targ_lt_Aw_Lock(o_aic_0_targ_lt_axi_m_awlock),
    .aic_0_targ_lt_Aw_Prot(o_aic_0_targ_lt_axi_m_awprot),
    .aic_0_targ_lt_Aw_Qos(o_aic_0_targ_lt_axi_m_awqos),
    .aic_0_targ_lt_Aw_Ready(i_aic_0_targ_lt_axi_m_awready),
    .aic_0_targ_lt_Aw_Size(o_aic_0_targ_lt_axi_m_awsize),
    .aic_0_targ_lt_Aw_Valid(o_aic_0_targ_lt_axi_m_awvalid),
    .aic_0_targ_lt_B_Id(i_aic_0_targ_lt_axi_m_bid),
    .aic_0_targ_lt_B_Ready(o_aic_0_targ_lt_axi_m_bready),
    .aic_0_targ_lt_B_Resp(i_aic_0_targ_lt_axi_m_bresp),
    .aic_0_targ_lt_B_Valid(i_aic_0_targ_lt_axi_m_bvalid),
    .aic_0_targ_lt_R_Data(i_aic_0_targ_lt_axi_m_rdata),
    .aic_0_targ_lt_R_Id(i_aic_0_targ_lt_axi_m_rid),
    .aic_0_targ_lt_R_Last(i_aic_0_targ_lt_axi_m_rlast),
    .aic_0_targ_lt_R_Ready(o_aic_0_targ_lt_axi_m_rready),
    .aic_0_targ_lt_R_Resp(i_aic_0_targ_lt_axi_m_rresp),
    .aic_0_targ_lt_R_Valid(i_aic_0_targ_lt_axi_m_rvalid),
    .aic_0_targ_lt_W_Data(o_aic_0_targ_lt_axi_m_wdata),
    .aic_0_targ_lt_W_Last(o_aic_0_targ_lt_axi_m_wlast),
    .aic_0_targ_lt_W_Ready(i_aic_0_targ_lt_axi_m_wready),
    .aic_0_targ_lt_W_Strb(o_aic_0_targ_lt_axi_m_wstrb),
    .aic_0_targ_lt_W_Valid(o_aic_0_targ_lt_axi_m_wvalid),
    .aic_0_targ_syscfg_PAddr(o_aic_0_targ_syscfg_apb_m_paddr),
    .aic_0_targ_syscfg_PEnable(o_aic_0_targ_syscfg_apb_m_penable),
    .aic_0_targ_syscfg_PProt(o_aic_0_targ_syscfg_apb_m_pprot),
    .aic_0_targ_syscfg_PRData(i_aic_0_targ_syscfg_apb_m_prdata),
    .aic_0_targ_syscfg_PReady(i_aic_0_targ_syscfg_apb_m_pready),
    .aic_0_targ_syscfg_PSel(o_aic_0_targ_syscfg_apb_m_psel),
    .aic_0_targ_syscfg_PSlvErr(i_aic_0_targ_syscfg_apb_m_pslverr),
    .aic_0_targ_syscfg_PStrb(o_aic_0_targ_syscfg_apb_m_pstrb),
    .aic_0_targ_syscfg_PWData(o_aic_0_targ_syscfg_apb_m_pwdata),
    .aic_0_targ_syscfg_PWrite(o_aic_0_targ_syscfg_apb_m_pwrite),
    .aic_1_aon_clk(i_aic_1_aon_clk),
    .aic_1_aon_rst_n(i_aic_1_aon_rst_n),
    .aic_1_clk(i_aic_1_clk),
    .aic_1_clken(i_aic_1_clken),
    .aic_1_init_ht_rd_Ar_Addr(aic_1_init_ht_axi_s_araddr_msb_fixed),
    .aic_1_init_ht_rd_Ar_Burst(i_aic_1_init_ht_axi_s_arburst),
    .aic_1_init_ht_rd_Ar_Cache(i_aic_1_init_ht_axi_s_arcache),
    .aic_1_init_ht_rd_Ar_Id(i_aic_1_init_ht_axi_s_arid),
    .aic_1_init_ht_rd_Ar_Len(i_aic_1_init_ht_axi_s_arlen),
    .aic_1_init_ht_rd_Ar_Lock(i_aic_1_init_ht_axi_s_arlock),
    .aic_1_init_ht_rd_Ar_Prot(i_aic_1_init_ht_axi_s_arprot),
    .aic_1_init_ht_rd_Ar_Ready(o_aic_1_init_ht_axi_s_arready),
    .aic_1_init_ht_rd_Ar_Size(i_aic_1_init_ht_axi_s_arsize),
    .aic_1_init_ht_rd_Ar_Valid(i_aic_1_init_ht_axi_s_arvalid),
    .aic_1_init_ht_rd_R_Data(o_aic_1_init_ht_axi_s_rdata),
    .aic_1_init_ht_rd_R_Id(o_aic_1_init_ht_axi_s_rid),
    .aic_1_init_ht_rd_R_Last(o_aic_1_init_ht_axi_s_rlast),
    .aic_1_init_ht_rd_R_Ready(i_aic_1_init_ht_axi_s_rready),
    .aic_1_init_ht_rd_R_Resp(o_aic_1_init_ht_axi_s_rresp),
    .aic_1_init_ht_rd_R_Valid(o_aic_1_init_ht_axi_s_rvalid),
    .aic_1_init_ht_wr_Aw_Addr(aic_1_init_ht_axi_s_awaddr_msb_fixed),
    .aic_1_init_ht_wr_Aw_Burst(i_aic_1_init_ht_axi_s_awburst),
    .aic_1_init_ht_wr_Aw_Cache(i_aic_1_init_ht_axi_s_awcache),
    .aic_1_init_ht_wr_Aw_Id(i_aic_1_init_ht_axi_s_awid),
    .aic_1_init_ht_wr_Aw_Len(i_aic_1_init_ht_axi_s_awlen),
    .aic_1_init_ht_wr_Aw_Lock(i_aic_1_init_ht_axi_s_awlock),
    .aic_1_init_ht_wr_Aw_Prot(i_aic_1_init_ht_axi_s_awprot),
    .aic_1_init_ht_wr_Aw_Ready(o_aic_1_init_ht_axi_s_awready),
    .aic_1_init_ht_wr_Aw_Size(i_aic_1_init_ht_axi_s_awsize),
    .aic_1_init_ht_wr_Aw_Valid(i_aic_1_init_ht_axi_s_awvalid),
    .aic_1_init_ht_wr_B_Id(o_aic_1_init_ht_axi_s_bid),
    .aic_1_init_ht_wr_B_Ready(i_aic_1_init_ht_axi_s_bready),
    .aic_1_init_ht_wr_B_Resp(o_aic_1_init_ht_axi_s_bresp),
    .aic_1_init_ht_wr_B_Valid(o_aic_1_init_ht_axi_s_bvalid),
    .aic_1_init_ht_wr_W_Data(i_aic_1_init_ht_axi_s_wdata),
    .aic_1_init_ht_wr_W_Last(i_aic_1_init_ht_axi_s_wlast),
    .aic_1_init_ht_wr_W_Ready(o_aic_1_init_ht_axi_s_wready),
    .aic_1_init_ht_wr_W_Strb(i_aic_1_init_ht_axi_s_wstrb),
    .aic_1_init_ht_wr_W_Valid(i_aic_1_init_ht_axi_s_wvalid),
    .aic_1_init_lt_Ar_Addr(aic_1_init_lt_axi_s_araddr_msb_fixed),
    .aic_1_init_lt_Ar_Burst(i_aic_1_init_lt_axi_s_arburst),
    .aic_1_init_lt_Ar_Cache(i_aic_1_init_lt_axi_s_arcache),
    .aic_1_init_lt_Ar_Id(i_aic_1_init_lt_axi_s_arid),
    .aic_1_init_lt_Ar_Len(i_aic_1_init_lt_axi_s_arlen),
    .aic_1_init_lt_Ar_Lock(i_aic_1_init_lt_axi_s_arlock),
    .aic_1_init_lt_Ar_Prot(i_aic_1_init_lt_axi_s_arprot),
    .aic_1_init_lt_Ar_Qos(i_aic_1_init_lt_axi_s_arqos),
    .aic_1_init_lt_Ar_Ready(o_aic_1_init_lt_axi_s_arready),
    .aic_1_init_lt_Ar_Size(i_aic_1_init_lt_axi_s_arsize),
    .aic_1_init_lt_Ar_Valid(i_aic_1_init_lt_axi_s_arvalid),
    .aic_1_init_lt_Aw_Addr(aic_1_init_lt_axi_s_awaddr_msb_fixed),
    .aic_1_init_lt_Aw_Burst(i_aic_1_init_lt_axi_s_awburst),
    .aic_1_init_lt_Aw_Cache(i_aic_1_init_lt_axi_s_awcache),
    .aic_1_init_lt_Aw_Id(i_aic_1_init_lt_axi_s_awid),
    .aic_1_init_lt_Aw_Len(i_aic_1_init_lt_axi_s_awlen),
    .aic_1_init_lt_Aw_Lock(i_aic_1_init_lt_axi_s_awlock),
    .aic_1_init_lt_Aw_Prot(i_aic_1_init_lt_axi_s_awprot),
    .aic_1_init_lt_Aw_Qos(i_aic_1_init_lt_axi_s_awqos),
    .aic_1_init_lt_Aw_Ready(o_aic_1_init_lt_axi_s_awready),
    .aic_1_init_lt_Aw_Size(i_aic_1_init_lt_axi_s_awsize),
    .aic_1_init_lt_Aw_Valid(i_aic_1_init_lt_axi_s_awvalid),
    .aic_1_init_lt_B_Id(o_aic_1_init_lt_axi_s_bid),
    .aic_1_init_lt_B_Ready(i_aic_1_init_lt_axi_s_bready),
    .aic_1_init_lt_B_Resp(o_aic_1_init_lt_axi_s_bresp),
    .aic_1_init_lt_B_Valid(o_aic_1_init_lt_axi_s_bvalid),
    .aic_1_init_lt_R_Data(o_aic_1_init_lt_axi_s_rdata),
    .aic_1_init_lt_R_Id(o_aic_1_init_lt_axi_s_rid),
    .aic_1_init_lt_R_Last(o_aic_1_init_lt_axi_s_rlast),
    .aic_1_init_lt_R_Ready(i_aic_1_init_lt_axi_s_rready),
    .aic_1_init_lt_R_Resp(o_aic_1_init_lt_axi_s_rresp),
    .aic_1_init_lt_R_Valid(o_aic_1_init_lt_axi_s_rvalid),
    .aic_1_init_lt_W_Data(i_aic_1_init_lt_axi_s_wdata),
    .aic_1_init_lt_W_Last(i_aic_1_init_lt_axi_s_wlast),
    .aic_1_init_lt_W_Ready(o_aic_1_init_lt_axi_s_wready),
    .aic_1_init_lt_W_Strb(i_aic_1_init_lt_axi_s_wstrb),
    .aic_1_init_lt_W_Valid(i_aic_1_init_lt_axi_s_wvalid),
    .aic_1_pwr_Idle(o_aic_1_pwr_idle_val),
    .aic_1_pwr_IdleAck(o_aic_1_pwr_idle_ack),
    .aic_1_pwr_IdleReq(i_aic_1_pwr_idle_req),
    .aic_1_rst_n(i_aic_1_rst_n),
    .aic_1_targ_lt_Ar_Addr(aic_1_targ_lt_axi_m_araddr_msb_fixed),
    .aic_1_targ_lt_Ar_Burst(o_aic_1_targ_lt_axi_m_arburst),
    .aic_1_targ_lt_Ar_Cache(o_aic_1_targ_lt_axi_m_arcache),
    .aic_1_targ_lt_Ar_Id(o_aic_1_targ_lt_axi_m_arid),
    .aic_1_targ_lt_Ar_Len(o_aic_1_targ_lt_axi_m_arlen),
    .aic_1_targ_lt_Ar_Lock(o_aic_1_targ_lt_axi_m_arlock),
    .aic_1_targ_lt_Ar_Prot(o_aic_1_targ_lt_axi_m_arprot),
    .aic_1_targ_lt_Ar_Qos(o_aic_1_targ_lt_axi_m_arqos),
    .aic_1_targ_lt_Ar_Ready(i_aic_1_targ_lt_axi_m_arready),
    .aic_1_targ_lt_Ar_Size(o_aic_1_targ_lt_axi_m_arsize),
    .aic_1_targ_lt_Ar_Valid(o_aic_1_targ_lt_axi_m_arvalid),
    .aic_1_targ_lt_Aw_Addr(aic_1_targ_lt_axi_m_awaddr_msb_fixed),
    .aic_1_targ_lt_Aw_Burst(o_aic_1_targ_lt_axi_m_awburst),
    .aic_1_targ_lt_Aw_Cache(o_aic_1_targ_lt_axi_m_awcache),
    .aic_1_targ_lt_Aw_Id(o_aic_1_targ_lt_axi_m_awid),
    .aic_1_targ_lt_Aw_Len(o_aic_1_targ_lt_axi_m_awlen),
    .aic_1_targ_lt_Aw_Lock(o_aic_1_targ_lt_axi_m_awlock),
    .aic_1_targ_lt_Aw_Prot(o_aic_1_targ_lt_axi_m_awprot),
    .aic_1_targ_lt_Aw_Qos(o_aic_1_targ_lt_axi_m_awqos),
    .aic_1_targ_lt_Aw_Ready(i_aic_1_targ_lt_axi_m_awready),
    .aic_1_targ_lt_Aw_Size(o_aic_1_targ_lt_axi_m_awsize),
    .aic_1_targ_lt_Aw_Valid(o_aic_1_targ_lt_axi_m_awvalid),
    .aic_1_targ_lt_B_Id(i_aic_1_targ_lt_axi_m_bid),
    .aic_1_targ_lt_B_Ready(o_aic_1_targ_lt_axi_m_bready),
    .aic_1_targ_lt_B_Resp(i_aic_1_targ_lt_axi_m_bresp),
    .aic_1_targ_lt_B_Valid(i_aic_1_targ_lt_axi_m_bvalid),
    .aic_1_targ_lt_R_Data(i_aic_1_targ_lt_axi_m_rdata),
    .aic_1_targ_lt_R_Id(i_aic_1_targ_lt_axi_m_rid),
    .aic_1_targ_lt_R_Last(i_aic_1_targ_lt_axi_m_rlast),
    .aic_1_targ_lt_R_Ready(o_aic_1_targ_lt_axi_m_rready),
    .aic_1_targ_lt_R_Resp(i_aic_1_targ_lt_axi_m_rresp),
    .aic_1_targ_lt_R_Valid(i_aic_1_targ_lt_axi_m_rvalid),
    .aic_1_targ_lt_W_Data(o_aic_1_targ_lt_axi_m_wdata),
    .aic_1_targ_lt_W_Last(o_aic_1_targ_lt_axi_m_wlast),
    .aic_1_targ_lt_W_Ready(i_aic_1_targ_lt_axi_m_wready),
    .aic_1_targ_lt_W_Strb(o_aic_1_targ_lt_axi_m_wstrb),
    .aic_1_targ_lt_W_Valid(o_aic_1_targ_lt_axi_m_wvalid),
    .aic_1_targ_syscfg_PAddr(o_aic_1_targ_syscfg_apb_m_paddr),
    .aic_1_targ_syscfg_PEnable(o_aic_1_targ_syscfg_apb_m_penable),
    .aic_1_targ_syscfg_PProt(o_aic_1_targ_syscfg_apb_m_pprot),
    .aic_1_targ_syscfg_PRData(i_aic_1_targ_syscfg_apb_m_prdata),
    .aic_1_targ_syscfg_PReady(i_aic_1_targ_syscfg_apb_m_pready),
    .aic_1_targ_syscfg_PSel(o_aic_1_targ_syscfg_apb_m_psel),
    .aic_1_targ_syscfg_PSlvErr(i_aic_1_targ_syscfg_apb_m_pslverr),
    .aic_1_targ_syscfg_PStrb(o_aic_1_targ_syscfg_apb_m_pstrb),
    .aic_1_targ_syscfg_PWData(o_aic_1_targ_syscfg_apb_m_pwdata),
    .aic_1_targ_syscfg_PWrite(o_aic_1_targ_syscfg_apb_m_pwrite),
    .aic_2_aon_clk(i_aic_2_aon_clk),
    .aic_2_aon_rst_n(i_aic_2_aon_rst_n),
    .aic_2_clk(i_aic_2_clk),
    .aic_2_clken(i_aic_2_clken),
    .aic_2_init_ht_rd_Ar_Addr(aic_2_init_ht_axi_s_araddr_msb_fixed),
    .aic_2_init_ht_rd_Ar_Burst(i_aic_2_init_ht_axi_s_arburst),
    .aic_2_init_ht_rd_Ar_Cache(i_aic_2_init_ht_axi_s_arcache),
    .aic_2_init_ht_rd_Ar_Id(i_aic_2_init_ht_axi_s_arid),
    .aic_2_init_ht_rd_Ar_Len(i_aic_2_init_ht_axi_s_arlen),
    .aic_2_init_ht_rd_Ar_Lock(i_aic_2_init_ht_axi_s_arlock),
    .aic_2_init_ht_rd_Ar_Prot(i_aic_2_init_ht_axi_s_arprot),
    .aic_2_init_ht_rd_Ar_Ready(o_aic_2_init_ht_axi_s_arready),
    .aic_2_init_ht_rd_Ar_Size(i_aic_2_init_ht_axi_s_arsize),
    .aic_2_init_ht_rd_Ar_Valid(i_aic_2_init_ht_axi_s_arvalid),
    .aic_2_init_ht_rd_R_Data(o_aic_2_init_ht_axi_s_rdata),
    .aic_2_init_ht_rd_R_Id(o_aic_2_init_ht_axi_s_rid),
    .aic_2_init_ht_rd_R_Last(o_aic_2_init_ht_axi_s_rlast),
    .aic_2_init_ht_rd_R_Ready(i_aic_2_init_ht_axi_s_rready),
    .aic_2_init_ht_rd_R_Resp(o_aic_2_init_ht_axi_s_rresp),
    .aic_2_init_ht_rd_R_Valid(o_aic_2_init_ht_axi_s_rvalid),
    .aic_2_init_ht_wr_Aw_Addr(aic_2_init_ht_axi_s_awaddr_msb_fixed),
    .aic_2_init_ht_wr_Aw_Burst(i_aic_2_init_ht_axi_s_awburst),
    .aic_2_init_ht_wr_Aw_Cache(i_aic_2_init_ht_axi_s_awcache),
    .aic_2_init_ht_wr_Aw_Id(i_aic_2_init_ht_axi_s_awid),
    .aic_2_init_ht_wr_Aw_Len(i_aic_2_init_ht_axi_s_awlen),
    .aic_2_init_ht_wr_Aw_Lock(i_aic_2_init_ht_axi_s_awlock),
    .aic_2_init_ht_wr_Aw_Prot(i_aic_2_init_ht_axi_s_awprot),
    .aic_2_init_ht_wr_Aw_Ready(o_aic_2_init_ht_axi_s_awready),
    .aic_2_init_ht_wr_Aw_Size(i_aic_2_init_ht_axi_s_awsize),
    .aic_2_init_ht_wr_Aw_Valid(i_aic_2_init_ht_axi_s_awvalid),
    .aic_2_init_ht_wr_B_Id(o_aic_2_init_ht_axi_s_bid),
    .aic_2_init_ht_wr_B_Ready(i_aic_2_init_ht_axi_s_bready),
    .aic_2_init_ht_wr_B_Resp(o_aic_2_init_ht_axi_s_bresp),
    .aic_2_init_ht_wr_B_Valid(o_aic_2_init_ht_axi_s_bvalid),
    .aic_2_init_ht_wr_W_Data(i_aic_2_init_ht_axi_s_wdata),
    .aic_2_init_ht_wr_W_Last(i_aic_2_init_ht_axi_s_wlast),
    .aic_2_init_ht_wr_W_Ready(o_aic_2_init_ht_axi_s_wready),
    .aic_2_init_ht_wr_W_Strb(i_aic_2_init_ht_axi_s_wstrb),
    .aic_2_init_ht_wr_W_Valid(i_aic_2_init_ht_axi_s_wvalid),
    .aic_2_init_lt_Ar_Addr(aic_2_init_lt_axi_s_araddr_msb_fixed),
    .aic_2_init_lt_Ar_Burst(i_aic_2_init_lt_axi_s_arburst),
    .aic_2_init_lt_Ar_Cache(i_aic_2_init_lt_axi_s_arcache),
    .aic_2_init_lt_Ar_Id(i_aic_2_init_lt_axi_s_arid),
    .aic_2_init_lt_Ar_Len(i_aic_2_init_lt_axi_s_arlen),
    .aic_2_init_lt_Ar_Lock(i_aic_2_init_lt_axi_s_arlock),
    .aic_2_init_lt_Ar_Prot(i_aic_2_init_lt_axi_s_arprot),
    .aic_2_init_lt_Ar_Qos(i_aic_2_init_lt_axi_s_arqos),
    .aic_2_init_lt_Ar_Ready(o_aic_2_init_lt_axi_s_arready),
    .aic_2_init_lt_Ar_Size(i_aic_2_init_lt_axi_s_arsize),
    .aic_2_init_lt_Ar_Valid(i_aic_2_init_lt_axi_s_arvalid),
    .aic_2_init_lt_Aw_Addr(aic_2_init_lt_axi_s_awaddr_msb_fixed),
    .aic_2_init_lt_Aw_Burst(i_aic_2_init_lt_axi_s_awburst),
    .aic_2_init_lt_Aw_Cache(i_aic_2_init_lt_axi_s_awcache),
    .aic_2_init_lt_Aw_Id(i_aic_2_init_lt_axi_s_awid),
    .aic_2_init_lt_Aw_Len(i_aic_2_init_lt_axi_s_awlen),
    .aic_2_init_lt_Aw_Lock(i_aic_2_init_lt_axi_s_awlock),
    .aic_2_init_lt_Aw_Prot(i_aic_2_init_lt_axi_s_awprot),
    .aic_2_init_lt_Aw_Qos(i_aic_2_init_lt_axi_s_awqos),
    .aic_2_init_lt_Aw_Ready(o_aic_2_init_lt_axi_s_awready),
    .aic_2_init_lt_Aw_Size(i_aic_2_init_lt_axi_s_awsize),
    .aic_2_init_lt_Aw_Valid(i_aic_2_init_lt_axi_s_awvalid),
    .aic_2_init_lt_B_Id(o_aic_2_init_lt_axi_s_bid),
    .aic_2_init_lt_B_Ready(i_aic_2_init_lt_axi_s_bready),
    .aic_2_init_lt_B_Resp(o_aic_2_init_lt_axi_s_bresp),
    .aic_2_init_lt_B_Valid(o_aic_2_init_lt_axi_s_bvalid),
    .aic_2_init_lt_R_Data(o_aic_2_init_lt_axi_s_rdata),
    .aic_2_init_lt_R_Id(o_aic_2_init_lt_axi_s_rid),
    .aic_2_init_lt_R_Last(o_aic_2_init_lt_axi_s_rlast),
    .aic_2_init_lt_R_Ready(i_aic_2_init_lt_axi_s_rready),
    .aic_2_init_lt_R_Resp(o_aic_2_init_lt_axi_s_rresp),
    .aic_2_init_lt_R_Valid(o_aic_2_init_lt_axi_s_rvalid),
    .aic_2_init_lt_W_Data(i_aic_2_init_lt_axi_s_wdata),
    .aic_2_init_lt_W_Last(i_aic_2_init_lt_axi_s_wlast),
    .aic_2_init_lt_W_Ready(o_aic_2_init_lt_axi_s_wready),
    .aic_2_init_lt_W_Strb(i_aic_2_init_lt_axi_s_wstrb),
    .aic_2_init_lt_W_Valid(i_aic_2_init_lt_axi_s_wvalid),
    .aic_2_pwr_Idle(o_aic_2_pwr_idle_val),
    .aic_2_pwr_IdleAck(o_aic_2_pwr_idle_ack),
    .aic_2_pwr_IdleReq(i_aic_2_pwr_idle_req),
    .aic_2_rst_n(i_aic_2_rst_n),
    .aic_2_targ_lt_Ar_Addr(aic_2_targ_lt_axi_m_araddr_msb_fixed),
    .aic_2_targ_lt_Ar_Burst(o_aic_2_targ_lt_axi_m_arburst),
    .aic_2_targ_lt_Ar_Cache(o_aic_2_targ_lt_axi_m_arcache),
    .aic_2_targ_lt_Ar_Id(o_aic_2_targ_lt_axi_m_arid),
    .aic_2_targ_lt_Ar_Len(o_aic_2_targ_lt_axi_m_arlen),
    .aic_2_targ_lt_Ar_Lock(o_aic_2_targ_lt_axi_m_arlock),
    .aic_2_targ_lt_Ar_Prot(o_aic_2_targ_lt_axi_m_arprot),
    .aic_2_targ_lt_Ar_Qos(o_aic_2_targ_lt_axi_m_arqos),
    .aic_2_targ_lt_Ar_Ready(i_aic_2_targ_lt_axi_m_arready),
    .aic_2_targ_lt_Ar_Size(o_aic_2_targ_lt_axi_m_arsize),
    .aic_2_targ_lt_Ar_Valid(o_aic_2_targ_lt_axi_m_arvalid),
    .aic_2_targ_lt_Aw_Addr(aic_2_targ_lt_axi_m_awaddr_msb_fixed),
    .aic_2_targ_lt_Aw_Burst(o_aic_2_targ_lt_axi_m_awburst),
    .aic_2_targ_lt_Aw_Cache(o_aic_2_targ_lt_axi_m_awcache),
    .aic_2_targ_lt_Aw_Id(o_aic_2_targ_lt_axi_m_awid),
    .aic_2_targ_lt_Aw_Len(o_aic_2_targ_lt_axi_m_awlen),
    .aic_2_targ_lt_Aw_Lock(o_aic_2_targ_lt_axi_m_awlock),
    .aic_2_targ_lt_Aw_Prot(o_aic_2_targ_lt_axi_m_awprot),
    .aic_2_targ_lt_Aw_Qos(o_aic_2_targ_lt_axi_m_awqos),
    .aic_2_targ_lt_Aw_Ready(i_aic_2_targ_lt_axi_m_awready),
    .aic_2_targ_lt_Aw_Size(o_aic_2_targ_lt_axi_m_awsize),
    .aic_2_targ_lt_Aw_Valid(o_aic_2_targ_lt_axi_m_awvalid),
    .aic_2_targ_lt_B_Id(i_aic_2_targ_lt_axi_m_bid),
    .aic_2_targ_lt_B_Ready(o_aic_2_targ_lt_axi_m_bready),
    .aic_2_targ_lt_B_Resp(i_aic_2_targ_lt_axi_m_bresp),
    .aic_2_targ_lt_B_Valid(i_aic_2_targ_lt_axi_m_bvalid),
    .aic_2_targ_lt_R_Data(i_aic_2_targ_lt_axi_m_rdata),
    .aic_2_targ_lt_R_Id(i_aic_2_targ_lt_axi_m_rid),
    .aic_2_targ_lt_R_Last(i_aic_2_targ_lt_axi_m_rlast),
    .aic_2_targ_lt_R_Ready(o_aic_2_targ_lt_axi_m_rready),
    .aic_2_targ_lt_R_Resp(i_aic_2_targ_lt_axi_m_rresp),
    .aic_2_targ_lt_R_Valid(i_aic_2_targ_lt_axi_m_rvalid),
    .aic_2_targ_lt_W_Data(o_aic_2_targ_lt_axi_m_wdata),
    .aic_2_targ_lt_W_Last(o_aic_2_targ_lt_axi_m_wlast),
    .aic_2_targ_lt_W_Ready(i_aic_2_targ_lt_axi_m_wready),
    .aic_2_targ_lt_W_Strb(o_aic_2_targ_lt_axi_m_wstrb),
    .aic_2_targ_lt_W_Valid(o_aic_2_targ_lt_axi_m_wvalid),
    .aic_2_targ_syscfg_PAddr(o_aic_2_targ_syscfg_apb_m_paddr),
    .aic_2_targ_syscfg_PEnable(o_aic_2_targ_syscfg_apb_m_penable),
    .aic_2_targ_syscfg_PProt(o_aic_2_targ_syscfg_apb_m_pprot),
    .aic_2_targ_syscfg_PRData(i_aic_2_targ_syscfg_apb_m_prdata),
    .aic_2_targ_syscfg_PReady(i_aic_2_targ_syscfg_apb_m_pready),
    .aic_2_targ_syscfg_PSel(o_aic_2_targ_syscfg_apb_m_psel),
    .aic_2_targ_syscfg_PSlvErr(i_aic_2_targ_syscfg_apb_m_pslverr),
    .aic_2_targ_syscfg_PStrb(o_aic_2_targ_syscfg_apb_m_pstrb),
    .aic_2_targ_syscfg_PWData(o_aic_2_targ_syscfg_apb_m_pwdata),
    .aic_2_targ_syscfg_PWrite(o_aic_2_targ_syscfg_apb_m_pwrite),
    .aic_3_aon_clk(i_aic_3_aon_clk),
    .aic_3_aon_rst_n(i_aic_3_aon_rst_n),
    .aic_3_clk(i_aic_3_clk),
    .aic_3_clken(i_aic_3_clken),
    .aic_3_init_ht_rd_Ar_Addr(aic_3_init_ht_axi_s_araddr_msb_fixed),
    .aic_3_init_ht_rd_Ar_Burst(i_aic_3_init_ht_axi_s_arburst),
    .aic_3_init_ht_rd_Ar_Cache(i_aic_3_init_ht_axi_s_arcache),
    .aic_3_init_ht_rd_Ar_Id(i_aic_3_init_ht_axi_s_arid),
    .aic_3_init_ht_rd_Ar_Len(i_aic_3_init_ht_axi_s_arlen),
    .aic_3_init_ht_rd_Ar_Lock(i_aic_3_init_ht_axi_s_arlock),
    .aic_3_init_ht_rd_Ar_Prot(i_aic_3_init_ht_axi_s_arprot),
    .aic_3_init_ht_rd_Ar_Ready(o_aic_3_init_ht_axi_s_arready),
    .aic_3_init_ht_rd_Ar_Size(i_aic_3_init_ht_axi_s_arsize),
    .aic_3_init_ht_rd_Ar_Valid(i_aic_3_init_ht_axi_s_arvalid),
    .aic_3_init_ht_rd_R_Data(o_aic_3_init_ht_axi_s_rdata),
    .aic_3_init_ht_rd_R_Id(o_aic_3_init_ht_axi_s_rid),
    .aic_3_init_ht_rd_R_Last(o_aic_3_init_ht_axi_s_rlast),
    .aic_3_init_ht_rd_R_Ready(i_aic_3_init_ht_axi_s_rready),
    .aic_3_init_ht_rd_R_Resp(o_aic_3_init_ht_axi_s_rresp),
    .aic_3_init_ht_rd_R_Valid(o_aic_3_init_ht_axi_s_rvalid),
    .aic_3_init_ht_wr_Aw_Addr(aic_3_init_ht_axi_s_awaddr_msb_fixed),
    .aic_3_init_ht_wr_Aw_Burst(i_aic_3_init_ht_axi_s_awburst),
    .aic_3_init_ht_wr_Aw_Cache(i_aic_3_init_ht_axi_s_awcache),
    .aic_3_init_ht_wr_Aw_Id(i_aic_3_init_ht_axi_s_awid),
    .aic_3_init_ht_wr_Aw_Len(i_aic_3_init_ht_axi_s_awlen),
    .aic_3_init_ht_wr_Aw_Lock(i_aic_3_init_ht_axi_s_awlock),
    .aic_3_init_ht_wr_Aw_Prot(i_aic_3_init_ht_axi_s_awprot),
    .aic_3_init_ht_wr_Aw_Ready(o_aic_3_init_ht_axi_s_awready),
    .aic_3_init_ht_wr_Aw_Size(i_aic_3_init_ht_axi_s_awsize),
    .aic_3_init_ht_wr_Aw_Valid(i_aic_3_init_ht_axi_s_awvalid),
    .aic_3_init_ht_wr_B_Id(o_aic_3_init_ht_axi_s_bid),
    .aic_3_init_ht_wr_B_Ready(i_aic_3_init_ht_axi_s_bready),
    .aic_3_init_ht_wr_B_Resp(o_aic_3_init_ht_axi_s_bresp),
    .aic_3_init_ht_wr_B_Valid(o_aic_3_init_ht_axi_s_bvalid),
    .aic_3_init_ht_wr_W_Data(i_aic_3_init_ht_axi_s_wdata),
    .aic_3_init_ht_wr_W_Last(i_aic_3_init_ht_axi_s_wlast),
    .aic_3_init_ht_wr_W_Ready(o_aic_3_init_ht_axi_s_wready),
    .aic_3_init_ht_wr_W_Strb(i_aic_3_init_ht_axi_s_wstrb),
    .aic_3_init_ht_wr_W_Valid(i_aic_3_init_ht_axi_s_wvalid),
    .aic_3_init_lt_Ar_Addr(aic_3_init_lt_axi_s_araddr_msb_fixed),
    .aic_3_init_lt_Ar_Burst(i_aic_3_init_lt_axi_s_arburst),
    .aic_3_init_lt_Ar_Cache(i_aic_3_init_lt_axi_s_arcache),
    .aic_3_init_lt_Ar_Id(i_aic_3_init_lt_axi_s_arid),
    .aic_3_init_lt_Ar_Len(i_aic_3_init_lt_axi_s_arlen),
    .aic_3_init_lt_Ar_Lock(i_aic_3_init_lt_axi_s_arlock),
    .aic_3_init_lt_Ar_Prot(i_aic_3_init_lt_axi_s_arprot),
    .aic_3_init_lt_Ar_Qos(i_aic_3_init_lt_axi_s_arqos),
    .aic_3_init_lt_Ar_Ready(o_aic_3_init_lt_axi_s_arready),
    .aic_3_init_lt_Ar_Size(i_aic_3_init_lt_axi_s_arsize),
    .aic_3_init_lt_Ar_Valid(i_aic_3_init_lt_axi_s_arvalid),
    .aic_3_init_lt_Aw_Addr(aic_3_init_lt_axi_s_awaddr_msb_fixed),
    .aic_3_init_lt_Aw_Burst(i_aic_3_init_lt_axi_s_awburst),
    .aic_3_init_lt_Aw_Cache(i_aic_3_init_lt_axi_s_awcache),
    .aic_3_init_lt_Aw_Id(i_aic_3_init_lt_axi_s_awid),
    .aic_3_init_lt_Aw_Len(i_aic_3_init_lt_axi_s_awlen),
    .aic_3_init_lt_Aw_Lock(i_aic_3_init_lt_axi_s_awlock),
    .aic_3_init_lt_Aw_Prot(i_aic_3_init_lt_axi_s_awprot),
    .aic_3_init_lt_Aw_Qos(i_aic_3_init_lt_axi_s_awqos),
    .aic_3_init_lt_Aw_Ready(o_aic_3_init_lt_axi_s_awready),
    .aic_3_init_lt_Aw_Size(i_aic_3_init_lt_axi_s_awsize),
    .aic_3_init_lt_Aw_Valid(i_aic_3_init_lt_axi_s_awvalid),
    .aic_3_init_lt_B_Id(o_aic_3_init_lt_axi_s_bid),
    .aic_3_init_lt_B_Ready(i_aic_3_init_lt_axi_s_bready),
    .aic_3_init_lt_B_Resp(o_aic_3_init_lt_axi_s_bresp),
    .aic_3_init_lt_B_Valid(o_aic_3_init_lt_axi_s_bvalid),
    .aic_3_init_lt_R_Data(o_aic_3_init_lt_axi_s_rdata),
    .aic_3_init_lt_R_Id(o_aic_3_init_lt_axi_s_rid),
    .aic_3_init_lt_R_Last(o_aic_3_init_lt_axi_s_rlast),
    .aic_3_init_lt_R_Ready(i_aic_3_init_lt_axi_s_rready),
    .aic_3_init_lt_R_Resp(o_aic_3_init_lt_axi_s_rresp),
    .aic_3_init_lt_R_Valid(o_aic_3_init_lt_axi_s_rvalid),
    .aic_3_init_lt_W_Data(i_aic_3_init_lt_axi_s_wdata),
    .aic_3_init_lt_W_Last(i_aic_3_init_lt_axi_s_wlast),
    .aic_3_init_lt_W_Ready(o_aic_3_init_lt_axi_s_wready),
    .aic_3_init_lt_W_Strb(i_aic_3_init_lt_axi_s_wstrb),
    .aic_3_init_lt_W_Valid(i_aic_3_init_lt_axi_s_wvalid),
    .aic_3_pwr_Idle(o_aic_3_pwr_idle_val),
    .aic_3_pwr_IdleAck(o_aic_3_pwr_idle_ack),
    .aic_3_pwr_IdleReq(i_aic_3_pwr_idle_req),
    .aic_3_rst_n(i_aic_3_rst_n),
    .aic_3_targ_lt_Ar_Addr(aic_3_targ_lt_axi_m_araddr_msb_fixed),
    .aic_3_targ_lt_Ar_Burst(o_aic_3_targ_lt_axi_m_arburst),
    .aic_3_targ_lt_Ar_Cache(o_aic_3_targ_lt_axi_m_arcache),
    .aic_3_targ_lt_Ar_Id(o_aic_3_targ_lt_axi_m_arid),
    .aic_3_targ_lt_Ar_Len(o_aic_3_targ_lt_axi_m_arlen),
    .aic_3_targ_lt_Ar_Lock(o_aic_3_targ_lt_axi_m_arlock),
    .aic_3_targ_lt_Ar_Prot(o_aic_3_targ_lt_axi_m_arprot),
    .aic_3_targ_lt_Ar_Qos(o_aic_3_targ_lt_axi_m_arqos),
    .aic_3_targ_lt_Ar_Ready(i_aic_3_targ_lt_axi_m_arready),
    .aic_3_targ_lt_Ar_Size(o_aic_3_targ_lt_axi_m_arsize),
    .aic_3_targ_lt_Ar_Valid(o_aic_3_targ_lt_axi_m_arvalid),
    .aic_3_targ_lt_Aw_Addr(aic_3_targ_lt_axi_m_awaddr_msb_fixed),
    .aic_3_targ_lt_Aw_Burst(o_aic_3_targ_lt_axi_m_awburst),
    .aic_3_targ_lt_Aw_Cache(o_aic_3_targ_lt_axi_m_awcache),
    .aic_3_targ_lt_Aw_Id(o_aic_3_targ_lt_axi_m_awid),
    .aic_3_targ_lt_Aw_Len(o_aic_3_targ_lt_axi_m_awlen),
    .aic_3_targ_lt_Aw_Lock(o_aic_3_targ_lt_axi_m_awlock),
    .aic_3_targ_lt_Aw_Prot(o_aic_3_targ_lt_axi_m_awprot),
    .aic_3_targ_lt_Aw_Qos(o_aic_3_targ_lt_axi_m_awqos),
    .aic_3_targ_lt_Aw_Ready(i_aic_3_targ_lt_axi_m_awready),
    .aic_3_targ_lt_Aw_Size(o_aic_3_targ_lt_axi_m_awsize),
    .aic_3_targ_lt_Aw_Valid(o_aic_3_targ_lt_axi_m_awvalid),
    .aic_3_targ_lt_B_Id(i_aic_3_targ_lt_axi_m_bid),
    .aic_3_targ_lt_B_Ready(o_aic_3_targ_lt_axi_m_bready),
    .aic_3_targ_lt_B_Resp(i_aic_3_targ_lt_axi_m_bresp),
    .aic_3_targ_lt_B_Valid(i_aic_3_targ_lt_axi_m_bvalid),
    .aic_3_targ_lt_R_Data(i_aic_3_targ_lt_axi_m_rdata),
    .aic_3_targ_lt_R_Id(i_aic_3_targ_lt_axi_m_rid),
    .aic_3_targ_lt_R_Last(i_aic_3_targ_lt_axi_m_rlast),
    .aic_3_targ_lt_R_Ready(o_aic_3_targ_lt_axi_m_rready),
    .aic_3_targ_lt_R_Resp(i_aic_3_targ_lt_axi_m_rresp),
    .aic_3_targ_lt_R_Valid(i_aic_3_targ_lt_axi_m_rvalid),
    .aic_3_targ_lt_W_Data(o_aic_3_targ_lt_axi_m_wdata),
    .aic_3_targ_lt_W_Last(o_aic_3_targ_lt_axi_m_wlast),
    .aic_3_targ_lt_W_Ready(i_aic_3_targ_lt_axi_m_wready),
    .aic_3_targ_lt_W_Strb(o_aic_3_targ_lt_axi_m_wstrb),
    .aic_3_targ_lt_W_Valid(o_aic_3_targ_lt_axi_m_wvalid),
    .aic_3_targ_syscfg_PAddr(o_aic_3_targ_syscfg_apb_m_paddr),
    .aic_3_targ_syscfg_PEnable(o_aic_3_targ_syscfg_apb_m_penable),
    .aic_3_targ_syscfg_PProt(o_aic_3_targ_syscfg_apb_m_pprot),
    .aic_3_targ_syscfg_PRData(i_aic_3_targ_syscfg_apb_m_prdata),
    .aic_3_targ_syscfg_PReady(i_aic_3_targ_syscfg_apb_m_pready),
    .aic_3_targ_syscfg_PSel(o_aic_3_targ_syscfg_apb_m_psel),
    .aic_3_targ_syscfg_PSlvErr(i_aic_3_targ_syscfg_apb_m_pslverr),
    .aic_3_targ_syscfg_PStrb(o_aic_3_targ_syscfg_apb_m_pstrb),
    .aic_3_targ_syscfg_PWData(o_aic_3_targ_syscfg_apb_m_pwdata),
    .aic_3_targ_syscfg_PWrite(o_aic_3_targ_syscfg_apb_m_pwrite),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Data(i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Head(i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Data(i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Head(i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Data(i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Head(i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Data(i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Head(i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Data(i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Head(i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Data(i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Head(i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Data(i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Head(i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Data(i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Head(i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Data(i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Head(i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Data(i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Head(i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Data(i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Head(i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Data(i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Head(i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Data(i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Head(i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Rdy(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Tail(i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Vld(i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Data(o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Head(o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Rdy(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Tail(o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Vld(o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Data(o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Head(o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Rdy(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Tail(o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Vld(o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Data(i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Head(i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Data(o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Head(o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Rdy(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Tail(o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Vld(o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Data(i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Head(i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Data(o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Head(o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Rdy(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Tail(o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Vld(o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Data(i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Head(i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Data(o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Head(o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Rdy(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Tail(o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Vld(o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Data(i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Head(i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Data(o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Head(o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Rdy(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Tail(o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Vld(o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Data(i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Head(i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Data(o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Head(o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Rdy(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Tail(o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Vld(o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Data(i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Head(i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Data(o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Head(o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Rdy(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Tail(o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Vld(o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Data(i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Head(i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Data(o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Head(o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Rdy(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Tail(o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Vld(o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Data(i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Head(i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Data(o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Head(o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Rdy(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Tail(o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Vld(o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Data(i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Head(i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Data(o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Head(o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Rdy(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Tail(o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Vld(o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Data(i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Head(i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Data(o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Head(o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Rdy(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Tail(o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Vld(o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Data(i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Head(i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Data(o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Head(o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Rdy(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Tail(o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Vld(o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Data(i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Head(i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Rdy(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Tail(i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Vld(i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Data(o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Head(o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Rdy(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Tail(o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Vld(o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Data(i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Head(i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Rdy(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Tail(i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Vld(i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld),
    .l2_0_aon_clk(i_l2_0_aon_clk),
    .l2_0_aon_rst_n(i_l2_0_aon_rst_n),
    .l2_0_clk(i_l2_0_clk),
    .l2_0_clken(i_l2_0_clken),
    .l2_0_pwr_Idle(o_l2_0_pwr_idle_val),
    .l2_0_pwr_IdleAck(o_l2_0_pwr_idle_ack),
    .l2_0_pwr_IdleReq(i_l2_0_pwr_idle_req),
    .l2_0_rst_n(i_l2_0_rst_n),
    .l2_0_targ_ht_rd_Ar_Addr(l2_0_targ_ht_axi_m_araddr_msb_fixed),
    .l2_0_targ_ht_rd_Ar_Burst(o_l2_0_targ_ht_axi_m_arburst),
    .l2_0_targ_ht_rd_Ar_Cache(o_l2_0_targ_ht_axi_m_arcache),
    .l2_0_targ_ht_rd_Ar_Id(o_l2_0_targ_ht_axi_m_arid),
    .l2_0_targ_ht_rd_Ar_Len(o_l2_0_targ_ht_axi_m_arlen),
    .l2_0_targ_ht_rd_Ar_Lock(o_l2_0_targ_ht_axi_m_arlock),
    .l2_0_targ_ht_rd_Ar_Prot(o_l2_0_targ_ht_axi_m_arprot),
    .l2_0_targ_ht_rd_Ar_Ready(i_l2_0_targ_ht_axi_m_arready),
    .l2_0_targ_ht_rd_Ar_Size(o_l2_0_targ_ht_axi_m_arsize),
    .l2_0_targ_ht_rd_Ar_Valid(o_l2_0_targ_ht_axi_m_arvalid),
    .l2_0_targ_ht_rd_R_Data(i_l2_0_targ_ht_axi_m_rdata),
    .l2_0_targ_ht_rd_R_Id(i_l2_0_targ_ht_axi_m_rid),
    .l2_0_targ_ht_rd_R_Last(i_l2_0_targ_ht_axi_m_rlast),
    .l2_0_targ_ht_rd_R_Ready(o_l2_0_targ_ht_axi_m_rready),
    .l2_0_targ_ht_rd_R_Resp(i_l2_0_targ_ht_axi_m_rresp),
    .l2_0_targ_ht_rd_R_Valid(i_l2_0_targ_ht_axi_m_rvalid),
    .l2_0_targ_ht_wr_Aw_Addr(l2_0_targ_ht_axi_m_awaddr_msb_fixed),
    .l2_0_targ_ht_wr_Aw_Burst(o_l2_0_targ_ht_axi_m_awburst),
    .l2_0_targ_ht_wr_Aw_Cache(o_l2_0_targ_ht_axi_m_awcache),
    .l2_0_targ_ht_wr_Aw_Id(o_l2_0_targ_ht_axi_m_awid),
    .l2_0_targ_ht_wr_Aw_Len(o_l2_0_targ_ht_axi_m_awlen),
    .l2_0_targ_ht_wr_Aw_Lock(o_l2_0_targ_ht_axi_m_awlock),
    .l2_0_targ_ht_wr_Aw_Prot(o_l2_0_targ_ht_axi_m_awprot),
    .l2_0_targ_ht_wr_Aw_Ready(i_l2_0_targ_ht_axi_m_awready),
    .l2_0_targ_ht_wr_Aw_Size(o_l2_0_targ_ht_axi_m_awsize),
    .l2_0_targ_ht_wr_Aw_Valid(o_l2_0_targ_ht_axi_m_awvalid),
    .l2_0_targ_ht_wr_B_Id(i_l2_0_targ_ht_axi_m_bid),
    .l2_0_targ_ht_wr_B_Ready(o_l2_0_targ_ht_axi_m_bready),
    .l2_0_targ_ht_wr_B_Resp(i_l2_0_targ_ht_axi_m_bresp),
    .l2_0_targ_ht_wr_B_Valid(i_l2_0_targ_ht_axi_m_bvalid),
    .l2_0_targ_ht_wr_W_Data(o_l2_0_targ_ht_axi_m_wdata),
    .l2_0_targ_ht_wr_W_Last(o_l2_0_targ_ht_axi_m_wlast),
    .l2_0_targ_ht_wr_W_Ready(i_l2_0_targ_ht_axi_m_wready),
    .l2_0_targ_ht_wr_W_Strb(o_l2_0_targ_ht_axi_m_wstrb),
    .l2_0_targ_ht_wr_W_Valid(o_l2_0_targ_ht_axi_m_wvalid),
    .l2_0_targ_syscfg_PAddr(o_l2_0_targ_syscfg_apb_m_paddr),
    .l2_0_targ_syscfg_PEnable(o_l2_0_targ_syscfg_apb_m_penable),
    .l2_0_targ_syscfg_PProt(o_l2_0_targ_syscfg_apb_m_pprot),
    .l2_0_targ_syscfg_PRData(i_l2_0_targ_syscfg_apb_m_prdata),
    .l2_0_targ_syscfg_PReady(i_l2_0_targ_syscfg_apb_m_pready),
    .l2_0_targ_syscfg_PSel(o_l2_0_targ_syscfg_apb_m_psel),
    .l2_0_targ_syscfg_PSlvErr(i_l2_0_targ_syscfg_apb_m_pslverr),
    .l2_0_targ_syscfg_PStrb(o_l2_0_targ_syscfg_apb_m_pstrb),
    .l2_0_targ_syscfg_PWData(o_l2_0_targ_syscfg_apb_m_pwdata),
    .l2_0_targ_syscfg_PWrite(o_l2_0_targ_syscfg_apb_m_pwrite),
    .l2_1_aon_clk(i_l2_1_aon_clk),
    .l2_1_aon_rst_n(i_l2_1_aon_rst_n),
    .l2_1_clk(i_l2_1_clk),
    .l2_1_clken(i_l2_1_clken),
    .l2_1_pwr_Idle(o_l2_1_pwr_idle_val),
    .l2_1_pwr_IdleAck(o_l2_1_pwr_idle_ack),
    .l2_1_pwr_IdleReq(i_l2_1_pwr_idle_req),
    .l2_1_rst_n(i_l2_1_rst_n),
    .l2_1_targ_ht_rd_Ar_Addr(l2_1_targ_ht_axi_m_araddr_msb_fixed),
    .l2_1_targ_ht_rd_Ar_Burst(o_l2_1_targ_ht_axi_m_arburst),
    .l2_1_targ_ht_rd_Ar_Cache(o_l2_1_targ_ht_axi_m_arcache),
    .l2_1_targ_ht_rd_Ar_Id(o_l2_1_targ_ht_axi_m_arid),
    .l2_1_targ_ht_rd_Ar_Len(o_l2_1_targ_ht_axi_m_arlen),
    .l2_1_targ_ht_rd_Ar_Lock(o_l2_1_targ_ht_axi_m_arlock),
    .l2_1_targ_ht_rd_Ar_Prot(o_l2_1_targ_ht_axi_m_arprot),
    .l2_1_targ_ht_rd_Ar_Ready(i_l2_1_targ_ht_axi_m_arready),
    .l2_1_targ_ht_rd_Ar_Size(o_l2_1_targ_ht_axi_m_arsize),
    .l2_1_targ_ht_rd_Ar_Valid(o_l2_1_targ_ht_axi_m_arvalid),
    .l2_1_targ_ht_rd_R_Data(i_l2_1_targ_ht_axi_m_rdata),
    .l2_1_targ_ht_rd_R_Id(i_l2_1_targ_ht_axi_m_rid),
    .l2_1_targ_ht_rd_R_Last(i_l2_1_targ_ht_axi_m_rlast),
    .l2_1_targ_ht_rd_R_Ready(o_l2_1_targ_ht_axi_m_rready),
    .l2_1_targ_ht_rd_R_Resp(i_l2_1_targ_ht_axi_m_rresp),
    .l2_1_targ_ht_rd_R_Valid(i_l2_1_targ_ht_axi_m_rvalid),
    .l2_1_targ_ht_wr_Aw_Addr(l2_1_targ_ht_axi_m_awaddr_msb_fixed),
    .l2_1_targ_ht_wr_Aw_Burst(o_l2_1_targ_ht_axi_m_awburst),
    .l2_1_targ_ht_wr_Aw_Cache(o_l2_1_targ_ht_axi_m_awcache),
    .l2_1_targ_ht_wr_Aw_Id(o_l2_1_targ_ht_axi_m_awid),
    .l2_1_targ_ht_wr_Aw_Len(o_l2_1_targ_ht_axi_m_awlen),
    .l2_1_targ_ht_wr_Aw_Lock(o_l2_1_targ_ht_axi_m_awlock),
    .l2_1_targ_ht_wr_Aw_Prot(o_l2_1_targ_ht_axi_m_awprot),
    .l2_1_targ_ht_wr_Aw_Ready(i_l2_1_targ_ht_axi_m_awready),
    .l2_1_targ_ht_wr_Aw_Size(o_l2_1_targ_ht_axi_m_awsize),
    .l2_1_targ_ht_wr_Aw_Valid(o_l2_1_targ_ht_axi_m_awvalid),
    .l2_1_targ_ht_wr_B_Id(i_l2_1_targ_ht_axi_m_bid),
    .l2_1_targ_ht_wr_B_Ready(o_l2_1_targ_ht_axi_m_bready),
    .l2_1_targ_ht_wr_B_Resp(i_l2_1_targ_ht_axi_m_bresp),
    .l2_1_targ_ht_wr_B_Valid(i_l2_1_targ_ht_axi_m_bvalid),
    .l2_1_targ_ht_wr_W_Data(o_l2_1_targ_ht_axi_m_wdata),
    .l2_1_targ_ht_wr_W_Last(o_l2_1_targ_ht_axi_m_wlast),
    .l2_1_targ_ht_wr_W_Ready(i_l2_1_targ_ht_axi_m_wready),
    .l2_1_targ_ht_wr_W_Strb(o_l2_1_targ_ht_axi_m_wstrb),
    .l2_1_targ_ht_wr_W_Valid(o_l2_1_targ_ht_axi_m_wvalid),
    .l2_1_targ_syscfg_PAddr(o_l2_1_targ_syscfg_apb_m_paddr),
    .l2_1_targ_syscfg_PEnable(o_l2_1_targ_syscfg_apb_m_penable),
    .l2_1_targ_syscfg_PProt(o_l2_1_targ_syscfg_apb_m_pprot),
    .l2_1_targ_syscfg_PRData(i_l2_1_targ_syscfg_apb_m_prdata),
    .l2_1_targ_syscfg_PReady(i_l2_1_targ_syscfg_apb_m_pready),
    .l2_1_targ_syscfg_PSel(o_l2_1_targ_syscfg_apb_m_psel),
    .l2_1_targ_syscfg_PSlvErr(i_l2_1_targ_syscfg_apb_m_pslverr),
    .l2_1_targ_syscfg_PStrb(o_l2_1_targ_syscfg_apb_m_pstrb),
    .l2_1_targ_syscfg_PWData(o_l2_1_targ_syscfg_apb_m_pwdata),
    .l2_1_targ_syscfg_PWrite(o_l2_1_targ_syscfg_apb_m_pwrite),
    .l2_2_aon_clk(i_l2_2_aon_clk),
    .l2_2_aon_rst_n(i_l2_2_aon_rst_n),
    .l2_2_clk(i_l2_2_clk),
    .l2_2_clken(i_l2_2_clken),
    .l2_2_pwr_Idle(o_l2_2_pwr_idle_val),
    .l2_2_pwr_IdleAck(o_l2_2_pwr_idle_ack),
    .l2_2_pwr_IdleReq(i_l2_2_pwr_idle_req),
    .l2_2_rst_n(i_l2_2_rst_n),
    .l2_2_targ_ht_rd_Ar_Addr(l2_2_targ_ht_axi_m_araddr_msb_fixed),
    .l2_2_targ_ht_rd_Ar_Burst(o_l2_2_targ_ht_axi_m_arburst),
    .l2_2_targ_ht_rd_Ar_Cache(o_l2_2_targ_ht_axi_m_arcache),
    .l2_2_targ_ht_rd_Ar_Id(o_l2_2_targ_ht_axi_m_arid),
    .l2_2_targ_ht_rd_Ar_Len(o_l2_2_targ_ht_axi_m_arlen),
    .l2_2_targ_ht_rd_Ar_Lock(o_l2_2_targ_ht_axi_m_arlock),
    .l2_2_targ_ht_rd_Ar_Prot(o_l2_2_targ_ht_axi_m_arprot),
    .l2_2_targ_ht_rd_Ar_Ready(i_l2_2_targ_ht_axi_m_arready),
    .l2_2_targ_ht_rd_Ar_Size(o_l2_2_targ_ht_axi_m_arsize),
    .l2_2_targ_ht_rd_Ar_Valid(o_l2_2_targ_ht_axi_m_arvalid),
    .l2_2_targ_ht_rd_R_Data(i_l2_2_targ_ht_axi_m_rdata),
    .l2_2_targ_ht_rd_R_Id(i_l2_2_targ_ht_axi_m_rid),
    .l2_2_targ_ht_rd_R_Last(i_l2_2_targ_ht_axi_m_rlast),
    .l2_2_targ_ht_rd_R_Ready(o_l2_2_targ_ht_axi_m_rready),
    .l2_2_targ_ht_rd_R_Resp(i_l2_2_targ_ht_axi_m_rresp),
    .l2_2_targ_ht_rd_R_Valid(i_l2_2_targ_ht_axi_m_rvalid),
    .l2_2_targ_ht_wr_Aw_Addr(l2_2_targ_ht_axi_m_awaddr_msb_fixed),
    .l2_2_targ_ht_wr_Aw_Burst(o_l2_2_targ_ht_axi_m_awburst),
    .l2_2_targ_ht_wr_Aw_Cache(o_l2_2_targ_ht_axi_m_awcache),
    .l2_2_targ_ht_wr_Aw_Id(o_l2_2_targ_ht_axi_m_awid),
    .l2_2_targ_ht_wr_Aw_Len(o_l2_2_targ_ht_axi_m_awlen),
    .l2_2_targ_ht_wr_Aw_Lock(o_l2_2_targ_ht_axi_m_awlock),
    .l2_2_targ_ht_wr_Aw_Prot(o_l2_2_targ_ht_axi_m_awprot),
    .l2_2_targ_ht_wr_Aw_Ready(i_l2_2_targ_ht_axi_m_awready),
    .l2_2_targ_ht_wr_Aw_Size(o_l2_2_targ_ht_axi_m_awsize),
    .l2_2_targ_ht_wr_Aw_Valid(o_l2_2_targ_ht_axi_m_awvalid),
    .l2_2_targ_ht_wr_B_Id(i_l2_2_targ_ht_axi_m_bid),
    .l2_2_targ_ht_wr_B_Ready(o_l2_2_targ_ht_axi_m_bready),
    .l2_2_targ_ht_wr_B_Resp(i_l2_2_targ_ht_axi_m_bresp),
    .l2_2_targ_ht_wr_B_Valid(i_l2_2_targ_ht_axi_m_bvalid),
    .l2_2_targ_ht_wr_W_Data(o_l2_2_targ_ht_axi_m_wdata),
    .l2_2_targ_ht_wr_W_Last(o_l2_2_targ_ht_axi_m_wlast),
    .l2_2_targ_ht_wr_W_Ready(i_l2_2_targ_ht_axi_m_wready),
    .l2_2_targ_ht_wr_W_Strb(o_l2_2_targ_ht_axi_m_wstrb),
    .l2_2_targ_ht_wr_W_Valid(o_l2_2_targ_ht_axi_m_wvalid),
    .l2_2_targ_syscfg_PAddr(o_l2_2_targ_syscfg_apb_m_paddr),
    .l2_2_targ_syscfg_PEnable(o_l2_2_targ_syscfg_apb_m_penable),
    .l2_2_targ_syscfg_PProt(o_l2_2_targ_syscfg_apb_m_pprot),
    .l2_2_targ_syscfg_PRData(i_l2_2_targ_syscfg_apb_m_prdata),
    .l2_2_targ_syscfg_PReady(i_l2_2_targ_syscfg_apb_m_pready),
    .l2_2_targ_syscfg_PSel(o_l2_2_targ_syscfg_apb_m_psel),
    .l2_2_targ_syscfg_PSlvErr(i_l2_2_targ_syscfg_apb_m_pslverr),
    .l2_2_targ_syscfg_PStrb(o_l2_2_targ_syscfg_apb_m_pstrb),
    .l2_2_targ_syscfg_PWData(o_l2_2_targ_syscfg_apb_m_pwdata),
    .l2_2_targ_syscfg_PWrite(o_l2_2_targ_syscfg_apb_m_pwrite),
    .l2_3_aon_clk(i_l2_3_aon_clk),
    .l2_3_aon_rst_n(i_l2_3_aon_rst_n),
    .l2_3_clk(i_l2_3_clk),
    .l2_3_clken(i_l2_3_clken),
    .l2_3_pwr_Idle(o_l2_3_pwr_idle_val),
    .l2_3_pwr_IdleAck(o_l2_3_pwr_idle_ack),
    .l2_3_pwr_IdleReq(i_l2_3_pwr_idle_req),
    .l2_3_rst_n(i_l2_3_rst_n),
    .l2_3_targ_ht_rd_Ar_Addr(l2_3_targ_ht_axi_m_araddr_msb_fixed),
    .l2_3_targ_ht_rd_Ar_Burst(o_l2_3_targ_ht_axi_m_arburst),
    .l2_3_targ_ht_rd_Ar_Cache(o_l2_3_targ_ht_axi_m_arcache),
    .l2_3_targ_ht_rd_Ar_Id(o_l2_3_targ_ht_axi_m_arid),
    .l2_3_targ_ht_rd_Ar_Len(o_l2_3_targ_ht_axi_m_arlen),
    .l2_3_targ_ht_rd_Ar_Lock(o_l2_3_targ_ht_axi_m_arlock),
    .l2_3_targ_ht_rd_Ar_Prot(o_l2_3_targ_ht_axi_m_arprot),
    .l2_3_targ_ht_rd_Ar_Ready(i_l2_3_targ_ht_axi_m_arready),
    .l2_3_targ_ht_rd_Ar_Size(o_l2_3_targ_ht_axi_m_arsize),
    .l2_3_targ_ht_rd_Ar_Valid(o_l2_3_targ_ht_axi_m_arvalid),
    .l2_3_targ_ht_rd_R_Data(i_l2_3_targ_ht_axi_m_rdata),
    .l2_3_targ_ht_rd_R_Id(i_l2_3_targ_ht_axi_m_rid),
    .l2_3_targ_ht_rd_R_Last(i_l2_3_targ_ht_axi_m_rlast),
    .l2_3_targ_ht_rd_R_Ready(o_l2_3_targ_ht_axi_m_rready),
    .l2_3_targ_ht_rd_R_Resp(i_l2_3_targ_ht_axi_m_rresp),
    .l2_3_targ_ht_rd_R_Valid(i_l2_3_targ_ht_axi_m_rvalid),
    .l2_3_targ_ht_wr_Aw_Addr(l2_3_targ_ht_axi_m_awaddr_msb_fixed),
    .l2_3_targ_ht_wr_Aw_Burst(o_l2_3_targ_ht_axi_m_awburst),
    .l2_3_targ_ht_wr_Aw_Cache(o_l2_3_targ_ht_axi_m_awcache),
    .l2_3_targ_ht_wr_Aw_Id(o_l2_3_targ_ht_axi_m_awid),
    .l2_3_targ_ht_wr_Aw_Len(o_l2_3_targ_ht_axi_m_awlen),
    .l2_3_targ_ht_wr_Aw_Lock(o_l2_3_targ_ht_axi_m_awlock),
    .l2_3_targ_ht_wr_Aw_Prot(o_l2_3_targ_ht_axi_m_awprot),
    .l2_3_targ_ht_wr_Aw_Ready(i_l2_3_targ_ht_axi_m_awready),
    .l2_3_targ_ht_wr_Aw_Size(o_l2_3_targ_ht_axi_m_awsize),
    .l2_3_targ_ht_wr_Aw_Valid(o_l2_3_targ_ht_axi_m_awvalid),
    .l2_3_targ_ht_wr_B_Id(i_l2_3_targ_ht_axi_m_bid),
    .l2_3_targ_ht_wr_B_Ready(o_l2_3_targ_ht_axi_m_bready),
    .l2_3_targ_ht_wr_B_Resp(i_l2_3_targ_ht_axi_m_bresp),
    .l2_3_targ_ht_wr_B_Valid(i_l2_3_targ_ht_axi_m_bvalid),
    .l2_3_targ_ht_wr_W_Data(o_l2_3_targ_ht_axi_m_wdata),
    .l2_3_targ_ht_wr_W_Last(o_l2_3_targ_ht_axi_m_wlast),
    .l2_3_targ_ht_wr_W_Ready(i_l2_3_targ_ht_axi_m_wready),
    .l2_3_targ_ht_wr_W_Strb(o_l2_3_targ_ht_axi_m_wstrb),
    .l2_3_targ_ht_wr_W_Valid(o_l2_3_targ_ht_axi_m_wvalid),
    .l2_3_targ_syscfg_PAddr(o_l2_3_targ_syscfg_apb_m_paddr),
    .l2_3_targ_syscfg_PEnable(o_l2_3_targ_syscfg_apb_m_penable),
    .l2_3_targ_syscfg_PProt(o_l2_3_targ_syscfg_apb_m_pprot),
    .l2_3_targ_syscfg_PRData(i_l2_3_targ_syscfg_apb_m_prdata),
    .l2_3_targ_syscfg_PReady(i_l2_3_targ_syscfg_apb_m_pready),
    .l2_3_targ_syscfg_PSel(o_l2_3_targ_syscfg_apb_m_psel),
    .l2_3_targ_syscfg_PSlvErr(i_l2_3_targ_syscfg_apb_m_pslverr),
    .l2_3_targ_syscfg_PStrb(o_l2_3_targ_syscfg_apb_m_pstrb),
    .l2_3_targ_syscfg_PWData(o_l2_3_targ_syscfg_apb_m_pwdata),
    .l2_3_targ_syscfg_PWrite(o_l2_3_targ_syscfg_apb_m_pwrite),
    .l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .noc_clk(i_noc_clk),
    .noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
);

endmodule
