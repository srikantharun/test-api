// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: Manuel Oliveira <manuel.oliveira@axelera.ai>


/// Package used by Read-Only monitor
///
package ro_monitor_pkg;

endpackage
