
typedef struct {
  bit [1:0]            access_type;
  bit [1:0]rd_wr;
  bit [31:0]           reg_addr;
  bit [31:0]           value;
} phy_init_value_t;

const phy_init_value_t phy_init_snps_data_details_pre[] = '{

'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10ff8, value: 'h0},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10ffc, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10b84, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10000, value: 'h3080808},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10010, value: 'h101},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10100, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10104, value: 'h5},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10108, value: 'h5},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10118, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20001},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10184, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h1018c, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10200, value: 'h3b7},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10220, value: 'h1f000301},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10224, value: 'h18},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10288, value: 'h2},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10300, value: 'h5b005b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10308, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10380, value: 'ha901a014},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10384, value: 'h80002000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10390, value: 'h83c0810},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10394, value: 'h3000041e},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10400, value: 'h2000030},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10500, value: 'h110111},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10508, value: 'h60008000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10510, value: 'h10005},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10518, value: 'h1000001},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10600, value: 'h643f5980},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10648, value: 'h600},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h1064c, value: 'h2037274},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10658, value: 'h89bbb8cf},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10660, value: 'hb7},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10984, value: 'h67},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c90, value: 'hc00b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c94, value: 'h3},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10cb0, value: 'h11},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10d00, value: 'h40030008},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10f00, value: 'h80208200},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h20004, value: 'hf00000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h20008, value: 'h2000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h20094, value: 'h2100500},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h20098, value: 'h66d04d7},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h2009c, value: 'h1110b06},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h200a0, value: 'h7607c9},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h200e0, value: 'h10105b10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h200f0, value: 'h466416f5},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h200f8, value: 'h73de8765},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h0, value: 'h280c3622},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h4, value: 'h7100830},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h8, value: 'h9131317},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hc, value: 'hc232f},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10, value: 'hf04030f},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h14, value: 'h2040c09},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h18, value: 'h12},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h1c, value: 'h3},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h24, value: 'h20310},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30, value: 'h30000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h34, value: 'hc100002},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h38, value: 'h390136},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h44, value: 'h780050},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h5c, value: 'h9d0009},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h60, value: 'h11180e},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h64, value: 'h2806},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h78, value: 'h1b151a},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h500, value: 'h510},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h504, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h508, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h50c, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h580, value: 'h33f021f},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h584, value: 'h80303},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h588, value: 'h183f1f},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h590, value: 'h200c0411},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h594, value: 'h410000f},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h598, value: 'h117},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h5a0, value: 'h20202},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h5a4, value: 'h201},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h5a8, value: 'h190000d},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h5ac, value: 'h5000a},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h5b4, value: 'h48000007},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h5b8, value: 'h147},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h600, value: 'hc03f0c34},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h604, value: 'h1300098},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h608, value: 'h6480000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h60c, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h650, value: 'hd0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h800, value: 'h1804d6},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h804, value: 'h280006d},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'ha80, value: 'h560},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hb00, value: 'hdb7fa538},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hb04, value: 'h1024100a},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hb08, value: 'h833},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hb80, value: 'hd000000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hc00, value: 'h18},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hc88, value: 'hf000000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hd00, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hd04, value: 'hb07},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hd08, value: 'h1302},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hd0c, value: 'h2990017},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hd30, value: 'h1efd6c},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hd34, value: 'h2100a159},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'hd80, value: 'h2},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h100500, value: 'h510},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h100504, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h100508, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10050c, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h200500, value: 'h510},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h200504, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h200508, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h20050c, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h300500, value: 'h510},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h300504, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h300508, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30050c, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30004, value: 'h19},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h3000c, value: 'h3f0903},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30010, value: 'h101},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30014, value: 'h1f030303},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30018, value: 'h3030300},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h3001c, value: 'h1f080808},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30020, value: 'h8080808},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30024, value: 'h8080808},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30028, value: 'h8080808},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h3002c, value: 'h808},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h30030, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10b84, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h20090, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10208, value: 'h1}
 };

const phy_init_value_t phy_init_snps_data_details[] = '{
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20001},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10100, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10510, value: 'h10004},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10c84, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10510, value: 'h10014},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10c84, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10208, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040088, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041088, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10141c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10151c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b1c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c1c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h11141c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h11151c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h111b1c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h111c1c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h12141c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h12151c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h121b1c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h121c1c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h13141c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h13151c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h131b1c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h131c1c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1010014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1011014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1012014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1013014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1014014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1015014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1017014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1018014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1019014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10b0c20, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10b0008, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0118, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f011c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0120, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0124, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1118, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f111c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1120, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1124, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1128, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f012c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f112c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2118, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f211c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2120, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2124, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3118, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f311c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3120, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3124, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3128, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f212c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f312c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4118, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f411c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4120, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4124, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5118, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f511c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5120, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5124, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5128, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f412c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f512c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6118, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f611c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6120, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6124, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7118, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f711c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7120, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7124, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7128, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f612c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f712c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040080, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041080, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1010014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1011014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1012014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1013014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1014014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1015014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1017014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1018014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1019014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c014, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10b0c20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10b0008, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0118, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f011c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0120, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0124, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1118, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f111c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1120, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1124, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1128, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f012c, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f112c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2118, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f211c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2120, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2124, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3118, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f311c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3120, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3124, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3128, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f212c, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f312c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4118, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f411c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4120, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4124, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5118, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f511c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5120, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5124, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5128, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f412c, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f512c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6118, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f611c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6120, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6124, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7118, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f711c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7120, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7124, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7128, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f612c, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f712c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1030294, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102025c, value: 'h7ff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102125c, value: 'h7ff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102225c, value: 'h7ff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102325c, value: 'h7ff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0c0c, value: 'h9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10b0c08, value: 'h26},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0c04, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0c3c, value: 'h1d},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10402b8, value: 'h1880},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10402b4, value: 'h1880},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10402b0, value: 'h1880},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10412b8, value: 'h1880},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10412b4, value: 'h1880},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10412b0, value: 'h1880},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d0218, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h108046c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102028c, value: 'h833},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102128c, value: 'h83f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102228c, value: 'h833},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102328c, value: 'h83f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d03c0, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d03c4, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d03c8, value: 'h7},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d03cc, value: 'h34},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1ccc, value: 'h2d},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d03d0, value: 'h5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d03dc, value: 'hf000},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1cdc, value: 'ha00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c7c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a20a4, value: 'hf},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h103001c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f01e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f11e8, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f21e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f31e8, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f41e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f51e8, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f61e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f71e8, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1011878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1012878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1013878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1014878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1015878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1016878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1018878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1019878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101d878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102387c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102487c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102587c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102687c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h104201c, value: 'hee66},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h104301c, value: 'hee66},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102201c, value: 'hee66},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102301c, value: 'hee66},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102401c, value: 'hee66},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102501c, value: 'hee66},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040280, value: 'h3fff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041280, value: 'h3fff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020224, value: 'h1fff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020228, value: 'h7ff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021224, value: 'h1fff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021228, value: 'h7ff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022224, value: 'h1fff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022228, value: 'h7ff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023224, value: 'h1fff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023228, value: 'h7ff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1030018, value: 'hf},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1030030, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0034, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1034, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2034, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3034, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4034, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5034, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6034, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7034, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h104009c, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10100fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10110fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10120fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10130fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10140fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10150fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h104109c, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10170fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10180fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10190fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a0fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b0fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c0fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h103022c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2004, value: 'h80a2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2018, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2018, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10b0ffc, value: 'h4101},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10b0c2c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1070020, value: 'h2e9a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2380, value: 'h64},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2384, value: 'h12c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2388, value: 'h7d0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a238c, value: 'h58},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2390, value: 'h14},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2394, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2398, value: 'h43},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a239c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a23a8, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a23ac, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a23b0, value: 'ha},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1030008, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1070100, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1030000, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10203ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10213ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10223ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10233ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f002c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f102c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f202c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f302c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f402c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f502c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f602c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f702c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020090, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021090, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022090, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023090, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020094, value: 'h2c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021094, value: 'h2c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022094, value: 'h2c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023094, value: 'h2c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102000c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102100c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102200c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102300c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0010, value: 'h320},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10b0c30, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200f8, value: 'h5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210f8, value: 'h5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220f8, value: 'h5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230f8, value: 'h5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h103000c, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h103002c, value: 'h1111},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020420, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021420, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022420, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023420, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080014, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h108003c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020038, value: 'h1300},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021038, value: 'h1300},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022038, value: 'h1300},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023038, value: 'h1300},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1030064, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f00b0, value: 'h33},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f10b0, value: 'h33},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f00b4, value: 'h303},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f10b4, value: 'h3333},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f20b0, value: 'h33},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f30b0, value: 'h33},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f20b4, value: 'h303},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f30b4, value: 'h3333},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f40b0, value: 'h33},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f50b0, value: 'h33},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f40b4, value: 'h303},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f50b4, value: 'h3333},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f60b0, value: 'h33},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f70b0, value: 'h33},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f60b4, value: 'h303},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f70b4, value: 'h3333},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10101c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10111c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10121c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10131c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10141c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10151c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10171c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10181c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10191c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a1c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b1c0, value: 'hff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c1c0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f00b8, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f10b8, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f00bc, value: 'h3300},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f10bc, value: 'h7700},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f20b8, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f30b8, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f20bc, value: 'h3300},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f30bc, value: 'h7700},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f40b8, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f50b8, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f40bc, value: 'h3300},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f50bc, value: 'h7700},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f60b8, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f70b8, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f60bc, value: 'h3300},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f70bc, value: 'h7700},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10101e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10111e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10121e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10131e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10141e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10151e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10171e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10181e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10191e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a1e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b1e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c1e4, value: 'h30},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0070, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1070, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2070, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3070, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4070, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5070, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6070, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7070, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10101b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10111b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10121b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10131b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10141b4, value: 'hf8},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10151b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10171b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10181b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10191b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a1b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b1b4, value: 'hf8},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c1b4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f00f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f10f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f20f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f30f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f40f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f50f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f60f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f70f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080100, value: 'h5b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080104, value: 'hf},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020294, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021294, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022294, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023294, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020824, value: 'h3232},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021824, value: 'h3232},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022824, value: 'h3232},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023824, value: 'h3232},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102083c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102183c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102283c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102383c, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1030014, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020020, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021020, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022020, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023020, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10801ac, value: 'h222},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080198, value: 'h20},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10803ac, value: 'h222},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080398, value: 'h20},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804d4, value: 'h100c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804d8, value: 'h100c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804dc, value: 'h41c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804e0, value: 'h1b20},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804e4, value: 'h1020},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804e8, value: 'h1020},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804ec, value: 'h430},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804f0, value: 'h2f34},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804f4, value: 'h1004},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804f8, value: 'h1004},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804fc, value: 'h414},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080500, value: 'h1318},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804b0, value: 'h83f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804b4, value: 'h83f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804c0, value: 'h83f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804b8, value: 'h81f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804bc, value: 'h81f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f004c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f104c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f204c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f304c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f404c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f504c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f604c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f704c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101178c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101278c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101378c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101478c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101578c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101678c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101878c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101978c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a78c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b78c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c78c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101d78c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f178c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f278c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f378c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f478c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f578c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f678c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f778c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f878c, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1011428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1012428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1013428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1014428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1015428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1016428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1018428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1019428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101d428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102202c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102302c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102402c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102502c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h104200c, value: 'h106a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h104300c, value: 'h106a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102200c, value: 'h106a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102300c, value: 'h106a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102400c, value: 'h106a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102500c, value: 'h106a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101140c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101240c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101340c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101440c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101540c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101640c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101840c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101940c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a40c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b40c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c40c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101d40c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102300c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102400c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102500c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102600c, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1010440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1011440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1012440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1013440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1014440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1015440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1017440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1018440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1019440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7440, value: 'h1f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a23a0, value: 'h13},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a23a4, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102042c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102142c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102242c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102342c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101018c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101118c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101218c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101318c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101418c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101518c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101718c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101818c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101918c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a18c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b18c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c18c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2028, value: 'h268},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a202c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2054, value: 'h268},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2058, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f018c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0190, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f021c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f118c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1190, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f121c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f218c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2190, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f221c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f318c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3190, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f321c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f418c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4190, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f421c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f518c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5190, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f521c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f618c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6190, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f621c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f718c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7190, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f721c, value: 'h68},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d0200, value: 'h7},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f00f0, value: 'h80},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f10f0, value: 'h80},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f20f0, value: 'h80},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f30f0, value: 'h80},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f40f0, value: 'h80},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f50f0, value: 'h80},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f60f0, value: 'h80},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f70f0, value: 'h80},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a205c, value: 'h53},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2060, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2064, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10403ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10413ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1070018, value: 'h3f0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020364, value: 'h9c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021364, value: 'h9c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022364, value: 'h9c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023364, value: 'h9c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102009c, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102109c, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102209c, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102309c, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040088, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041088, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040364, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040360, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040760, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040b60, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040f60, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041360, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041760, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041b60, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1042360, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1042760, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041364, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041360, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041760, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041b60, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041f60, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1042360, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1042760, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1042b60, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1043360, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1043760, value: 'h40},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020000, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021000, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022000, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023000, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080034, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200a8, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200ac, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210a8, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210ac, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220a8, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220ac, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230a8, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230ac, value: 'h200},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200a0, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200a4, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210a0, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210a4, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220a0, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220a4, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230a0, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230a4, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10201e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10201ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10205e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10205ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10209e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10209ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020de8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020dec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10215e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10215ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10219e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10219ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021de8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021dec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10215e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10215ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10219e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10219ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021de8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021dec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10225e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10225ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10229e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10229ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022de8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022dec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10225e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10225ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10229e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10229ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022de8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022dec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10235e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10235ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10239e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10239ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023de8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023dec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10241e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10241ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10235e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10235ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10239e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10239ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023de8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023dec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10241e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10241ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10245e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10245ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10249e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10249ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024de8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024dec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10251e8, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10251ec, value: 'hed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10201e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10201e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10205e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10205e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10209e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10209e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020de0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020de4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10215e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10215e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10219e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10219e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021de0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021de4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10215e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10215e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10219e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10219e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021de0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021de4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10225e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10225e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10229e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10229e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022de0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022de4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10225e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10225e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10229e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10229e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022de0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022de4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10235e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10235e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10239e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10239e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023de0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023de4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10241e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10241e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10235e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10235e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10239e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10239e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023de0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023de4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10241e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10241e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10245e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10245e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10249e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10249e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024de0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024de4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10251e0, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10251e4, value: 'h3b9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020080, value: 'h319},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020084, value: 'h319},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021080, value: 'h319},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021084, value: 'h319},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022080, value: 'h319},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022084, value: 'h319},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023080, value: 'h319},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023084, value: 'h319},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102004c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020440, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020444, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020448, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102044c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020840, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020844, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020848, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102084c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020c40, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020c44, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020c48, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020c4c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102104c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021440, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021444, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021448, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102144c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021840, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021844, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021848, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102184c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021c40, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021c44, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021c48, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021c4c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102204c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102104c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021440, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021444, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021448, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102144c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021840, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021844, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021848, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102184c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021c40, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021c44, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021c48, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021c4c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102204c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022440, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022444, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022448, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102244c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022840, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022844, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022848, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102284c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022c40, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022c44, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022c48, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022c4c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102304c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102204c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022440, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022444, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022448, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102244c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022840, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022844, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022848, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102284c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022c40, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022c44, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022c48, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022c4c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102304c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023440, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023444, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023448, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102344c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023840, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023844, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023848, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102384c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023c40, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023c44, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023c48, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023c4c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102404c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102304c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023440, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023444, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023448, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102344c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023840, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023844, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023848, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102384c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023c40, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023c44, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023c48, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023c4c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102404c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024440, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024444, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024448, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102444c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024840, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024844, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024848, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102484c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024c40, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024c44, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024c48, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1024c4c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1025040, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1025044, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1025048, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102504c, value: 'h12b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020030, value: 'hcc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020034, value: 'hcc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020050, value: 'h198},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020054, value: 'h198},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021030, value: 'hcc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021034, value: 'hcc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021050, value: 'h198},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021054, value: 'h198},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022030, value: 'hcc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022034, value: 'hcc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022050, value: 'h198},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022054, value: 'h198},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023030, value: 'hcc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023034, value: 'hcc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023050, value: 'h198},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023054, value: 'h198},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10801dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10301c4, value: 'h66},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101018c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101118c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101218c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101318c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101418c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101518c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101718c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101818c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101918c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101a18c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101b18c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h101c18c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f018c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0190, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f021c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f118c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1190, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f121c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f218c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2190, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f221c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f318c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3190, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f321c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f418c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4190, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f421c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f518c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5190, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f521c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f618c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6190, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f621c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f718c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7190, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f721c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2028, value: 'h262},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a202c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2054, value: 'h262},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2058, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102057c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102157c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102257c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102357c, value: 'h62},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1070024, value: 'h10},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020a80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020a84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020a88, value: 'ha},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020a8c, value: 'h3e},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020a90, value: 'h72},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021a80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021a84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021a88, value: 'ha},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021a8c, value: 'h3e},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021a90, value: 'h72},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022a80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022a84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022a88, value: 'ha},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022a8c, value: 'h3e},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022a90, value: 'h72},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023a80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023a84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023a88, value: 'ha},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023a8c, value: 'h3e},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023a90, value: 'h72},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020ab4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021ab4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022ab4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023ab4, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1020abc, value: 'h4c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1021abc, value: 'h4c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1022abc, value: 'h4c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1023abc, value: 'h4c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a201c, value: 'h9701},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2020, value: 'hb681},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10200fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10210fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10220fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10230fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0c40, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0c44, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1070020, value: 'h2d56},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1070018, value: 'h3f0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10201f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10211f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10221f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10231f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080504, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102009c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102109c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102209c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102309c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102083c, value: 'h8},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102183c, value: 'h8},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102283c, value: 'h8},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h102383c, value: 'h8},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f00fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f0234, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f10fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f1234, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f20fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f2234, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f30fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f3234, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f40fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f4234, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f50fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f5234, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f60fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f6234, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f70fc, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10f7234, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a240c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10801c8, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a2038, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10801cc, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a203c, value: 'h3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e0000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e039c, value: 'h600},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080628, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080c90, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080c94, value: 'h19},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080c98, value: 'h3c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080c9c, value: 'h5f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ca0, value: 'h77},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ca4, value: 'h9a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ca8, value: 'hbd},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cac, value: 'hd5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cb0, value: 'hf8},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cb4, value: 'h11b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cb8, value: 'h133},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cbc, value: 'h156},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cc0, value: 'h179},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cc4, value: 'h17d},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cc8, value: 'h17f},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ccc, value: 'h183},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cd0, value: 'h185},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cd4, value: 'h186},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cdc, value: 'h187},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ce0, value: 'h189},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ce8, value: 'h18a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cec, value: 'h1a3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cf0, value: 'h1ad},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080cf4, value: 'h1c5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080d38, value: 'h1d5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080d3c, value: 'h1ed},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080d40, value: 'h1f6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080d44, value: 'h208},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e2c, value: 'h18},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e30, value: 'h3b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e34, value: 'h5e},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e38, value: 'h76},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e3c, value: 'h99},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e40, value: 'hbc},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e44, value: 'hd4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e48, value: 'hf7},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e4c, value: 'h11a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e50, value: 'h132},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e54, value: 'h155},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e58, value: 'h178},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e5c, value: 'h17c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e60, value: 'h17e},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e64, value: 'h182},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e68, value: 'h184},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e6c, value: 'h185},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e70, value: 'h186},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e78, value: 'h188},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e7c, value: 'h189},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e84, value: 'h1a2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e88, value: 'h1ac},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e8c, value: 'h1c4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080e90, value: 'h1d4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ed4, value: 'h1ec},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ed8, value: 'h1f5},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080edc, value: 'h207},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080ee0, value: 'h218},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080800, value: 'h38c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080808, value: 'h3cd},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080810, value: 'hc0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080814, value: 'h246},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080818, value: 'h101},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h108081c, value: 'h287},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080820, value: 'h142},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080824, value: 'h2c8},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080828, value: 'h10},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080830, value: 'h13},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080838, value: 'h14},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080848, value: 'h2a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h108084c, value: 'h16},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080850, value: 'h2b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080854, value: 'h17},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080858, value: 'h2c},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h108085c, value: 'h18},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080860, value: 'h2d},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080864, value: 'h19},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080868, value: 'h11},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0070, value: 'h25a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0074, value: 'h25a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0078, value: 'h25a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a007c, value: 'h25a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0080, value: 'h28e},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0084, value: 'h25a},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0088, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a008c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0090, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0094, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a0098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a009c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a00ac, value: 'h28b},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c20, value: 'h7ffde000},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080514, value: 'h2},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1180514, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1280514, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1380514, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e039c, value: 'h400},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d0004, value: 'h5821},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c30, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c34, value: 'hfe},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c38, value: 'hffff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c3c, value: 'hf040},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c40, value: 'hf040},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c50, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c54, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c58, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c5c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c64, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c68, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10a1c6c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10803c0, value: 'hb6d},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10801f8, value: 'hc3},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10807bc, value: 'h7fff},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1040298, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1041298, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10806a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10804d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080508, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080510, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d0200, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e0000, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e0000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d0200, value: 'h7},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h103001c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040088, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041088, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10141c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10151c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h11141c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h11151c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h111b1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h111c1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h12141c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h12151c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h121b1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h121c1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h13141c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h13151c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h131b1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h131c1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10b0008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1030294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102025c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102125c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102225c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102325c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10c0c0c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10b0c08, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10c0c04, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10c0c3c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10402b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10402b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10402b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10412b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10412b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10412b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d0218, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h108046c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102028c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102128c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102228c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102328c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d03c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d03c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d03c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d03cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1ccc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d03d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d03dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1cdc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c7c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a20a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1011878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1012878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1013878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1014878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1015878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1016878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1018878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1019878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101d878, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102387c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102487c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102587c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102687c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h104201c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h104301c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102201c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102301c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102401c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102501c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020224, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020228, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021224, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021228, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022224, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022228, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023224, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023228, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1030018, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1030030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h104009c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10100fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10110fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10120fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10130fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10140fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10150fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h104109c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10170fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10180fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10190fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a0fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b0fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c0fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2018, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10b0ffc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10b0c2c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1070020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2380, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2384, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2388, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a238c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2390, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2394, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2398, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a239c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a23a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a23ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a23b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1030008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1070100, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1030000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10203ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10213ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10223ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10233ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f002c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f102c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f202c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f302c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f402c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f502c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f602c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f702c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020090, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021090, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022090, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023090, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020094, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021094, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022094, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023094, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102000c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102100c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102200c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102300c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10c0010, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10b0c30, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10200f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10210f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10220f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10230f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h103000c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h103002c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020420, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021420, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022420, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023420, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080014, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h108003c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020038, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021038, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022038, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023038, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1030064, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10101c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10111c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10121c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10131c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10171c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10181c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10191c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a1c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10101e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10111e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10121e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10131e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10141e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10151e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10171e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10181e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10191e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a1e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b1e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c1e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10101b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10111b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10121b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10131b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10141b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10151b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10171b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10181b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10191b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a1b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b1b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c1b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080100, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080104, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020824, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021824, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022824, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023824, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102083c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102183c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102283c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102383c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1030014, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10801ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080198, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10803ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080398, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804f4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080500, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f004c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f104c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f204c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f304c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f404c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f504c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f604c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f704c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101178c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101278c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101378c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101478c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101578c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101678c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101878c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101978c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a78c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b78c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c78c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101d78c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f178c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f278c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f378c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f478c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f578c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f678c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f778c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f878c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1011428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1012428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1013428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1014428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1015428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1016428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1018428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1019428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101d428, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102202c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102302c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102402c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102502c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h104200c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h104300c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102200c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102300c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102400c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102500c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101140c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101240c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101340c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101440c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101540c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101640c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101840c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101940c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a40c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b40c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c40c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101d40c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102300c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102400c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102500c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102600c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1010440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1011440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1012440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1013440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1014440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1015440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1017440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1018440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1019440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a23a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a23a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7008, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102042c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102142c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102242c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102342c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101018c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101118c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101218c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101318c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101418c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101518c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101718c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101818c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101918c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a18c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b18c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c18c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2028, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a202c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2058, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f018c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f021c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f118c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f121c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f218c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f221c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f318c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f321c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f418c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f421c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f518c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f521c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f618c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f621c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f718c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f721c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a205c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2060, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2064, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10403ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10413ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10c0c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1070018, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231f0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080504, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102009c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102109c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102209c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102309c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0234, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1234, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2234, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3234, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4234, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5234, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6234, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70fc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7234, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a240c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10801c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2038, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10801cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a203c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10e039c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080628, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080c90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080c94, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080c98, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080c9c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ca0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ca4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ca8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cb0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cb4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cb8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cc0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cc4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cc8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ccc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cd0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cd4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cdc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ce0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ce8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cf0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080cf4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080d38, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080d3c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080d40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080d44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e2c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e30, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e34, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e38, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e3c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e50, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e54, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e58, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e5c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e64, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e68, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e6c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e70, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e78, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e7c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e88, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080e90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ed4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ed8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080edc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080ee0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080810, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080818, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h108081c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080820, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080824, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080828, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080830, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080838, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h108084c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080850, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080854, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080858, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h108085c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080860, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080864, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080868, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0070, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0074, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0078, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a007c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0080, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0084, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0088, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a008c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0090, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0094, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a0098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a009c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a00ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080514, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1180514, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1280514, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1380514, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d0004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c30, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c34, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c38, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c3c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c50, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c54, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c58, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c5c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c64, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c68, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a1c6c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10803c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10801f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10807bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040298, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041298, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10806a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10804d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080508, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080510, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10c0c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10c0c50, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10c0c54, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10e00c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d00c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d00cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d00d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10d00d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10202f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10206f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020af8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020ef8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10212f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10216f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021af8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021ef8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10222f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10202c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020200, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020204, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020208, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102020c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020210, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020214, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020218, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102021c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020220, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020364, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10200c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10212f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10216f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021af8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021ef8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10222f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10226f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022af8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022ef8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10232f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10212c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021200, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021204, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021208, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102120c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021210, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021214, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021218, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102121c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021220, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021364, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10210c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10222f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10226f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022af8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022ef8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10232f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10236f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023af8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023ef8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10242f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10222c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022200, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022204, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022208, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102220c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022210, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022214, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022218, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102221c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022220, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022364, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10220c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10232f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10236f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023af8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023ef8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10242f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10246f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024af8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024ef8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10252f8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10232c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023200, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023204, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023208, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102320c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023210, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023214, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023218, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102321c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023220, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023364, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10230c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f009c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f109c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f00a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f10a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f209c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f309c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f20a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f30a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f409c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f509c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f40a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f50a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7098, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f609c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f709c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f60a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f70a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10301c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040364, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040360, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040760, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040b60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1040f60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041360, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041760, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041b60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041f60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1042360, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1042760, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041364, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041360, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041760, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041b60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1041f60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1042360, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1042760, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1042b60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1042f60, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1043360, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1043760, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1011980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1011984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1011580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1011584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1012980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1012984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1012580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1012584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1013980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1013984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1013580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1013584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1014980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1014984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1014580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1014584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1015980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1015984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1015580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1015584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1018980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1018984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1018580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1018584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1019980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1019984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1019580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1019584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101a584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101b584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h101c584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020ab4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020abc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020a80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020a84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020a88, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020a8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020a90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020080, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020084, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10200a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10200a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10200a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10200ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102004c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10201bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102018c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020444, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020448, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102044c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020720, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10205bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102058c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020590, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020840, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020844, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102084c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020b20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10209bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102098c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020990, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020de0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020de4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020de8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020dec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020f20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020da0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020da4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020da8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020dac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020db0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020db4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020db8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020dbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020d80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020d84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020d8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020d90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102104c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102118c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021444, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021448, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102144c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021720, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102158c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021590, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021840, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021844, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102184c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021b20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102198c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021990, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021de0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021de4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021de8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021dec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021f20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021da0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021da4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021da8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021dac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021db0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021db4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021db8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021dbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021d80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021d84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021d8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021d90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102204c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102218c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020050, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020064, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102006c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1020088, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102008c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102057c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021ab4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021abc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021a80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021a84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021a88, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021a8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021a90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021080, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021084, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10210a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10210a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10210a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10210ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102104c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10211bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102118c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021444, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021448, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102144c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021720, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10215bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102158c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021590, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021840, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021844, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102184c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021b20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10219bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102198c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021990, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021de0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021de4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021de8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021dec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021f20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021da0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021da4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021da8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021dac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021db0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021db4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021db8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021dbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021d80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021d84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021d8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021d90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102204c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102218c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022444, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022448, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102244c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022720, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102258c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022590, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022840, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022844, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102284c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022b20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102298c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022990, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022de0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022de4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022de8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022dec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022f20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022da0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022da4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022da8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022dac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022db0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022db4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022db8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022dbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022d80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022d84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022d8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022d90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102304c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102318c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021050, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021064, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102106c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1021088, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102108c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102157c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022ab4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022abc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022a80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022a84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022a88, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022a8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022a90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022080, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022084, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10220a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10220a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10220a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10220ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102204c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10221bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102218c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022444, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022448, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102244c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022720, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10225bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102258c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022590, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022840, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022844, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102284c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022b20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10229bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102298c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022990, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022de0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022de4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022de8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022dec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022f20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022da0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022da4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022da8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022dac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022db0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022db4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022db8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022dbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022d80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022d84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022d8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022d90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102304c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102318c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023444, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023448, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102344c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023720, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102358c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023590, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023840, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023844, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102384c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023b20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102398c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023990, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023de0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023de4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023de8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023dec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023f20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023da0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023da4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023da8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023dac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023db0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023db4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023db8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023dbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023d80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023d84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023d8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023d90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102404c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102418c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022050, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022064, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102206c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1022088, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102208c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102257c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023ab4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023abc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023a80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023a84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023a88, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023a8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023a90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023080, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023084, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10230a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10230a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10230a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10230ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102304c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10231bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102318c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023444, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023448, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102344c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023720, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10235bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102358c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023590, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023840, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023844, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102384c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023b20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10239bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102398c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023990, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023de0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023de4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023de8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023dec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023f20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023da0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023da4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023da8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023dac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023db0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023db4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023db8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023dbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023d80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023d84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023d8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023d90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102404c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10241bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102418c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024440, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024444, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024448, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102444c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024720, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10245bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102458c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024590, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024840, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024844, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024848, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102484c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024b20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10249bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024980, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024984, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102498c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024990, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024de0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024de4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024de8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024dec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024c40, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024c44, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024c48, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024c4c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024f20, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024da0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024da4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024da8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024dac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024db0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024db4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024db8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024dbc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024d80, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024d84, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024d8c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1024d90, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251e8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251ec, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1025040, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1025044, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1025048, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102504c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1025320, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251a0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251a4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251a8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251ac, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251b0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251b4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251b8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10251bc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1025180, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1025184, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102518c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1025190, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023030, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023050, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023054, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023064, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102306c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1023088, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102308c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h102357c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1070024, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080034, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f01e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f11e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f03c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f13c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f03c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f13c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f03c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f13c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f03cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f13cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f13d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f03d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f13d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0804, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1804, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f080c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f180c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1810, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f02c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f12c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0300, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1300, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0340, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1340, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1380, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0284, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1284, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f02c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f12c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0304, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1304, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0344, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1344, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1384, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0290, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1290, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f02d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f12d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0310, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1310, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0350, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1350, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1390, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f02d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f12d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0314, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1314, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f0354, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1354, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1394, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1540, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2540, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1544, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2544, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f15c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f25c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f15c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f25c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1600, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2600, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f1604, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2604, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f21e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f31e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f23c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f33c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f23c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f33c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f23c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f33c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f23cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f33cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f33d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f23d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f33d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2804, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3804, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f280c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f380c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3810, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f22c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f32c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2300, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3300, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2340, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3340, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3380, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2284, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3284, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f22c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f32c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2304, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3304, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2344, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3344, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3384, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2290, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3290, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f22d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f32d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2310, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3310, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2350, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3350, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3390, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f22d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f32d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2314, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3314, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f2354, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3354, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3394, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3540, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4540, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3544, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4544, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f35c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f45c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f35c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f45c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3600, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4600, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f3604, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4604, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f41e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f51e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f43c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f53c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f43c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f53c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f43c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f53c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f43cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f53cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f53d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f43d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f53d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4804, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5804, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f480c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f580c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5810, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f42c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f52c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4300, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5300, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4340, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5340, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5380, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4284, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5284, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f42c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f52c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4304, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5304, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4344, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5344, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5384, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4290, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5290, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f42d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f52d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4310, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5310, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4350, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5350, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5390, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f42d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f52d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4314, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5314, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f4354, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5354, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5394, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5540, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6540, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5544, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6544, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f55c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f65c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f55c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f65c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5600, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6600, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f5604, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6604, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71d8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f61e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71e0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f71e4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f63c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f73c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f63c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f73c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f63c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f73c8, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f63cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f73cc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f73d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f63d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f73d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7800, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6804, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7804, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7808, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f680c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f780c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7810, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7814, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7280, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f62c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f72c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6300, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7300, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6340, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7340, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7380, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6284, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7284, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f62c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f72c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6304, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7304, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6344, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7344, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7384, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6290, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7290, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f62d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f72d0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6310, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7310, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6350, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7350, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7390, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7294, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f62d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f72d4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6314, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7314, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f6354, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7354, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7394, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7540, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f8540, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7544, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f8544, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f8580, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f8584, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f75c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f85c0, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f75c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f85c4, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7600, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f8600, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f7604, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10f8604, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a201c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10a2020, value: 'h0},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10801dc, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h103001c, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10c0004, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10d0200, value: 'h4},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e0000, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e0000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1030014, value: 'h6},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h108019c, value: 'h9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h108039c, value: 'h9},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080100, value: 'h9},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080100, value: 'h5e},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1180100, value: 'h5e},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1180100, value: 'he},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1280100, value: 'he},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1280100, value: 'he},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1380100, value: 'he},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1380100, value: 'he},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080198, value: 'he},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080198, value: 'hb20},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1080398, value: 'hb20},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1080398, value: 'hb20},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10801ac, value: 'hb20},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10801ac, value: 'hb22},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h10803ac, value: 'hb22},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10803ac, value: 'hb22},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1180198, value: 'hb22},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1180198, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1180398, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1180398, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h11801ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h11801ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h11803ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h11803ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1280198, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1280198, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1280398, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1280398, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h12801ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h12801ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h12803ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h12803ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1380198, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1380198, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h1380398, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h1380398, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h13801ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h13801ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h2, reg_addr: 'h13803ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h13803ac, value: 'hb00},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h108003c, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e0000, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10510, value: 'h10034},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10c84, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10510, value: 'h1},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e0000, value: 'h0},
'{access_type: 'h2, rd_wr: 'h3, reg_addr: 'h10e0000, value: 'h1}};


const phy_init_value_t phy_init_snps_data_details_post[] = '{
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10514, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10510, value: 'h10014},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10c84, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10510, value: 'h10015},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10c80, value: 'h1},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10c84, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10014, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'ha80, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'ha80, value: 'h560},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h560},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h255b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h285b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2900},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2e00},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h255b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h285b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2900},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2e00},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10518, value: 'h1000000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h1000000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h121e},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h121e},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1b0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1b0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2bb},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2bb},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h381},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h381},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'ha58},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'ha58},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'hb44},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'hb44},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'hc12},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'hc12},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'hd00},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'hd00},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'he10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'he10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'hf13},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'hf13},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1128},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1128},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1300},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1300},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1402},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1402},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1640},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1640},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1700},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1700},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h18c6},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h18c6},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1980},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1980},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1c00},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h1c00},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h255b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h255b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h285b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h285b},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2904},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2904},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2e00},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000010},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h20},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10084, value: 'h2e00},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10080, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h80000020},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10518, value: 'h1000001},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10208, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20001},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20001},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10100, value: 'h1},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'ha80, value: 'h560},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10000, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10000, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h200e0, value: 'h10105b10},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10180, value: 'h20000},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10184, value: 'h0},
'{access_type: 'h1, rd_wr: 'h3, reg_addr: 'h10100, value: 'h5},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10090, value: 'h5},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10b88, value: 'h5},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10b88, value: 'h5},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10b88, value: 'h5},
'{access_type: 'h1, rd_wr: 'h2, reg_addr: 'h10b88, value: 'h5}
} ;
