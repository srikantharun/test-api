
// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description:
// Owner: Axelera (Axelera@axelera.ai)

`ifndef EUROPA_SV
`define EUROPA_SV

module europa

  import aic_common_pkg::*;
  import aic_ls_pkg::*;
  import apu_interrupt_map_pkg::*;
  import apu_pkg::*;
  import axe_tcl_sram_pkg::*;
  import axi_pkg::*;
  import chip_pkg::*;
  import dcd_pkg::*;
  import ddr_west_clock_gen_pkg::*;
  import dmc_pkg::*;
  import emmc_pkg::*;
  import l2_p_pkg::*;
  import lpddr_pkg::*;
  import pcie_pkg::*;
  import pve_pkg::*;
  import rot_pkg::*;
  import soc_mgmt_pkg::*;
  import soc_periph_pkg::*;
  import svs_monitor_pkg::*;
  import sys_spm_pkg::*;


(
  input wire    i_ref_clk,
  output wire    o_ref_clk,
  input logic   i_ref_clk_bypass,
  input wire    i_tck,
  output logic   o_spi_clk_out,
  inout wire    io_i2c_0_clk,
  inout wire    io_i2c_1_clk,
  output logic   o_sd_emmc_clk_out,
  input wire    i_por_rst_n,
  input wire    i_trst_n,
  input logic   i_uart_rx,
  output logic   o_uart_tx,
  input logic   i_uart_cts_n,
  output logic   o_uart_rts_n,
  output logic  [3:0] o_spi_ss_n,
  inout wire   [3:0] io_spi_sd,
  inout wire    io_i2c_0_data,
  inout wire    io_i2c_1_data,
  inout wire   [15:0] io_gpio,
  inout wire    io_sd_emmc_cmd,
  inout wire   [7:0] io_sd_emmc_data,
  inout wire    io_emmc_rebar,
  input logic   i_emmc_lpbk_dqs,
  input logic   i_sd_emmc_strobe,
  output logic   o_emmc_reset,
  output logic   o_emmc_power,
  input logic   i_sd_emmc_detect,
  input logic   i_sd_emmc_wp,
  output logic   o_sd_emmc_pu_pd,
  output logic  [15:0] o_observability,
  output logic   o_thermal_warning_n,
  output logic   o_thermal_shutdown_n,
  input logic   i_thermal_throttle,
  input logic   i_throttle,
  input logic  [2:0] i_boot_mode,
  input logic   i_tms,
  input logic   i_td_in,
  output logic   o_td_out,
  input wire    i_ssn_bus_0_clk,
  input wire    i_ssn_bus_1_clk,
  inout wire   [44:0] io_dft_test,
  inout wire    io_efuse_vqps,
  inout wire    io_efuse_vddwl,
  inout wire    io_pvt_test_out_ts,
  inout wire    io_otp_vtdo,
  inout wire    io_otp_vrefm,
  inout wire    io_otp_vpp,
  output wire    o_lpddr_ppp_0_bp_memreset_l,
  output wire    o_lpddr_ppp_1_bp_memreset_l,
  output wire    o_lpddr_ppp_2_bp_memreset_l,
  output wire    o_lpddr_ppp_3_bp_memreset_l,
  inout wire   [19:0] io_lpddr_ppp_0_bp_a,
  inout wire   [19:0] io_lpddr_ppp_1_bp_a,
  inout wire   [19:0] io_lpddr_ppp_2_bp_a,
  inout wire   [19:0] io_lpddr_ppp_3_bp_a,
  inout wire    io_lpddr_ppp_0_bp_ato,
  inout wire    io_lpddr_ppp_1_bp_ato,
  inout wire    io_lpddr_ppp_2_bp_ato,
  inout wire    io_lpddr_ppp_3_bp_ato,
  inout wire    io_lpddr_ppp_0_bp_ato_pll,
  inout wire    io_lpddr_ppp_1_bp_ato_pll,
  inout wire    io_lpddr_ppp_2_bp_ato_pll,
  inout wire    io_lpddr_ppp_3_bp_ato_pll,
  inout wire   [12:0] io_lpddr_ppp_0_bp_b0_d,
  inout wire   [12:0] io_lpddr_ppp_1_bp_b0_d,
  inout wire   [12:0] io_lpddr_ppp_2_bp_b0_d,
  inout wire   [12:0] io_lpddr_ppp_3_bp_b0_d,
  inout wire   [12:0] io_lpddr_ppp_0_bp_b1_d,
  inout wire   [12:0] io_lpddr_ppp_1_bp_b1_d,
  inout wire   [12:0] io_lpddr_ppp_2_bp_b1_d,
  inout wire   [12:0] io_lpddr_ppp_3_bp_b1_d,
  inout wire   [12:0] io_lpddr_ppp_0_bp_b2_d,
  inout wire   [12:0] io_lpddr_ppp_1_bp_b2_d,
  inout wire   [12:0] io_lpddr_ppp_2_bp_b2_d,
  inout wire   [12:0] io_lpddr_ppp_3_bp_b2_d,
  inout wire   [12:0] io_lpddr_ppp_0_bp_b3_d,
  inout wire   [12:0] io_lpddr_ppp_1_bp_b3_d,
  inout wire   [12:0] io_lpddr_ppp_2_bp_b3_d,
  inout wire   [12:0] io_lpddr_ppp_3_bp_b3_d,
  inout wire    io_lpddr_ppp_0_bp_ck0_c,
  inout wire    io_lpddr_ppp_1_bp_ck0_c,
  inout wire    io_lpddr_ppp_2_bp_ck0_c,
  inout wire    io_lpddr_ppp_3_bp_ck0_c,
  inout wire    io_lpddr_ppp_0_bp_ck0_t,
  inout wire    io_lpddr_ppp_1_bp_ck0_t,
  inout wire    io_lpddr_ppp_2_bp_ck0_t,
  inout wire    io_lpddr_ppp_3_bp_ck0_t,
  inout wire    io_lpddr_ppp_0_bp_ck1_c,
  inout wire    io_lpddr_ppp_1_bp_ck1_c,
  inout wire    io_lpddr_ppp_2_bp_ck1_c,
  inout wire    io_lpddr_ppp_3_bp_ck1_c,
  inout wire    io_lpddr_ppp_0_bp_ck1_t,
  inout wire    io_lpddr_ppp_1_bp_ck1_t,
  inout wire    io_lpddr_ppp_2_bp_ck1_t,
  inout wire    io_lpddr_ppp_3_bp_ck1_t,
  inout wire    io_lpddr_ppp_0_bp_zn,
  inout wire    io_lpddr_ppp_1_bp_zn,
  inout wire    io_lpddr_ppp_2_bp_zn,
  inout wire    io_lpddr_ppp_3_bp_zn,
  output wire    o_lpddr_graph_0_bp_memreset_l,
  output wire    o_lpddr_graph_1_bp_memreset_l,
  output wire    o_lpddr_graph_2_bp_memreset_l,
  output wire    o_lpddr_graph_3_bp_memreset_l,
  inout wire   [19:0] io_lpddr_graph_0_bp_a,
  inout wire   [19:0] io_lpddr_graph_1_bp_a,
  inout wire   [19:0] io_lpddr_graph_2_bp_a,
  inout wire   [19:0] io_lpddr_graph_3_bp_a,
  inout wire    io_lpddr_graph_0_bp_ato,
  inout wire    io_lpddr_graph_1_bp_ato,
  inout wire    io_lpddr_graph_2_bp_ato,
  inout wire    io_lpddr_graph_3_bp_ato,
  inout wire    io_lpddr_graph_0_bp_ato_pll,
  inout wire    io_lpddr_graph_1_bp_ato_pll,
  inout wire    io_lpddr_graph_2_bp_ato_pll,
  inout wire    io_lpddr_graph_3_bp_ato_pll,
  inout wire   [12:0] io_lpddr_graph_0_bp_b0_d,
  inout wire   [12:0] io_lpddr_graph_1_bp_b0_d,
  inout wire   [12:0] io_lpddr_graph_2_bp_b0_d,
  inout wire   [12:0] io_lpddr_graph_3_bp_b0_d,
  inout wire   [12:0] io_lpddr_graph_0_bp_b1_d,
  inout wire   [12:0] io_lpddr_graph_1_bp_b1_d,
  inout wire   [12:0] io_lpddr_graph_2_bp_b1_d,
  inout wire   [12:0] io_lpddr_graph_3_bp_b1_d,
  inout wire   [12:0] io_lpddr_graph_0_bp_b2_d,
  inout wire   [12:0] io_lpddr_graph_1_bp_b2_d,
  inout wire   [12:0] io_lpddr_graph_2_bp_b2_d,
  inout wire   [12:0] io_lpddr_graph_3_bp_b2_d,
  inout wire   [12:0] io_lpddr_graph_0_bp_b3_d,
  inout wire   [12:0] io_lpddr_graph_1_bp_b3_d,
  inout wire   [12:0] io_lpddr_graph_2_bp_b3_d,
  inout wire   [12:0] io_lpddr_graph_3_bp_b3_d,
  inout wire    io_lpddr_graph_0_bp_ck0_c,
  inout wire    io_lpddr_graph_1_bp_ck0_c,
  inout wire    io_lpddr_graph_2_bp_ck0_c,
  inout wire    io_lpddr_graph_3_bp_ck0_c,
  inout wire    io_lpddr_graph_0_bp_ck0_t,
  inout wire    io_lpddr_graph_1_bp_ck0_t,
  inout wire    io_lpddr_graph_2_bp_ck0_t,
  inout wire    io_lpddr_graph_3_bp_ck0_t,
  inout wire    io_lpddr_graph_0_bp_ck1_c,
  inout wire    io_lpddr_graph_1_bp_ck1_c,
  inout wire    io_lpddr_graph_2_bp_ck1_c,
  inout wire    io_lpddr_graph_3_bp_ck1_c,
  inout wire    io_lpddr_graph_0_bp_ck1_t,
  inout wire    io_lpddr_graph_1_bp_ck1_t,
  inout wire    io_lpddr_graph_2_bp_ck1_t,
  inout wire    io_lpddr_graph_3_bp_ck1_t,
  inout wire    io_lpddr_graph_0_bp_zn,
  inout wire    io_lpddr_graph_1_bp_zn,
  inout wire    io_lpddr_graph_2_bp_zn,
  inout wire    io_lpddr_graph_3_bp_zn,
  inout wire    io_pcie_resref,
  input wire    i_ref_pad_clk_p,
  input wire    i_ref_pad_clk_m,
  input wire    i_pcie_perst_n,
  input logic   i_pcie_rxm_00,
  input logic   i_pcie_rxm_01,
  input logic   i_pcie_rxm_02,
  input logic   i_pcie_rxm_03,
  input logic   i_pcie_rxp_00,
  input logic   i_pcie_rxp_01,
  input logic   i_pcie_rxp_02,
  input logic   i_pcie_rxp_03,
  output logic   o_pcie_txm_00,
  output logic   o_pcie_txm_01,
  output logic   o_pcie_txm_02,
  output logic   o_pcie_txm_03,
  output logic   o_pcie_txp_00,
  output logic   o_pcie_txp_01,
  output logic   o_pcie_txp_02,
  output logic   o_pcie_txp_03
);


  logic  [1:0] u_aipu_to_u_europa_io__o_ref_clk_sel_freq;
  wire   u_aipu_to_u_europa_io__o_spi_clk_out;
  logic   u_aipu_to_u_europa_io__o_uart_tx;
  logic   u_aipu_to_u_europa_io__o_uart_rts_n;
  logic  [1:0] u_aipu_to_u_europa_io__o_uart_drive;
  logic   u_aipu_to_u_europa_io__o_uart_schmitt;
  logic   u_aipu_to_u_europa_io__o_uart_cts_n_pd_en;
  logic   u_aipu_to_u_europa_io__o_uart_rx_pd_en;
  logic  [3:0] u_aipu_to_u_europa_io__o_spi_ss_n;
  logic  [3:0] u_aipu_to_u_europa_io__o_spi_sd;
  logic  [3:0] u_aipu_to_u_europa_io__o_spi_sd_oe_n;
  logic  [1:0] u_aipu_to_u_europa_io__o_spi_drive;
  logic   u_aipu_to_u_europa_io__o_spi_schmitt;
  logic  [3:0] u_aipu_to_u_europa_io__o_spi_sd_pd_en;
  logic   u_aipu_to_u_europa_io__o_i2c_0_clk_oe;
  logic   u_aipu_to_u_europa_io__o_i2c_1_clk_oe;
  logic   u_aipu_to_u_europa_io__o_i2c_0_data_oe;
  logic   u_aipu_to_u_europa_io__o_i2c_1_data_oe;
  logic  [1:0] u_aipu_to_u_europa_io__o_i2c_drive;
  logic   u_aipu_to_u_europa_io__o_i2c_schmitt;
  logic  [15:0] u_aipu_to_u_europa_io__o_gpio;
  logic  [15:0] u_aipu_to_u_europa_io__o_gpio_oe;
  logic  [1:0] u_aipu_to_u_europa_io__o_gpio_drive;
  logic   u_aipu_to_u_europa_io__o_gpio_schmitt;
  logic  [15:0] u_aipu_to_u_europa_io__o_gpio_pd_en;
  logic   u_aipu_to_u_europa_io__o_mem_webar_opad;
  logic   u_aipu_to_u_europa_io__o_mem_webar_oepad;
  logic   u_aipu_to_u_europa_io__o_mem_ale_opad;
  logic   u_aipu_to_u_europa_io__o_mem_ale_oepad;
  logic   u_aipu_to_u_europa_io__o_mem_ctrl_0_iepad;
  logic   u_aipu_to_u_europa_io__o_mem_ctrl_1_oepad;
  logic   u_aipu_to_u_europa_io__o_mem_ctrl_1_opad;
  logic   u_aipu_to_u_europa_io__o_mem_dqs_iepad;
  logic   u_aipu_to_u_europa_io__o_mem_rstbar_oepad;
  logic   u_aipu_to_u_europa_io__o_mem_rstbar_opad;
  logic   u_aipu_to_u_europa_io__o_mem_wpbar_iepad;
  logic   u_aipu_to_u_europa_io__o_mem_lpbk_dqs_iepad;
  logic   u_aipu_to_u_europa_io__o_mem_rebar_oepad;
  logic   u_aipu_to_u_europa_io__o_mem_rebar_iepad;
  logic   u_aipu_to_u_europa_io__o_mem_rebar_opad;
  logic   u_aipu_to_u_europa_io__o_mem_cmd_oepad;
  logic   u_aipu_to_u_europa_io__o_mem_cmd_iepad;
  logic   u_aipu_to_u_europa_io__o_mem_cmd_opad;
  logic  [7:0] u_aipu_to_u_europa_io__o_mem_data_opad;
  logic  [7:0] u_aipu_to_u_europa_io__o_mem_data_oepad;
  logic  [7:0] u_aipu_to_u_europa_io__o_mem_data_iepad;
  logic  [15:0] u_aipu_to_u_europa_io__o_observability;
  logic   u_aipu_to_u_europa_io__o_thermal_warning_n;
  logic   u_aipu_to_u_europa_io__o_thermal_shutdown_n;
  logic  [2:0] u_aipu_to_u_europa_io__o_bootmode_pull_en;
  logic   u_aipu_to_u_europa_io__o_td;
  logic  [1:0] u_aipu_to_u_europa_io__o_dft_drive;
  logic   u_aipu_to_u_europa_io__o_dft_schmitt;
  logic  [44:0] u_aipu_to_u_europa_io__o_dft_test;
  logic  [44:0] u_aipu_to_u_europa_io__o_dft_test_oe;
  logic  [2:0] u_aipu_to_u_europa_io__o_emmc_drive;
  logic   u_aipu_to_u_europa_io__o_emmc_schmitt;
  logic  [1:0] u_aipu_to_u_europa_io__o_jtag_drive;
  logic  [1:0] u_aipu_to_u_europa_io__o_obs_drive;
  logic   u_aipu_to_u_europa_io__o_clk_schmitt;
  logic   u_aipu_to_u_europa_io__o_rst_schmitt;
  logic   u_europa_io_to_u_aipu__o_ref_clk;
  logic   u_europa_io_to_u_aipu__o_tck;
  logic   u_europa_io_to_u_aipu__o_ssn_bus_0_clk;
  logic   u_europa_io_to_u_aipu__o_ssn_bus_1_clk;
  logic   u_europa_io_to_u_aipu__o_por_rst_n;
  logic   u_europa_io_to_u_aipu__o_trst_n;
  logic   u_europa_io_to_u_aipu__o_uart_rx;
  logic   u_europa_io_to_u_aipu__o_uart_cts_n;
  logic  [3:0] u_europa_io_to_u_aipu__o_spi_sd;
  logic   u_europa_io_to_u_aipu__o_i2c_0_clk;
  logic   u_europa_io_to_u_aipu__o_i2c_1_clk;
  logic   u_europa_io_to_u_aipu__o_i2c_0_data;
  logic   u_europa_io_to_u_aipu__o_i2c_1_data;
  logic  [15:0] u_europa_io_to_u_aipu__o_gpio;
  logic   u_europa_io_to_u_aipu__o_sd_emmc_detect;
  logic   u_europa_io_to_u_aipu__o_sd_emmc_strobe;
  logic   u_europa_io_to_u_aipu__o_sd_emmc_wp;
  logic   u_europa_io_to_u_aipu__o_emmc_lpbk_dqs;
  logic   u_europa_io_to_u_aipu__o_emmc_rebar;
  logic   u_europa_io_to_u_aipu__o_sd_emmc_cmd;
  logic  [7:0] u_europa_io_to_u_aipu__o_sd_emmc_data;
  logic   u_europa_io_to_u_aipu__o_thermal_throttle;
  logic   u_europa_io_to_u_aipu__o_throttle;
  logic  [2:0] u_europa_io_to_u_aipu__o_boot_mode;
  logic   u_europa_io_to_u_aipu__o_tms;
  logic   u_europa_io_to_u_aipu__o_td;
  logic  [44:0] u_europa_io_to_u_aipu__o_dft_test;
  logic   u_europa_io_to_u_aipu__o_pcie_perst_n;



aipu u_aipu (
  .i_ref_clk (u_europa_io_to_u_aipu__o_ref_clk),
  .i_tck (u_europa_io_to_u_aipu__o_tck),
  .o_spi_clk_out (u_aipu_to_u_europa_io__o_spi_clk_out),
  .i_ssn_bus_0_clk (u_europa_io_to_u_aipu__o_ssn_bus_0_clk),
  .i_ssn_bus_1_clk (u_europa_io_to_u_aipu__o_ssn_bus_1_clk),
  .i_por_rst_n (u_europa_io_to_u_aipu__o_por_rst_n),
  .i_trst_n (u_europa_io_to_u_aipu__o_trst_n),
  .i_uart_rx (u_europa_io_to_u_aipu__o_uart_rx),
  .o_uart_tx (u_aipu_to_u_europa_io__o_uart_tx),
  .i_uart_cts_n (u_europa_io_to_u_aipu__o_uart_cts_n),
  .o_uart_rts_n (u_aipu_to_u_europa_io__o_uart_rts_n),
  .o_spi_ss_n (u_aipu_to_u_europa_io__o_spi_ss_n),
  .i_spi_sd (u_europa_io_to_u_aipu__o_spi_sd),
  .o_spi_sd (u_aipu_to_u_europa_io__o_spi_sd),
  .o_spi_sd_oe_n (u_aipu_to_u_europa_io__o_spi_sd_oe_n),
  .i_i2c_0_clk (u_europa_io_to_u_aipu__o_i2c_0_clk),
  .o_i2c_0_clk_oe (u_aipu_to_u_europa_io__o_i2c_0_clk_oe),
  .i_i2c_1_clk (u_europa_io_to_u_aipu__o_i2c_1_clk),
  .o_i2c_1_clk_oe (u_aipu_to_u_europa_io__o_i2c_1_clk_oe),
  .i_i2c_0_data (u_europa_io_to_u_aipu__o_i2c_0_data),
  .o_i2c_0_data_oe (u_aipu_to_u_europa_io__o_i2c_0_data_oe),
  .i_i2c_1_data (u_europa_io_to_u_aipu__o_i2c_1_data),
  .o_i2c_1_data_oe (u_aipu_to_u_europa_io__o_i2c_1_data_oe),
  .i_gpio (u_europa_io_to_u_aipu__o_gpio),
  .o_gpio (u_aipu_to_u_europa_io__o_gpio),
  .o_gpio_oe (u_aipu_to_u_europa_io__o_gpio_oe),
  .o_mem_ale_oepad (u_aipu_to_u_europa_io__o_mem_ale_oepad),
  .o_mem_ale_opad (u_aipu_to_u_europa_io__o_mem_ale_opad),
  .i_mem_cmd_ipad (u_europa_io_to_u_aipu__o_sd_emmc_cmd),
  .o_mem_cmd_oepad (u_aipu_to_u_europa_io__o_mem_cmd_oepad),
  .o_mem_cmd_iepad (u_aipu_to_u_europa_io__o_mem_cmd_iepad),
  .o_mem_cmd_opad (u_aipu_to_u_europa_io__o_mem_cmd_opad),
  .o_mem_ctrl_0_iepad (u_aipu_to_u_europa_io__o_mem_ctrl_0_iepad),
  .i_mem_ctrl_0_ipad (u_europa_io_to_u_aipu__o_sd_emmc_detect),
  .o_mem_ctrl_1_oepad (u_aipu_to_u_europa_io__o_mem_ctrl_1_oepad),
  .o_mem_ctrl_1_opad (u_aipu_to_u_europa_io__o_mem_ctrl_1_opad),
  .o_mem_rstbar_oepad (u_aipu_to_u_europa_io__o_mem_rstbar_oepad),
  .o_mem_rstbar_opad (u_aipu_to_u_europa_io__o_mem_rstbar_opad),
  .i_mem_lpbk_dqs_ipad (u_europa_io_to_u_aipu__o_emmc_lpbk_dqs),
  .o_mem_lpbk_dqs_iepad (u_aipu_to_u_europa_io__o_mem_lpbk_dqs_iepad),
  .i_mem_dqs_ipad (u_europa_io_to_u_aipu__o_sd_emmc_strobe),
  .o_mem_dqs_iepad (u_aipu_to_u_europa_io__o_mem_dqs_iepad),
  .o_mem_rebar_oepad (u_aipu_to_u_europa_io__o_mem_rebar_oepad),
  .o_mem_rebar_iepad (u_aipu_to_u_europa_io__o_mem_rebar_iepad),
  .o_mem_rebar_opad (u_aipu_to_u_europa_io__o_mem_rebar_opad),
  .i_mem_rebar_ipad (u_europa_io_to_u_aipu__o_emmc_rebar),
  .i_mem_data_ipad (u_europa_io_to_u_aipu__o_sd_emmc_data),
  .o_mem_data_oepad (u_aipu_to_u_europa_io__o_mem_data_oepad),
  .o_mem_data_iepad (u_aipu_to_u_europa_io__o_mem_data_iepad),
  .o_mem_data_opad (u_aipu_to_u_europa_io__o_mem_data_opad),
  .o_mem_webar_oepad (u_aipu_to_u_europa_io__o_mem_webar_oepad),
  .o_mem_webar_opad (u_aipu_to_u_europa_io__o_mem_webar_opad),
  .o_mem_wpbar_iepad (u_aipu_to_u_europa_io__o_mem_wpbar_iepad),
  .i_mem_wpbar_ipad (u_europa_io_to_u_aipu__o_sd_emmc_wp),
  .o_ref_clk_sel_freq (u_aipu_to_u_europa_io__o_ref_clk_sel_freq),
  .o_jtag_drive (u_aipu_to_u_europa_io__o_jtag_drive),
  .o_uart_drive (u_aipu_to_u_europa_io__o_uart_drive),
  .o_spi_drive (u_aipu_to_u_europa_io__o_spi_drive),
  .o_i2c_drive (u_aipu_to_u_europa_io__o_i2c_drive),
  .o_gpio_drive (u_aipu_to_u_europa_io__o_gpio_drive),
  .o_obs_drive (u_aipu_to_u_europa_io__o_obs_drive),
  .o_dft_drive (u_aipu_to_u_europa_io__o_dft_drive),
  .o_emmc_drive (u_aipu_to_u_europa_io__o_emmc_drive),
  .o_clk_schmitt (u_aipu_to_u_europa_io__o_clk_schmitt),
  .o_rst_schmitt (u_aipu_to_u_europa_io__o_rst_schmitt),
  .o_spi_schmitt (u_aipu_to_u_europa_io__o_spi_schmitt),
  .o_uart_schmitt (u_aipu_to_u_europa_io__o_uart_schmitt),
  .o_i2c_schmitt (u_aipu_to_u_europa_io__o_i2c_schmitt),
  .o_gpio_schmitt (u_aipu_to_u_europa_io__o_gpio_schmitt),
  .o_emmc_schmitt (u_aipu_to_u_europa_io__o_emmc_schmitt),
  .o_dft_schmitt (u_aipu_to_u_europa_io__o_dft_schmitt),
  .o_bootmode_pull_en (u_aipu_to_u_europa_io__o_bootmode_pull_en),
  .o_spi_sd_pd_en (u_aipu_to_u_europa_io__o_spi_sd_pd_en),
  .o_uart_cts_n_pd_en (u_aipu_to_u_europa_io__o_uart_cts_n_pd_en),
  .o_uart_rx_pd_en (u_aipu_to_u_europa_io__o_uart_rx_pd_en),
  .o_gpio_pd_en (u_aipu_to_u_europa_io__o_gpio_pd_en),
  .o_observability (u_aipu_to_u_europa_io__o_observability),
  .o_thermal_warning_n (u_aipu_to_u_europa_io__o_thermal_warning_n),
  .o_thermal_shutdown_n (u_aipu_to_u_europa_io__o_thermal_shutdown_n),
  .i_thermal_throttle (u_europa_io_to_u_aipu__o_thermal_throttle),
  .i_throttle (u_europa_io_to_u_aipu__o_throttle),
  .i_boot_mode (u_europa_io_to_u_aipu__o_boot_mode),
  .i_tms (u_europa_io_to_u_aipu__o_tms),
  .i_td (u_europa_io_to_u_aipu__o_td),
  .o_td (u_aipu_to_u_europa_io__o_td),
  .i_dft_test (u_europa_io_to_u_aipu__o_dft_test),
  .o_dft_test (u_aipu_to_u_europa_io__o_dft_test),
  .o_dft_test_oe (u_aipu_to_u_europa_io__o_dft_test_oe),
  .io_efuse_vqps (io_efuse_vqps),
  .io_efuse_vddwl (io_efuse_vddwl),
  .io_pvt_test_out_ts (io_pvt_test_out_ts),
  .io_otp_vtdo (io_otp_vtdo),
  .io_otp_vrefm (io_otp_vrefm),
  .io_otp_vpp (io_otp_vpp),
  .o_lpddr_ppp_0_bp_memreset_l (o_lpddr_ppp_0_bp_memreset_l),
  .o_lpddr_ppp_1_bp_memreset_l (o_lpddr_ppp_1_bp_memreset_l),
  .o_lpddr_ppp_2_bp_memreset_l (o_lpddr_ppp_2_bp_memreset_l),
  .o_lpddr_ppp_3_bp_memreset_l (o_lpddr_ppp_3_bp_memreset_l),
  .io_lpddr_ppp_0_bp_a (io_lpddr_ppp_0_bp_a),
  .io_lpddr_ppp_1_bp_a (io_lpddr_ppp_1_bp_a),
  .io_lpddr_ppp_2_bp_a (io_lpddr_ppp_2_bp_a),
  .io_lpddr_ppp_3_bp_a (io_lpddr_ppp_3_bp_a),
  .io_lpddr_ppp_0_bp_ato (io_lpddr_ppp_0_bp_ato),
  .io_lpddr_ppp_1_bp_ato (io_lpddr_ppp_1_bp_ato),
  .io_lpddr_ppp_2_bp_ato (io_lpddr_ppp_2_bp_ato),
  .io_lpddr_ppp_3_bp_ato (io_lpddr_ppp_3_bp_ato),
  .io_lpddr_ppp_0_bp_ato_pll (io_lpddr_ppp_0_bp_ato_pll),
  .io_lpddr_ppp_1_bp_ato_pll (io_lpddr_ppp_1_bp_ato_pll),
  .io_lpddr_ppp_2_bp_ato_pll (io_lpddr_ppp_2_bp_ato_pll),
  .io_lpddr_ppp_3_bp_ato_pll (io_lpddr_ppp_3_bp_ato_pll),
  .io_lpddr_ppp_0_bp_b0_d (io_lpddr_ppp_0_bp_b0_d),
  .io_lpddr_ppp_1_bp_b0_d (io_lpddr_ppp_1_bp_b0_d),
  .io_lpddr_ppp_2_bp_b0_d (io_lpddr_ppp_2_bp_b0_d),
  .io_lpddr_ppp_3_bp_b0_d (io_lpddr_ppp_3_bp_b0_d),
  .io_lpddr_ppp_0_bp_b1_d (io_lpddr_ppp_0_bp_b1_d),
  .io_lpddr_ppp_1_bp_b1_d (io_lpddr_ppp_1_bp_b1_d),
  .io_lpddr_ppp_2_bp_b1_d (io_lpddr_ppp_2_bp_b1_d),
  .io_lpddr_ppp_3_bp_b1_d (io_lpddr_ppp_3_bp_b1_d),
  .io_lpddr_ppp_0_bp_b2_d (io_lpddr_ppp_0_bp_b2_d),
  .io_lpddr_ppp_1_bp_b2_d (io_lpddr_ppp_1_bp_b2_d),
  .io_lpddr_ppp_2_bp_b2_d (io_lpddr_ppp_2_bp_b2_d),
  .io_lpddr_ppp_3_bp_b2_d (io_lpddr_ppp_3_bp_b2_d),
  .io_lpddr_ppp_0_bp_b3_d (io_lpddr_ppp_0_bp_b3_d),
  .io_lpddr_ppp_1_bp_b3_d (io_lpddr_ppp_1_bp_b3_d),
  .io_lpddr_ppp_2_bp_b3_d (io_lpddr_ppp_2_bp_b3_d),
  .io_lpddr_ppp_3_bp_b3_d (io_lpddr_ppp_3_bp_b3_d),
  .io_lpddr_ppp_0_bp_ck0_c (io_lpddr_ppp_0_bp_ck0_c),
  .io_lpddr_ppp_1_bp_ck0_c (io_lpddr_ppp_1_bp_ck0_c),
  .io_lpddr_ppp_2_bp_ck0_c (io_lpddr_ppp_2_bp_ck0_c),
  .io_lpddr_ppp_3_bp_ck0_c (io_lpddr_ppp_3_bp_ck0_c),
  .io_lpddr_ppp_0_bp_ck0_t (io_lpddr_ppp_0_bp_ck0_t),
  .io_lpddr_ppp_1_bp_ck0_t (io_lpddr_ppp_1_bp_ck0_t),
  .io_lpddr_ppp_2_bp_ck0_t (io_lpddr_ppp_2_bp_ck0_t),
  .io_lpddr_ppp_3_bp_ck0_t (io_lpddr_ppp_3_bp_ck0_t),
  .io_lpddr_ppp_0_bp_ck1_c (io_lpddr_ppp_0_bp_ck1_c),
  .io_lpddr_ppp_1_bp_ck1_c (io_lpddr_ppp_1_bp_ck1_c),
  .io_lpddr_ppp_2_bp_ck1_c (io_lpddr_ppp_2_bp_ck1_c),
  .io_lpddr_ppp_3_bp_ck1_c (io_lpddr_ppp_3_bp_ck1_c),
  .io_lpddr_ppp_0_bp_ck1_t (io_lpddr_ppp_0_bp_ck1_t),
  .io_lpddr_ppp_1_bp_ck1_t (io_lpddr_ppp_1_bp_ck1_t),
  .io_lpddr_ppp_2_bp_ck1_t (io_lpddr_ppp_2_bp_ck1_t),
  .io_lpddr_ppp_3_bp_ck1_t (io_lpddr_ppp_3_bp_ck1_t),
  .io_lpddr_ppp_0_bp_zn (io_lpddr_ppp_0_bp_zn),
  .io_lpddr_ppp_1_bp_zn (io_lpddr_ppp_1_bp_zn),
  .io_lpddr_ppp_2_bp_zn (io_lpddr_ppp_2_bp_zn),
  .io_lpddr_ppp_3_bp_zn (io_lpddr_ppp_3_bp_zn),
  .o_lpddr_graph_0_bp_memreset_l (o_lpddr_graph_0_bp_memreset_l),
  .o_lpddr_graph_1_bp_memreset_l (o_lpddr_graph_1_bp_memreset_l),
  .o_lpddr_graph_2_bp_memreset_l (o_lpddr_graph_2_bp_memreset_l),
  .o_lpddr_graph_3_bp_memreset_l (o_lpddr_graph_3_bp_memreset_l),
  .io_lpddr_graph_0_bp_a (io_lpddr_graph_0_bp_a),
  .io_lpddr_graph_1_bp_a (io_lpddr_graph_1_bp_a),
  .io_lpddr_graph_2_bp_a (io_lpddr_graph_2_bp_a),
  .io_lpddr_graph_3_bp_a (io_lpddr_graph_3_bp_a),
  .io_lpddr_graph_0_bp_ato (io_lpddr_graph_0_bp_ato),
  .io_lpddr_graph_1_bp_ato (io_lpddr_graph_1_bp_ato),
  .io_lpddr_graph_2_bp_ato (io_lpddr_graph_2_bp_ato),
  .io_lpddr_graph_3_bp_ato (io_lpddr_graph_3_bp_ato),
  .io_lpddr_graph_0_bp_ato_pll (io_lpddr_graph_0_bp_ato_pll),
  .io_lpddr_graph_1_bp_ato_pll (io_lpddr_graph_1_bp_ato_pll),
  .io_lpddr_graph_2_bp_ato_pll (io_lpddr_graph_2_bp_ato_pll),
  .io_lpddr_graph_3_bp_ato_pll (io_lpddr_graph_3_bp_ato_pll),
  .io_lpddr_graph_0_bp_b0_d (io_lpddr_graph_0_bp_b0_d),
  .io_lpddr_graph_1_bp_b0_d (io_lpddr_graph_1_bp_b0_d),
  .io_lpddr_graph_2_bp_b0_d (io_lpddr_graph_2_bp_b0_d),
  .io_lpddr_graph_3_bp_b0_d (io_lpddr_graph_3_bp_b0_d),
  .io_lpddr_graph_0_bp_b1_d (io_lpddr_graph_0_bp_b1_d),
  .io_lpddr_graph_1_bp_b1_d (io_lpddr_graph_1_bp_b1_d),
  .io_lpddr_graph_2_bp_b1_d (io_lpddr_graph_2_bp_b1_d),
  .io_lpddr_graph_3_bp_b1_d (io_lpddr_graph_3_bp_b1_d),
  .io_lpddr_graph_0_bp_b2_d (io_lpddr_graph_0_bp_b2_d),
  .io_lpddr_graph_1_bp_b2_d (io_lpddr_graph_1_bp_b2_d),
  .io_lpddr_graph_2_bp_b2_d (io_lpddr_graph_2_bp_b2_d),
  .io_lpddr_graph_3_bp_b2_d (io_lpddr_graph_3_bp_b2_d),
  .io_lpddr_graph_0_bp_b3_d (io_lpddr_graph_0_bp_b3_d),
  .io_lpddr_graph_1_bp_b3_d (io_lpddr_graph_1_bp_b3_d),
  .io_lpddr_graph_2_bp_b3_d (io_lpddr_graph_2_bp_b3_d),
  .io_lpddr_graph_3_bp_b3_d (io_lpddr_graph_3_bp_b3_d),
  .io_lpddr_graph_0_bp_ck0_c (io_lpddr_graph_0_bp_ck0_c),
  .io_lpddr_graph_1_bp_ck0_c (io_lpddr_graph_1_bp_ck0_c),
  .io_lpddr_graph_2_bp_ck0_c (io_lpddr_graph_2_bp_ck0_c),
  .io_lpddr_graph_3_bp_ck0_c (io_lpddr_graph_3_bp_ck0_c),
  .io_lpddr_graph_0_bp_ck0_t (io_lpddr_graph_0_bp_ck0_t),
  .io_lpddr_graph_1_bp_ck0_t (io_lpddr_graph_1_bp_ck0_t),
  .io_lpddr_graph_2_bp_ck0_t (io_lpddr_graph_2_bp_ck0_t),
  .io_lpddr_graph_3_bp_ck0_t (io_lpddr_graph_3_bp_ck0_t),
  .io_lpddr_graph_0_bp_ck1_c (io_lpddr_graph_0_bp_ck1_c),
  .io_lpddr_graph_1_bp_ck1_c (io_lpddr_graph_1_bp_ck1_c),
  .io_lpddr_graph_2_bp_ck1_c (io_lpddr_graph_2_bp_ck1_c),
  .io_lpddr_graph_3_bp_ck1_c (io_lpddr_graph_3_bp_ck1_c),
  .io_lpddr_graph_0_bp_ck1_t (io_lpddr_graph_0_bp_ck1_t),
  .io_lpddr_graph_1_bp_ck1_t (io_lpddr_graph_1_bp_ck1_t),
  .io_lpddr_graph_2_bp_ck1_t (io_lpddr_graph_2_bp_ck1_t),
  .io_lpddr_graph_3_bp_ck1_t (io_lpddr_graph_3_bp_ck1_t),
  .io_lpddr_graph_0_bp_zn (io_lpddr_graph_0_bp_zn),
  .io_lpddr_graph_1_bp_zn (io_lpddr_graph_1_bp_zn),
  .io_lpddr_graph_2_bp_zn (io_lpddr_graph_2_bp_zn),
  .io_lpddr_graph_3_bp_zn (io_lpddr_graph_3_bp_zn),
  .i_pcie_perst_n (u_europa_io_to_u_aipu__o_pcie_perst_n),
  .io_pcie_resref (io_pcie_resref),
  .i_ref_pad_clk_p (i_ref_pad_clk_p),
  .i_ref_pad_clk_m (i_ref_pad_clk_m),
  .i_pcie_rxm_00 (i_pcie_rxm_00),
  .i_pcie_rxm_01 (i_pcie_rxm_01),
  .i_pcie_rxm_02 (i_pcie_rxm_02),
  .i_pcie_rxm_03 (i_pcie_rxm_03),
  .i_pcie_rxp_00 (i_pcie_rxp_00),
  .i_pcie_rxp_01 (i_pcie_rxp_01),
  .i_pcie_rxp_02 (i_pcie_rxp_02),
  .i_pcie_rxp_03 (i_pcie_rxp_03),
  .o_pcie_txm_00 (o_pcie_txm_00),
  .o_pcie_txm_01 (o_pcie_txm_01),
  .o_pcie_txm_02 (o_pcie_txm_02),
  .o_pcie_txm_03 (o_pcie_txm_03),
  .o_pcie_txp_00 (o_pcie_txp_00),
  .o_pcie_txp_01 (o_pcie_txp_01),
  .o_pcie_txp_02 (o_pcie_txp_02),
  .o_pcie_txp_03 (o_pcie_txp_03)
);
europa_io u_europa_io (
  .o_ref_clk (u_europa_io_to_u_aipu__o_ref_clk),
  .i_ref_clk_sel_freq (u_aipu_to_u_europa_io__o_ref_clk_sel_freq),
  .o_pad_ref_clk (o_ref_clk),
  .i_pad_ref_clk (i_ref_clk),
  .i_pad_ref_clk_bypass (i_ref_clk_bypass),
  .o_tck (u_europa_io_to_u_aipu__o_tck),
  .i_clk_schmitt (u_aipu_to_u_europa_io__o_clk_schmitt),
  .i_pad_tck (i_tck),
  .i_spi_clk (u_aipu_to_u_europa_io__o_spi_clk_out),
  .i_spi_drive (u_aipu_to_u_europa_io__o_spi_drive),
  .o_pad_spi_clk_out (o_spi_clk_out),
  .i_sd_emmc_clk (u_aipu_to_u_europa_io__o_mem_webar_opad),
  .i_sd_emmc_clk_oe (u_aipu_to_u_europa_io__o_mem_webar_oepad),
  .i_emmc_drive (u_aipu_to_u_europa_io__o_emmc_drive),
  .i_emmc_schmitt (u_aipu_to_u_europa_io__o_emmc_schmitt),
  .o_pad_sd_emmc_clk_out (o_sd_emmc_clk_out),
  .o_ssn_bus_0_clk (u_europa_io_to_u_aipu__o_ssn_bus_0_clk),
  .i_dft_pulldown ('0),
  .i_dft_drive (u_aipu_to_u_europa_io__o_dft_drive),
  .i_pad_ssn_bus_0_clk (i_ssn_bus_0_clk),
  .o_ssn_bus_1_clk (u_europa_io_to_u_aipu__o_ssn_bus_1_clk),
  .i_pad_ssn_bus_1_clk (i_ssn_bus_1_clk),
  .o_por_rst_n (u_europa_io_to_u_aipu__o_por_rst_n),
  .i_rst_schmitt (u_aipu_to_u_europa_io__o_rst_schmitt),
  .i_pad_por_rst_n (i_por_rst_n),
  .o_pcie_perst_n (u_europa_io_to_u_aipu__o_pcie_perst_n),
  .i_pad_pcie_perst_n (i_pcie_perst_n),
  .o_trst_n (u_europa_io_to_u_aipu__o_trst_n),
  .i_pad_trst_n (i_trst_n),
  .o_uart_rx (u_europa_io_to_u_aipu__o_uart_rx),
  .i_uart_rx_pd_en (u_aipu_to_u_europa_io__o_uart_rx_pd_en),
  .i_uart_schmitt (u_aipu_to_u_europa_io__o_uart_schmitt),
  .o_dft_uart_rx_inp (),
  .i_dft_uart_rx_inp_en ('0),
  .i_dft_uart_rx_pull_type ('0),
  .i_dft_uart_rx_pull_en ('0),
  .i_dft_uart_rx_schmitt ('0),
  .i_dft_uart_rx_drive ('0),
  .i_pad_uart_rx (i_uart_rx),
  .i_uart_tx (u_aipu_to_u_europa_io__o_uart_tx),
  .i_uart_drive (u_aipu_to_u_europa_io__o_uart_drive),
  .i_dft_uart_tx_oup ('0),
  .i_dft_uart_tx_oup_en ('0),
  .i_dft_uart_tx_pull_type ('0),
  .i_dft_uart_tx_pull_en ('0),
  .i_dft_uart_tx_schmitt ('0),
  .i_dft_uart_tx_drive ('0),
  .o_pad_uart_tx (o_uart_tx),
  .o_uart_cts_n (u_europa_io_to_u_aipu__o_uart_cts_n),
  .i_uart_cts_n_pd_en (u_aipu_to_u_europa_io__o_uart_cts_n_pd_en),
  .o_dft_uart_cts_n_inp (),
  .i_dft_uart_cts_n_inp_en ('0),
  .i_dft_uart_cts_n_pull_type ('0),
  .i_dft_uart_cts_n_pull_en ('0),
  .i_dft_uart_cts_n_schmitt ('0),
  .i_dft_uart_cts_n_drive ('0),
  .i_pad_uart_cts_n (i_uart_cts_n),
  .i_uart_rts_n (u_aipu_to_u_europa_io__o_uart_rts_n),
  .i_dft_uart_rts_n_oup ('0),
  .i_dft_uart_rts_n_oup_en ('0),
  .i_dft_uart_rts_n_pull_type ('0),
  .i_dft_uart_rts_n_pull_en ('0),
  .i_dft_uart_rts_n_schmitt ('0),
  .i_dft_uart_rts_n_drive ('0),
  .o_pad_uart_rts_n (o_uart_rts_n),
  .i_spi_ss_n (u_aipu_to_u_europa_io__o_spi_ss_n),
  .i_dft_spi_ss_n_oup ('0),
  .i_dft_spi_ss_n_oup_en ('0),
  .i_dft_spi_ss_n_pull_type ('0),
  .i_dft_spi_ss_n_pull_en ('0),
  .i_dft_spi_ss_n_schmitt ('0),
  .i_dft_spi_ss_n_drive ('0),
  .o_pad_spi_ss_n (o_spi_ss_n),
  .i_spi_sd (u_aipu_to_u_europa_io__o_spi_sd),
  .i_spi_sd_oe_n (u_aipu_to_u_europa_io__o_spi_sd_oe_n),
  .o_spi_sd (u_europa_io_to_u_aipu__o_spi_sd),
  .i_spi_sd_pd_en (u_aipu_to_u_europa_io__o_spi_sd_pd_en),
  .i_spi_schmitt (u_aipu_to_u_europa_io__o_spi_schmitt),
  .i_dft_spi_sd_oup ('0),
  .i_dft_spi_sd_oup_en ('0),
  .o_dft_spi_sd_inp (),
  .i_dft_spi_sd_inp_en ('0),
  .i_dft_spi_sd_pull_type ('0),
  .i_dft_spi_sd_pull_en ('0),
  .i_dft_spi_sd_schmitt ('0),
  .i_dft_spi_sd_drive ('0),
  .io_pad_spi_sd (io_spi_sd),
  .i_i2c_0_clk_oe (u_aipu_to_u_europa_io__o_i2c_0_clk_oe),
  .o_i2c_0_clk (u_europa_io_to_u_aipu__o_i2c_0_clk),
  .i_i2c_drive (u_aipu_to_u_europa_io__o_i2c_drive),
  .i_i2c_schmitt (u_aipu_to_u_europa_io__o_i2c_schmitt),
  .i_dft_i2c_0_clk_oup ('0),
  .i_dft_i2c_0_clk_oup_en ('0),
  .o_dft_i2c_0_clk_inp (),
  .i_dft_i2c_0_clk_inp_en ('0),
  .i_dft_i2c_0_clk_pull_type ('0),
  .i_dft_i2c_0_clk_pull_en ('0),
  .i_dft_i2c_0_clk_schmitt ('0),
  .i_dft_i2c_0_clk_drive ('0),
  .io_pad_i2c_0_clk (io_i2c_0_clk),
  .i_i2c_1_clk_oe (u_aipu_to_u_europa_io__o_i2c_1_clk_oe),
  .o_i2c_1_clk (u_europa_io_to_u_aipu__o_i2c_1_clk),
  .i_dft_i2c_1_clk_oup ('0),
  .i_dft_i2c_1_clk_oup_en ('0),
  .o_dft_i2c_1_clk_inp (),
  .i_dft_i2c_1_clk_inp_en ('0),
  .i_dft_i2c_1_clk_pull_type ('0),
  .i_dft_i2c_1_clk_pull_en ('0),
  .i_dft_i2c_1_clk_schmitt ('0),
  .i_dft_i2c_1_clk_drive ('0),
  .io_pad_i2c_1_clk (io_i2c_1_clk),
  .i_i2c_0_data_oe (u_aipu_to_u_europa_io__o_i2c_0_data_oe),
  .o_i2c_0_data (u_europa_io_to_u_aipu__o_i2c_0_data),
  .i_dft_i2c_0_data_oup ('0),
  .i_dft_i2c_0_data_oup_en ('0),
  .o_dft_i2c_0_data_inp (),
  .i_dft_i2c_0_data_inp_en ('0),
  .i_dft_i2c_0_data_pull_type ('0),
  .i_dft_i2c_0_data_pull_en ('0),
  .i_dft_i2c_0_data_schmitt ('0),
  .i_dft_i2c_0_data_drive ('0),
  .io_pad_i2c_0_data (io_i2c_0_data),
  .i_i2c_1_data_oe (u_aipu_to_u_europa_io__o_i2c_1_data_oe),
  .o_i2c_1_data (u_europa_io_to_u_aipu__o_i2c_1_data),
  .i_dft_i2c_1_data_oup ('0),
  .i_dft_i2c_1_data_oup_en ('0),
  .o_dft_i2c_1_data_inp (),
  .i_dft_i2c_1_data_inp_en ('0),
  .i_dft_i2c_1_data_pull_type ('0),
  .i_dft_i2c_1_data_pull_en ('0),
  .i_dft_i2c_1_data_schmitt ('0),
  .i_dft_i2c_1_data_drive ('0),
  .io_pad_i2c_1_data (io_i2c_1_data),
  .i_gpio (u_aipu_to_u_europa_io__o_gpio),
  .i_gpio_oe (u_aipu_to_u_europa_io__o_gpio_oe),
  .o_gpio (u_europa_io_to_u_aipu__o_gpio),
  .i_gpio_pd_en (u_aipu_to_u_europa_io__o_gpio_pd_en),
  .i_gpio_drive (u_aipu_to_u_europa_io__o_gpio_drive),
  .i_gpio_schmitt (u_aipu_to_u_europa_io__o_gpio_schmitt),
  .i_dft_gpio_oup ('0),
  .i_dft_gpio_oup_en ('0),
  .o_dft_gpio_inp (),
  .i_dft_gpio_inp_en ('0),
  .i_dft_gpio_pull_type ('0),
  .i_dft_gpio_pull_en ('0),
  .i_dft_gpio_schmitt ('0),
  .i_dft_gpio_drive ('0),
  .io_pad_gpio (io_gpio),
  .i_sd_emmc_cmd (u_aipu_to_u_europa_io__o_mem_cmd_opad),
  .i_sd_emmc_cmd_oe (u_aipu_to_u_europa_io__o_mem_cmd_oepad),
  .o_sd_emmc_cmd (u_europa_io_to_u_aipu__o_sd_emmc_cmd),
  .i_sd_emmc_cmd_ie (u_aipu_to_u_europa_io__o_mem_cmd_iepad),
  .io_pad_sd_emmc_cmd (io_sd_emmc_cmd),
  .i_sd_emmc_data (u_aipu_to_u_europa_io__o_mem_data_opad),
  .i_sd_emmc_data_oe (u_aipu_to_u_europa_io__o_mem_data_oepad),
  .o_sd_emmc_data (u_europa_io_to_u_aipu__o_sd_emmc_data),
  .i_sd_emmc_data_ie (u_aipu_to_u_europa_io__o_mem_data_iepad),
  .io_pad_sd_emmc_data (io_sd_emmc_data),
  .o_sd_emmc_strobe (u_europa_io_to_u_aipu__o_sd_emmc_strobe),
  .i_sd_emmc_strobe_ie (u_aipu_to_u_europa_io__o_mem_dqs_iepad),
  .i_pad_sd_emmc_strobe (i_sd_emmc_strobe),
  .i_emmc_reset (u_aipu_to_u_europa_io__o_mem_rstbar_opad),
  .i_emmc_reset_oe (u_aipu_to_u_europa_io__o_mem_rstbar_oepad),
  .o_pad_emmc_reset (o_emmc_reset),
  .i_emmc_power (u_aipu_to_u_europa_io__o_mem_ctrl_1_opad),
  .i_emmc_power_oe (u_aipu_to_u_europa_io__o_mem_ctrl_1_oepad),
  .o_pad_emmc_power (o_emmc_power),
  .o_sd_emmc_detect (u_europa_io_to_u_aipu__o_sd_emmc_detect),
  .i_sd_emmc_detect_ie (u_aipu_to_u_europa_io__o_mem_ctrl_0_iepad),
  .o_dft_sd_emmc_detect_inp (),
  .i_dft_sd_emmc_detect_inp_en ('0),
  .i_dft_sd_emmc_detect_pull_type ('0),
  .i_dft_sd_emmc_detect_pull_en ('0),
  .i_dft_sd_emmc_detect_schmitt ('0),
  .i_dft_sd_emmc_detect_drive ('0),
  .i_pad_sd_emmc_detect (i_sd_emmc_detect),
  .o_sd_emmc_wp (u_europa_io_to_u_aipu__o_sd_emmc_wp),
  .i_sd_emmc_wp_ie (u_aipu_to_u_europa_io__o_mem_wpbar_iepad),
  .o_dft_sd_emmc_wp_inp (),
  .i_dft_sd_emmc_wp_inp_en ('0),
  .i_dft_sd_emmc_wp_pull_type ('0),
  .i_dft_sd_emmc_wp_pull_en ('0),
  .i_dft_sd_emmc_wp_schmitt ('0),
  .i_dft_sd_emmc_wp_drive ('0),
  .i_pad_sd_emmc_wp (i_sd_emmc_wp),
  .i_sd_emmc_pu_pd (u_aipu_to_u_europa_io__o_mem_ale_opad),
  .i_sd_emmc_pu_pd_oe (u_aipu_to_u_europa_io__o_mem_ale_oepad),
  .o_pad_sd_emmc_pu_pd (o_sd_emmc_pu_pd),
  .i_emmc_rebar (u_aipu_to_u_europa_io__o_mem_rebar_opad),
  .i_emmc_rebar_oe (u_aipu_to_u_europa_io__o_mem_rebar_oepad),
  .o_emmc_rebar (u_europa_io_to_u_aipu__o_emmc_rebar),
  .i_emmc_rebar_ie (u_aipu_to_u_europa_io__o_mem_rebar_iepad),
  .io_pad_emmc_rebar (io_emmc_rebar),
  .o_emmc_lpbk_dqs (u_europa_io_to_u_aipu__o_emmc_lpbk_dqs),
  .i_emmc_lpbk_dqs_ie (u_aipu_to_u_europa_io__o_mem_lpbk_dqs_iepad),
  .i_pad_emmc_lpbk_dqs (i_emmc_lpbk_dqs),
  .i_observability (u_aipu_to_u_europa_io__o_observability),
  .i_obs_drive (u_aipu_to_u_europa_io__o_obs_drive),
  .i_dft_observability_oup ('0),
  .i_dft_observability_oup_en ('0),
  .i_dft_observability_pull_type ('0),
  .i_dft_observability_pull_en ('0),
  .i_dft_observability_schmitt ('0),
  .i_dft_observability_drive ('0),
  .o_pad_observability (o_observability),
  .i_thermal_warning_n (u_aipu_to_u_europa_io__o_thermal_warning_n),
  .o_pad_thermal_warning_n (o_thermal_warning_n),
  .i_thermal_shutdown_n (u_aipu_to_u_europa_io__o_thermal_shutdown_n),
  .o_pad_thermal_shutdown_n (o_thermal_shutdown_n),
  .o_thermal_throttle (u_europa_io_to_u_aipu__o_thermal_throttle),
  .i_pad_thermal_throttle (i_thermal_throttle),
  .o_throttle (u_europa_io_to_u_aipu__o_throttle),
  .o_dft_throttle_inp (),
  .i_dft_throttle_inp_en ('0),
  .i_dft_throttle_pull_type ('0),
  .i_dft_throttle_pull_en ('0),
  .i_dft_throttle_schmitt ('0),
  .i_dft_throttle_drive ('0),
  .i_pad_throttle (i_throttle),
  .o_boot_mode (u_europa_io_to_u_aipu__o_boot_mode),
  .i_bootmode_pull_en (u_aipu_to_u_europa_io__o_bootmode_pull_en),
  .i_pad_boot_mode (i_boot_mode),
  .o_tms (u_europa_io_to_u_aipu__o_tms),
  .i_pad_tms (i_tms),
  .o_td (u_europa_io_to_u_aipu__o_td),
  .i_pad_td_in (i_td_in),
  .i_td (u_aipu_to_u_europa_io__o_td),
  .i_jtag_drive (u_aipu_to_u_europa_io__o_jtag_drive),
  .o_pad_td_out (o_td_out),
  .i_dft_test (u_aipu_to_u_europa_io__o_dft_test),
  .i_dft_test_oe (u_aipu_to_u_europa_io__o_dft_test_oe),
  .o_dft_test (u_europa_io_to_u_aipu__o_dft_test),
  .i_dft_pull_en ('0),
  .i_dft_pull_type ('0),
  .i_dft_schmitt (u_aipu_to_u_europa_io__o_dft_schmitt),
  .io_pad_dft_test (io_dft_test),
  .i_dft_enable ('0)
);


endmodule
`endif  // EUROPA_SV
