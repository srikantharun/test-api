bind pcie_p Axi4PC # (
				.DATA_WIDTH(PCIE_LP_AXI_DATA_WIDTH),
                .ADDR_WIDTH(PCIE_LP_AXI_ADDR_WIDTH),
				.RID_WIDTH  (PCIE_LP_AXI_ID_WIDTH),
				.WID_WIDTH  (PCIE_LP_AXI_ID_WIDTH),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
        .AWREADY_MAXWAITS ( 50 ),
        .ARREADY_MAXWAITS ( 50 ),
        .WREADY_MAXWAITS ( 50 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_AIP_PCIE_lp_s_protocol_checker
				(
				.ACLK(pcie_ctrl_axi_s_clk),
				.ARESETn(pcie_ctrl_axi_s_rst_n),
				.ARVALID(pcie_ctrl_axi_s_arvalid),
				.ARADDR(pcie_ctrl_axi_s_araddr ),
				.ARLEN(pcie_ctrl_axi_s_arlen),
				.ARSIZE( pcie_ctrl_axi_s_arsize),
				.ARBURST( pcie_ctrl_axi_s_arburst ),
				.ARLOCK( pcie_ctrl_axi_s_arlock),
				.ARCACHE( pcie_ctrl_axi_s_arcache ),
				.ARPROT( pcie_ctrl_axi_s_arprot ),
				.ARID( pcie_ctrl_axi_s_arid ),
				.ARREADY( pcie_ctrl_axi_s_arready ),
				.RREADY( pcie_ctrl_axi_s_rready ),
				.RVALID( pcie_ctrl_axi_s_rvalid ),
				.RLAST( pcie_ctrl_axi_s_rlast ),
				.RDATA( pcie_ctrl_axi_s_rdata ),
				.RRESP( pcie_ctrl_axi_s_rresp ),
				.RID( pcie_ctrl_axi_s_rid ),
				.AWVALID( pcie_ctrl_axi_s_awvalid ),
				.AWADDR( pcie_ctrl_axi_s_awaddr ),
				.AWLEN( pcie_ctrl_axi_s_awlen),
				.AWSIZE( pcie_ctrl_axi_s_awsize ),
				.AWBURST( pcie_ctrl_axi_s_awburst ),
				.AWLOCK( pcie_ctrl_axi_s_awlock ),
				.AWCACHE( pcie_ctrl_axi_s_awcache ),
				.AWPROT( pcie_ctrl_axi_s_awprot ),
				.AWID( pcie_ctrl_axi_s_awid ),
				.AWREADY( pcie_ctrl_axi_s_awready ),
				.WVALID( pcie_ctrl_axi_s_wvalid ),
				.WLAST( pcie_ctrl_axi_s_wlast ),
				.WDATA( pcie_ctrl_axi_s_wdata ),
				.WSTRB( pcie_ctrl_axi_s_wstrb ),
				.WREADY( pcie_ctrl_axi_s_wready),
				.BREADY( pcie_ctrl_axi_s_bready ),
				.BVALID( pcie_ctrl_axi_s_bvalid ),
				.BRESP( pcie_ctrl_axi_s_bresp ),
				.BID( pcie_ctrl_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);





bind pcie_p Axi4PC # (
				.DATA_WIDTH(PCIE_LP_AXI_DATA_WIDTH),
                .ADDR_WIDTH(PCIE_LP_AXI_ADDR_WIDTH),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (PCIE_LP_AXI_ID_WIDTH),
				.WID_WIDTH  (PCIE_LP_AXI_ID_WIDTH),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
        .AWREADY_MAXWAITS ( 50 ),
        .ARREADY_MAXWAITS ( 50 ),
        .WREADY_MAXWAITS ( 50 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_AIP_PCIE_lp_m_protocol_checker
				(
				.ACLK(pcie_ctrl_axi_m_clk),
				.ARESETn(pcie_ctrl_axi_m_rst_n),
				.ARVALID(pcie_ctrl_axi_m_arvalid),
				.ARADDR(pcie_ctrl_axi_m_araddr ),
				.ARLEN(pcie_ctrl_axi_m_arlen),
				.ARSIZE( pcie_ctrl_axi_m_arsize),
				.ARBURST( pcie_ctrl_axi_m_arburst ),
				.ARLOCK( pcie_ctrl_axi_m_arlock),
				.ARCACHE( pcie_ctrl_axi_m_arcache ),
				.ARPROT( pcie_ctrl_axi_m_arprot ),
				.ARID( pcie_ctrl_axi_m_arid ),
				.ARREADY( pcie_ctrl_axi_m_arready ),
				.RREADY( pcie_ctrl_axi_m_rready ),
				.RVALID( pcie_ctrl_axi_m_rvalid ),
				.RLAST( pcie_ctrl_axi_m_rlast ),
				.RDATA( pcie_ctrl_axi_m_rdata ),
				.RRESP( pcie_ctrl_axi_m_rresp ),
				.RID( pcie_ctrl_axi_m_rid ),
				.AWVALID( pcie_ctrl_axi_m_awvalid ),
				.AWADDR( pcie_ctrl_axi_m_awaddr ),
				.AWLEN( pcie_ctrl_axi_m_awlen),
				.AWSIZE( pcie_ctrl_axi_m_awsize ),
				.AWBURST( pcie_ctrl_axi_m_awburst ),
				.AWLOCK( pcie_ctrl_axi_m_awlock ),
				.AWCACHE( pcie_ctrl_axi_m_awcache ),
				.AWPROT( pcie_ctrl_axi_m_awprot ),
				.AWID( pcie_ctrl_axi_m_awid ),
				.AWREADY( pcie_ctrl_axi_m_awready ),
				.WVALID( pcie_ctrl_axi_m_wvalid ),
				.WLAST( pcie_ctrl_axi_m_wlast ),
				.WDATA( pcie_ctrl_axi_m_wdata ),
				.WSTRB( pcie_ctrl_axi_m_wstrb ),
				.WREADY( pcie_ctrl_axi_m_wready),
				.BREADY( pcie_ctrl_axi_m_bready ),
				.BVALID( pcie_ctrl_axi_m_bvalid ),
				.BRESP( pcie_ctrl_axi_m_bresp ),
				.BID( pcie_ctrl_axi_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


bind pcie_p Axi4PC # (
				.DATA_WIDTH(PCIE_DBI_AXI_DATA_WIDTH),
                .ADDR_WIDTH(PCIE_DBI_AXI_ADDR_WIDTH),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (PCIE_DBI_AXI_ID_WIDTH),
				.WID_WIDTH  (PCIE_DBI_AXI_ID_WIDTH),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
        .AWREADY_MAXWAITS ( 50 ),
        .ARREADY_MAXWAITS ( 50 ),
        .WREADY_MAXWAITS ( 50 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_AIP_PCIE_lp_dbi_protocol_checker
				(
				.ACLK(pcie_ctrl_dbi_axi_s_clk),
				.ARESETn(pcie_ctrl_dbi_axi_s_rst_n),
				.ARVALID(pcie_ctrl_dbi_axi_s_arvalid),
				.ARADDR(pcie_ctrl_dbi_axi_s_araddr ),
				.ARLEN(pcie_ctrl_dbi_axi_s_arlen),
				.ARSIZE( pcie_ctrl_dbi_axi_s_arsize),
				.ARBURST( pcie_ctrl_dbi_axi_s_arburst ),
				.ARLOCK( pcie_ctrl_dbi_axi_s_arlock),
				.ARCACHE( pcie_ctrl_dbi_axi_s_arcache ),
				.ARPROT( pcie_ctrl_dbi_axi_s_arprot ),
				.ARID( pcie_ctrl_dbi_axi_s_arid ),
				.ARREADY( pcie_ctrl_dbi_axi_s_arready ),
				.RREADY( pcie_ctrl_dbi_axi_s_rready ),
				.RVALID( pcie_ctrl_dbi_axi_s_rvalid ),
				.RLAST( pcie_ctrl_dbi_axi_s_rlast ),
				.RDATA( pcie_ctrl_dbi_axi_s_rdata ),
				.RRESP( pcie_ctrl_dbi_axi_s_rresp ),
				.RID( pcie_ctrl_dbi_axi_s_rid ),
				.AWVALID( pcie_ctrl_dbi_axi_s_awvalid ),
				.AWADDR( pcie_ctrl_dbi_axi_s_awaddr ),
				.AWLEN( pcie_ctrl_dbi_axi_s_awlen),
				.AWSIZE( pcie_ctrl_dbi_axi_s_awsize ),
				.AWBURST( pcie_ctrl_dbi_axi_s_awburst ),
				.AWLOCK( pcie_ctrl_dbi_axi_s_awlock ),
				.AWCACHE( pcie_ctrl_dbi_axi_s_awcache ),
				.AWPROT( pcie_ctrl_dbi_axi_s_awprot ),
				.AWID( pcie_ctrl_dbi_axi_s_awid ),
				.AWREADY( pcie_ctrl_dbi_axi_s_awready ),
				.WVALID( pcie_ctrl_dbi_axi_s_wvalid ),
				.WLAST( pcie_ctrl_dbi_axi_s_wlast ),
				.WDATA(  pcie_ctrl_dbi_axi_s_wdata ),
				.WSTRB( pcie_ctrl_dbi_axi_s_wstrb ),
				.WREADY( pcie_ctrl_dbi_axi_s_wready),
				.BREADY( pcie_ctrl_dbi_axi_s_bready ),
				.BVALID( pcie_ctrl_dbi_axi_s_bvalid ),
				.BRESP( pcie_ctrl_dbi_axi_s_bresp ),
				.BID( pcie_ctrl_dbi_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

