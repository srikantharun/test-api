// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_h_west
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_h_west (
    output logic [182:0]  o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld,
    input  logic [182:0]  i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld,
    output logic [398:0]  o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld,
    input  logic [398:0]  i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld,
    output logic [398:0]  o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld,
    input  logic [398:0]  i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld,
    output logic [398:0]  o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld,
    input  logic [398:0]  i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld,
    output logic [398:0]  o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld,
    input  logic [398:0]  i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld,
    output logic [146:0]  o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld,
    input  logic [146:0]  i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w0_req_mainpde,
    output logic          lnk_buff_512_to_256_west_to_ddr_w0_req_mainprn,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w0_req_mainret,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w0_req_mainse,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainpde,
    output logic          lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainprn,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainret,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainse,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w1_req_mainpde,
    output logic          lnk_buff_512_to_256_west_to_ddr_w1_req_mainprn,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w1_req_mainret,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w1_req_mainse,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainpde,
    output logic          lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainprn,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainret,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainse,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w2_req_mainpde,
    output logic          lnk_buff_512_to_256_west_to_ddr_w2_req_mainprn,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w2_req_mainret,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w2_req_mainse,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainpde,
    output logic          lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainprn,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainret,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainse,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w3_req_mainpde,
    output logic          lnk_buff_512_to_256_west_to_ddr_w3_req_mainprn,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w3_req_mainret,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w3_req_mainse,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainpde,
    output logic          lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainprn,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainret,
    input  logic          lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainse,
    input  wire           i_noc_clk,
    input  wire           i_noc_rst_n,
    input  logic          scan_en
);

    noc_art_h_west u_noc_art_h_west (
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Data(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Head(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Rdy(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Tail(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Vld(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Data(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Head(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Rdy(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Tail(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Vld(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Data(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Head(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Rdy(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Tail(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Vld(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Data(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Head(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Rdy(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Tail(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Vld(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Data(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Head(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Rdy(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Tail(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Vld(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Data(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Head(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Rdy(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Tail(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Vld(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Data(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Head(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Rdy(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Tail(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Vld(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Data(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Head(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Rdy(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Tail(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Vld(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Data(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Head(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Rdy(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Tail(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Vld(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Data(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Head(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Rdy(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Tail(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Vld(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Data(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Head(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Rdy(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Tail(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_Vld(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Data(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Head(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Rdy(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Tail(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_Vld(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Data(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Head(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Rdy(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Tail(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_Vld(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Data(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Head(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Rdy(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Tail(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_Vld(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Data(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Head(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Rdy(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Tail(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_Vld(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Data(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Head(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Rdy(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Tail(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_Vld(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Data(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Head(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Rdy(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Tail(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_Vld(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Data(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Head(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Rdy(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Tail(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_Vld(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Data(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Head(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Rdy(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Tail(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail),
    .dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_Vld(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Data(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Head(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Rdy(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Tail(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail),
    .dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_Vld(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_mainpde(lnk_buff_512_to_256_west_to_ddr_w0_req_mainpde),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_mainprn(lnk_buff_512_to_256_west_to_ddr_w0_req_mainprn),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_mainret(lnk_buff_512_to_256_west_to_ddr_w0_req_mainret),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_mainse(lnk_buff_512_to_256_west_to_ddr_w0_req_mainse),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainpde(lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainpde),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainprn(lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainprn),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainret(lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainret),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainse(lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainse),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_mainpde(lnk_buff_512_to_256_west_to_ddr_w1_req_mainpde),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_mainprn(lnk_buff_512_to_256_west_to_ddr_w1_req_mainprn),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_mainret(lnk_buff_512_to_256_west_to_ddr_w1_req_mainret),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_mainse(lnk_buff_512_to_256_west_to_ddr_w1_req_mainse),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainpde(lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainpde),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainprn(lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainprn),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainret(lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainret),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainse(lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainse),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_mainpde(lnk_buff_512_to_256_west_to_ddr_w2_req_mainpde),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_mainprn(lnk_buff_512_to_256_west_to_ddr_w2_req_mainprn),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_mainret(lnk_buff_512_to_256_west_to_ddr_w2_req_mainret),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_mainse(lnk_buff_512_to_256_west_to_ddr_w2_req_mainse),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainpde(lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainpde),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainprn(lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainprn),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainret(lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainret),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainse(lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainse),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_mainpde(lnk_buff_512_to_256_west_to_ddr_w3_req_mainpde),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_mainprn(lnk_buff_512_to_256_west_to_ddr_w3_req_mainprn),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_mainret(lnk_buff_512_to_256_west_to_ddr_w3_req_mainret),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_mainse(lnk_buff_512_to_256_west_to_ddr_w3_req_mainse),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainpde(lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainpde),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainprn(lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainprn),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainret(lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainret),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainse(lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainse),
    .noc_clk(i_noc_clk),
    .noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
    );

endmodule
