// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description:
// All available sequences
// Owner: abond

`include "axe_dma_channel_seq_prologue.svh"
`include "axe_dma_channel_seq_epilogue.svh"
`include "axe_dma_channel_seq_base.svh"
