// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: Manuel Oliveira <manuel.oliveira@axelera.ai>

/// Bind SVA in ai_core
///

bind ai_core ai_core_sva u_ai_core_sva (.*);
