// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_v_center
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_v_center (
    output logic [686:0]                      o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld,
    output logic [182:0]                      o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data,
    output logic                              o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld,
    input  logic [182:0]                      i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld,
    output logic [182:0]                      o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data,
    output logic                              o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld,
    input  logic [182:0]                      i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld,
    input  logic [108:0]                      i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld,
    output logic [146:0]                      o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld,
    output logic [182:0]                      o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data,
    output logic                              o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head,
    input  logic                              i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy,
    output logic                              o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail,
    output logic                              o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld,
    input  logic [182:0]                      i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head,
    output logic                              o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld,
    input  logic [182:0]                      i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld,
    output logic [686:0]                      o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data,
    input  logic                              i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head,
    output logic                              o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy,
    input  logic                              i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail,
    input  logic                              i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld,
    output logic [182:0]                      o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data,
    output logic                              o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head,
    input  logic                              i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy,
    output logic                              o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail,
    output logic                              o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld,
    input  logic [686:0]                      i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld,
    input  logic [182:0]                      i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data,
    input  logic                              i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head,
    output logic                              o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy,
    input  logic                              i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail,
    input  logic                              i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld,
    output logic [182:0]                      o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data,
    output logic                              o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head,
    input  logic                              i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail,
    output logic                              o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld,
    input  logic [182:0]                      i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data,
    input  logic                              i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head,
    output logic                              o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy,
    input  logic                              i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail,
    input  logic                              i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld,
    output logic [182:0]                      o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data,
    output logic                              o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head,
    input  logic                              i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail,
    output logic                              o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld,
    input  logic [686:0]                      i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld,
    output logic [108:0]                      o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld,
    input  logic [146:0]                      i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld,
    output logic [686:0]                      o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld,
    input  logic [182:0]                      i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data,
    input  logic                              i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head,
    output logic                              o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy,
    input  logic                              i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail,
    input  logic                              i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld,
    output logic [182:0]                      o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data,
    output logic                              o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head,
    input  logic                              i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy,
    output logic                              o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail,
    output logic                              o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld,
    input  logic                              i_l2_addr_mode_port_b0,
    input  logic                              i_l2_addr_mode_port_b1,
    input  logic                              i_l2_intr_mode_port_b0,
    input  logic                              i_l2_intr_mode_port_b1,
    input  logic                              i_lpddr_graph_addr_mode_port_b0,
    input  logic                              i_lpddr_graph_addr_mode_port_b1,
    input  logic                              i_lpddr_graph_intr_mode_port_b0,
    input  logic                              i_lpddr_graph_intr_mode_port_b1,
    input  logic                              i_lpddr_ppp_addr_mode_port_b0,
    input  logic                              i_lpddr_ppp_addr_mode_port_b1,
    input  logic                              i_lpddr_ppp_intr_mode_port_b0,
    input  logic                              i_lpddr_ppp_intr_mode_port_b1,
    input  wire                               i_noc_clk,
    input  wire                               i_noc_rst_n,
    input  logic                              scan_en,
    input  wire                               i_sdma_0_aon_clk,
    input  wire                               i_sdma_0_aon_rst_n,
    input  wire                               i_sdma_0_clk,
    input  wire                               i_sdma_0_clken,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_ht_0_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_ht_0_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_ht_0_axi_s_arcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_0_init_ht_0_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_ht_0_axi_s_arlen,
    input  logic                              i_sdma_0_init_ht_0_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_ht_0_axi_s_arprot,
    output logic                              o_sdma_0_init_ht_0_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_ht_0_axi_s_arsize,
    input  logic                              i_sdma_0_init_ht_0_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t       o_sdma_0_init_ht_0_axi_s_rdata,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_0_init_ht_0_axi_s_rid,
    output logic                              o_sdma_0_init_ht_0_axi_s_rlast,
    input  logic                              i_sdma_0_init_ht_0_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_ht_0_axi_s_rresp,
    output logic                              o_sdma_0_init_ht_0_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_ht_0_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_ht_0_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_ht_0_axi_s_awcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_0_init_ht_0_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_ht_0_axi_s_awlen,
    input  logic                              i_sdma_0_init_ht_0_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_ht_0_axi_s_awprot,
    output logic                              o_sdma_0_init_ht_0_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_ht_0_axi_s_awsize,
    input  logic                              i_sdma_0_init_ht_0_axi_s_awvalid,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_0_init_ht_0_axi_s_bid,
    input  logic                              i_sdma_0_init_ht_0_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_ht_0_axi_s_bresp,
    output logic                              o_sdma_0_init_ht_0_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t       i_sdma_0_init_ht_0_axi_s_wdata,
    input  logic                              i_sdma_0_init_ht_0_axi_s_wlast,
    output logic                              o_sdma_0_init_ht_0_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t      i_sdma_0_init_ht_0_axi_s_wstrb,
    input  logic                              i_sdma_0_init_ht_0_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_ht_1_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_ht_1_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_ht_1_axi_s_arcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_0_init_ht_1_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_ht_1_axi_s_arlen,
    input  logic                              i_sdma_0_init_ht_1_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_ht_1_axi_s_arprot,
    output logic                              o_sdma_0_init_ht_1_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_ht_1_axi_s_arsize,
    input  logic                              i_sdma_0_init_ht_1_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t       o_sdma_0_init_ht_1_axi_s_rdata,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_0_init_ht_1_axi_s_rid,
    output logic                              o_sdma_0_init_ht_1_axi_s_rlast,
    input  logic                              i_sdma_0_init_ht_1_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_ht_1_axi_s_rresp,
    output logic                              o_sdma_0_init_ht_1_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_ht_1_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_ht_1_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_ht_1_axi_s_awcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_0_init_ht_1_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_ht_1_axi_s_awlen,
    input  logic                              i_sdma_0_init_ht_1_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_ht_1_axi_s_awprot,
    output logic                              o_sdma_0_init_ht_1_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_ht_1_axi_s_awsize,
    input  logic                              i_sdma_0_init_ht_1_axi_s_awvalid,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_0_init_ht_1_axi_s_bid,
    input  logic                              i_sdma_0_init_ht_1_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_ht_1_axi_s_bresp,
    output logic                              o_sdma_0_init_ht_1_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t       i_sdma_0_init_ht_1_axi_s_wdata,
    input  logic                              i_sdma_0_init_ht_1_axi_s_wlast,
    output logic                              o_sdma_0_init_ht_1_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t      i_sdma_0_init_ht_1_axi_s_wstrb,
    input  logic                              i_sdma_0_init_ht_1_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_lt_axi_s_arcache,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_0_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_lt_axi_s_arlen,
    input  logic                              i_sdma_0_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                 i_sdma_0_init_lt_axi_s_arqos,
    output logic                              o_sdma_0_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_lt_axi_s_arsize,
    input  logic                              i_sdma_0_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_0_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_0_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_0_init_lt_axi_s_awcache,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_0_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_0_init_lt_axi_s_awlen,
    input  logic                              i_sdma_0_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_0_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                 i_sdma_0_init_lt_axi_s_awqos,
    output logic                              o_sdma_0_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_0_init_lt_axi_s_awsize,
    input  logic                              i_sdma_0_init_lt_axi_s_awvalid,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_0_init_lt_axi_s_bid,
    input  logic                              i_sdma_0_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_lt_axi_s_bresp,
    output logic                              o_sdma_0_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t       o_sdma_0_init_lt_axi_s_rdata,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_0_init_lt_axi_s_rid,
    output logic                              o_sdma_0_init_lt_axi_s_rlast,
    input  logic                              i_sdma_0_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_0_init_lt_axi_s_rresp,
    output logic                              o_sdma_0_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t       i_sdma_0_init_lt_axi_s_wdata,
    input  logic                              i_sdma_0_init_lt_axi_s_wlast,
    output logic                              o_sdma_0_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t      i_sdma_0_init_lt_axi_s_wstrb,
    input  logic                              i_sdma_0_init_lt_axi_s_wvalid,
    output logic                              o_sdma_0_pwr_idle_val,
    output logic                              o_sdma_0_pwr_idle_ack,
    input  logic                              i_sdma_0_pwr_idle_req,
    input  wire                               i_sdma_0_rst_n,
    output chip_pkg::chip_axi_addr_t          o_sdma_0_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t               o_sdma_0_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t               o_sdma_0_targ_lt_axi_m_arcache,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_0_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                 o_sdma_0_targ_lt_axi_m_arlen,
    output logic                              o_sdma_0_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                o_sdma_0_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                 o_sdma_0_targ_lt_axi_m_arqos,
    input  logic                              i_sdma_0_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                o_sdma_0_targ_lt_axi_m_arsize,
    output logic                              o_sdma_0_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t          o_sdma_0_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t               o_sdma_0_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t               o_sdma_0_targ_lt_axi_m_awcache,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_0_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                 o_sdma_0_targ_lt_axi_m_awlen,
    output logic                              o_sdma_0_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                o_sdma_0_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                 o_sdma_0_targ_lt_axi_m_awqos,
    input  logic                              i_sdma_0_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                o_sdma_0_targ_lt_axi_m_awsize,
    output logic                              o_sdma_0_targ_lt_axi_m_awvalid,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_0_targ_lt_axi_m_bid,
    output logic                              o_sdma_0_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                i_sdma_0_targ_lt_axi_m_bresp,
    input  logic                              i_sdma_0_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t       i_sdma_0_targ_lt_axi_m_rdata,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_0_targ_lt_axi_m_rid,
    input  logic                              i_sdma_0_targ_lt_axi_m_rlast,
    output logic                              o_sdma_0_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                i_sdma_0_targ_lt_axi_m_rresp,
    input  logic                              i_sdma_0_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t       o_sdma_0_targ_lt_axi_m_wdata,
    output logic                              o_sdma_0_targ_lt_axi_m_wlast,
    input  logic                              i_sdma_0_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t      o_sdma_0_targ_lt_axi_m_wstrb,
    output logic                              o_sdma_0_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t       o_sdma_0_targ_syscfg_apb_m_paddr,
    output logic                              o_sdma_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t            o_sdma_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t   i_sdma_0_targ_syscfg_apb_m_prdata,
    input  logic                              i_sdma_0_targ_syscfg_apb_m_pready,
    output logic                              o_sdma_0_targ_syscfg_apb_m_psel,
    input  logic                              i_sdma_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t   o_sdma_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t   o_sdma_0_targ_syscfg_apb_m_pwdata,
    output logic                              o_sdma_0_targ_syscfg_apb_m_pwrite,
    input  wire                               i_sdma_1_aon_clk,
    input  wire                               i_sdma_1_aon_rst_n,
    input  wire                               i_sdma_1_clk,
    input  wire                               i_sdma_1_clken,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_ht_0_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_ht_0_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_ht_0_axi_s_arcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_1_init_ht_0_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_ht_0_axi_s_arlen,
    input  logic                              i_sdma_1_init_ht_0_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_ht_0_axi_s_arprot,
    output logic                              o_sdma_1_init_ht_0_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_ht_0_axi_s_arsize,
    input  logic                              i_sdma_1_init_ht_0_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t       o_sdma_1_init_ht_0_axi_s_rdata,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_1_init_ht_0_axi_s_rid,
    output logic                              o_sdma_1_init_ht_0_axi_s_rlast,
    input  logic                              i_sdma_1_init_ht_0_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_ht_0_axi_s_rresp,
    output logic                              o_sdma_1_init_ht_0_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_ht_0_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_ht_0_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_ht_0_axi_s_awcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_1_init_ht_0_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_ht_0_axi_s_awlen,
    input  logic                              i_sdma_1_init_ht_0_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_ht_0_axi_s_awprot,
    output logic                              o_sdma_1_init_ht_0_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_ht_0_axi_s_awsize,
    input  logic                              i_sdma_1_init_ht_0_axi_s_awvalid,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_1_init_ht_0_axi_s_bid,
    input  logic                              i_sdma_1_init_ht_0_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_ht_0_axi_s_bresp,
    output logic                              o_sdma_1_init_ht_0_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t       i_sdma_1_init_ht_0_axi_s_wdata,
    input  logic                              i_sdma_1_init_ht_0_axi_s_wlast,
    output logic                              o_sdma_1_init_ht_0_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t      i_sdma_1_init_ht_0_axi_s_wstrb,
    input  logic                              i_sdma_1_init_ht_0_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_ht_1_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_ht_1_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_ht_1_axi_s_arcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_1_init_ht_1_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_ht_1_axi_s_arlen,
    input  logic                              i_sdma_1_init_ht_1_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_ht_1_axi_s_arprot,
    output logic                              o_sdma_1_init_ht_1_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_ht_1_axi_s_arsize,
    input  logic                              i_sdma_1_init_ht_1_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t       o_sdma_1_init_ht_1_axi_s_rdata,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_1_init_ht_1_axi_s_rid,
    output logic                              o_sdma_1_init_ht_1_axi_s_rlast,
    input  logic                              i_sdma_1_init_ht_1_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_ht_1_axi_s_rresp,
    output logic                              o_sdma_1_init_ht_1_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_ht_1_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_ht_1_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_ht_1_axi_s_awcache,
    input  sdma_pkg::sdma_axi_ht_id_t         i_sdma_1_init_ht_1_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_ht_1_axi_s_awlen,
    input  logic                              i_sdma_1_init_ht_1_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_ht_1_axi_s_awprot,
    output logic                              o_sdma_1_init_ht_1_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_ht_1_axi_s_awsize,
    input  logic                              i_sdma_1_init_ht_1_axi_s_awvalid,
    output sdma_pkg::sdma_axi_ht_id_t         o_sdma_1_init_ht_1_axi_s_bid,
    input  logic                              i_sdma_1_init_ht_1_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_ht_1_axi_s_bresp,
    output logic                              o_sdma_1_init_ht_1_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t       i_sdma_1_init_ht_1_axi_s_wdata,
    input  logic                              i_sdma_1_init_ht_1_axi_s_wlast,
    output logic                              o_sdma_1_init_ht_1_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t      i_sdma_1_init_ht_1_axi_s_wstrb,
    input  logic                              i_sdma_1_init_ht_1_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_lt_axi_s_arcache,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_1_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_lt_axi_s_arlen,
    input  logic                              i_sdma_1_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                 i_sdma_1_init_lt_axi_s_arqos,
    output logic                              o_sdma_1_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_lt_axi_s_arsize,
    input  logic                              i_sdma_1_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t          i_sdma_1_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t               i_sdma_1_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t               i_sdma_1_init_lt_axi_s_awcache,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_1_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                 i_sdma_1_init_lt_axi_s_awlen,
    input  logic                              i_sdma_1_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                i_sdma_1_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                 i_sdma_1_init_lt_axi_s_awqos,
    output logic                              o_sdma_1_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                i_sdma_1_init_lt_axi_s_awsize,
    input  logic                              i_sdma_1_init_lt_axi_s_awvalid,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_1_init_lt_axi_s_bid,
    input  logic                              i_sdma_1_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_lt_axi_s_bresp,
    output logic                              o_sdma_1_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t       o_sdma_1_init_lt_axi_s_rdata,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_1_init_lt_axi_s_rid,
    output logic                              o_sdma_1_init_lt_axi_s_rlast,
    input  logic                              i_sdma_1_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                o_sdma_1_init_lt_axi_s_rresp,
    output logic                              o_sdma_1_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t       i_sdma_1_init_lt_axi_s_wdata,
    input  logic                              i_sdma_1_init_lt_axi_s_wlast,
    output logic                              o_sdma_1_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t      i_sdma_1_init_lt_axi_s_wstrb,
    input  logic                              i_sdma_1_init_lt_axi_s_wvalid,
    output logic                              o_sdma_1_pwr_idle_val,
    output logic                              o_sdma_1_pwr_idle_ack,
    input  logic                              i_sdma_1_pwr_idle_req,
    input  wire                               i_sdma_1_rst_n,
    output chip_pkg::chip_axi_addr_t          o_sdma_1_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t               o_sdma_1_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t               o_sdma_1_targ_lt_axi_m_arcache,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_1_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                 o_sdma_1_targ_lt_axi_m_arlen,
    output logic                              o_sdma_1_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                o_sdma_1_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                 o_sdma_1_targ_lt_axi_m_arqos,
    input  logic                              i_sdma_1_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                o_sdma_1_targ_lt_axi_m_arsize,
    output logic                              o_sdma_1_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t          o_sdma_1_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t               o_sdma_1_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t               o_sdma_1_targ_lt_axi_m_awcache,
    output sdma_pkg::sdma_axi_lt_id_t         o_sdma_1_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                 o_sdma_1_targ_lt_axi_m_awlen,
    output logic                              o_sdma_1_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                o_sdma_1_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                 o_sdma_1_targ_lt_axi_m_awqos,
    input  logic                              i_sdma_1_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                o_sdma_1_targ_lt_axi_m_awsize,
    output logic                              o_sdma_1_targ_lt_axi_m_awvalid,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_1_targ_lt_axi_m_bid,
    output logic                              o_sdma_1_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                i_sdma_1_targ_lt_axi_m_bresp,
    input  logic                              i_sdma_1_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t       i_sdma_1_targ_lt_axi_m_rdata,
    input  sdma_pkg::sdma_axi_lt_id_t         i_sdma_1_targ_lt_axi_m_rid,
    input  logic                              i_sdma_1_targ_lt_axi_m_rlast,
    output logic                              o_sdma_1_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                i_sdma_1_targ_lt_axi_m_rresp,
    input  logic                              i_sdma_1_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t       o_sdma_1_targ_lt_axi_m_wdata,
    output logic                              o_sdma_1_targ_lt_axi_m_wlast,
    input  logic                              i_sdma_1_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t      o_sdma_1_targ_lt_axi_m_wstrb,
    output logic                              o_sdma_1_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t       o_sdma_1_targ_syscfg_apb_m_paddr,
    output logic                              o_sdma_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t            o_sdma_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t   i_sdma_1_targ_syscfg_apb_m_prdata,
    input  logic                              i_sdma_1_targ_syscfg_apb_m_pready,
    output logic                              o_sdma_1_targ_syscfg_apb_m_psel,
    input  logic                              i_sdma_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t   o_sdma_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t   o_sdma_1_targ_syscfg_apb_m_pwdata,
    output logic                              o_sdma_1_targ_syscfg_apb_m_pwrite
);

    // Automated Address MSB fix: extra nets declaration
    logic[40:0] sdma_0_init_ht_0_axi_s_araddr_msb_fixed;
    logic[40:0] sdma_0_init_ht_0_axi_s_awaddr_msb_fixed;
    logic[40:0] sdma_0_init_ht_1_axi_s_araddr_msb_fixed;
    logic[40:0] sdma_0_init_ht_1_axi_s_awaddr_msb_fixed;
    logic[40:0] sdma_0_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] sdma_0_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] sdma_0_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] sdma_0_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] sdma_1_init_ht_0_axi_s_araddr_msb_fixed;
    logic[40:0] sdma_1_init_ht_0_axi_s_awaddr_msb_fixed;
    logic[40:0] sdma_1_init_ht_1_axi_s_araddr_msb_fixed;
    logic[40:0] sdma_1_init_ht_1_axi_s_awaddr_msb_fixed;
    logic[40:0] sdma_1_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] sdma_1_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] sdma_1_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] sdma_1_targ_lt_axi_m_awaddr_msb_fixed;

    // Automated Address MSB fix: Initiator-side assignments to extend addresses by 1 bit
    noc_common_addr_msb_setter u_addr_msb_fix_sdma_0_init_ht_0 (
        .i_axi_araddr_40b (i_sdma_0_init_ht_0_axi_s_araddr),
        .o_axi_araddr_41b (sdma_0_init_ht_0_axi_s_araddr_msb_fixed)
    );
    assign sdma_0_init_ht_0_axi_s_awaddr_msb_fixed = {1'b0, i_sdma_0_init_ht_0_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_sdma_0_init_ht_1 (
        .i_axi_araddr_40b (i_sdma_0_init_ht_1_axi_s_araddr),
        .o_axi_araddr_41b (sdma_0_init_ht_1_axi_s_araddr_msb_fixed)
    );
    assign sdma_0_init_ht_1_axi_s_awaddr_msb_fixed = {1'b0, i_sdma_0_init_ht_1_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_sdma_0_init_lt (
        .i_axi_araddr_40b (i_sdma_0_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (sdma_0_init_lt_axi_s_araddr_msb_fixed)
    );
    assign sdma_0_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_sdma_0_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_sdma_1_init_ht_0 (
        .i_axi_araddr_40b (i_sdma_1_init_ht_0_axi_s_araddr),
        .o_axi_araddr_41b (sdma_1_init_ht_0_axi_s_araddr_msb_fixed)
    );
    assign sdma_1_init_ht_0_axi_s_awaddr_msb_fixed = {1'b0, i_sdma_1_init_ht_0_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_sdma_1_init_ht_1 (
        .i_axi_araddr_40b (i_sdma_1_init_ht_1_axi_s_araddr),
        .o_axi_araddr_41b (sdma_1_init_ht_1_axi_s_araddr_msb_fixed)
    );
    assign sdma_1_init_ht_1_axi_s_awaddr_msb_fixed = {1'b0, i_sdma_1_init_ht_1_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_sdma_1_init_lt (
        .i_axi_araddr_40b (i_sdma_1_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (sdma_1_init_lt_axi_s_araddr_msb_fixed)
    );
    assign sdma_1_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_sdma_1_init_lt_axi_s_awaddr};

    // Automated Address MSB fix: Target-side assignments to drop unused MSB
    assign o_sdma_0_targ_lt_axi_m_araddr = sdma_0_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_sdma_0_targ_lt_axi_m_awaddr = sdma_0_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_sdma_1_targ_lt_axi_m_araddr = sdma_1_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_sdma_1_targ_lt_axi_m_awaddr = sdma_1_targ_lt_axi_m_awaddr_msb_fixed[39:0];


    noc_art_v_center u_noc_art_v_center (
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Data(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data),
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Head(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head),
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Data(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Head(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Data(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Head(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Data(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Head(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Data(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Head(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Rdy(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Tail(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail),
    .dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_Vld(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Data(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Head(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Rdy(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Tail(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail),
    .dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_Vld(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Data(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Head(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Data(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Head(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Data(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Head(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Data(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Head(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Data(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Head(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Data(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Head(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Data(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Head(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Data(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Head(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Data(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Head(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Data(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Head(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Data(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Head(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Data(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Head(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Data(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Head(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Rdy(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Tail(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Vld(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Data(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Head(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Rdy(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Tail(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Vld(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Data(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Head(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Data(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Head(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Data(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Head(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Data(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Head(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Data(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Head(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Data(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Head(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Data(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Head(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Data(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Head(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Data(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Head(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Data(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Head(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Data(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Head(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Rdy(i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Tail(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_Vld(o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Data(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Head(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Data(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Head(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Rdy(i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Tail(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_Vld(o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Data(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Head(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Rdy(o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Tail(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_Vld(i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Data(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Head(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Rdy(i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Tail(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail),
    .dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_Vld(o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Data(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Head(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Rdy(o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Tail(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail),
    .dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_Vld(i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Data(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Head(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Rdy(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Tail(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail),
    .dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_Vld(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Data(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Head(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Rdy(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Tail(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail),
    .dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_Vld(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Data(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Head(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Rdy(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Tail(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail),
    .dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_Vld(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Data(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Head(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Rdy(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Tail(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail),
    .dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_Vld(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Data(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Head(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Rdy(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Tail(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail),
    .dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_Vld(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Data(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Head(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Rdy(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Tail(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail),
    .dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_Vld(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Data(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Head(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Rdy(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Tail(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail),
    .dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_Vld(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Data(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Head(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Rdy(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Tail(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail),
    .dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_Vld(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Data(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Head(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Rdy(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Tail(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail),
    .dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_Vld(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Data(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Head(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Rdy(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Tail(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail),
    .dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_Vld(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Data(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Head(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Rdy(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Tail(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_Vld(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Data(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Head(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Rdy(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Tail(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_Vld(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Data(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Head(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Rdy(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Tail(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail),
    .dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_Vld(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Data(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Head(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Rdy(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Tail(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail),
    .dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_Vld(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Data(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Head(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Rdy(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Tail(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail),
    .dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_Vld(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Data(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Head(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Rdy(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Tail(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail),
    .dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_Vld(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Data(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Head(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Rdy(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Tail(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Vld(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Data(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Head(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Data(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Head(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Rdy(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Tail(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Vld(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Data(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Head(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Data(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Head(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Rdy(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Tail(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Vld(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Data(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Head(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Data(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Head(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Rdy(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Tail(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Vld(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Data(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Head(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Data(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Head(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Rdy(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Tail(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Vld(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Data(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Head(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Data(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Head(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Rdy(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Tail(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Vld(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Data(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Head(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Data(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Head(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Rdy(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Tail(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Vld(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Data(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Head(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Data(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Head(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Rdy(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Tail(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Vld(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Data(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Head(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Data(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Head(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Rdy(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Tail(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Vld(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Data(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Head(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Data(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Head(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Rdy(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Tail(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Vld(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Data(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Head(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Data(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Head(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Rdy(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Tail(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Vld(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Data(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Head(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Data(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Head(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Rdy(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Tail(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Vld(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Data(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Head(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Rdy(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Tail(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Vld(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Data(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Head(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Rdy(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Tail(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Vld(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Data(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Head(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Rdy(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Tail(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Vld(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Data(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Head(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Rdy(o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Tail(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_Vld(i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Data(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Head(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Data(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Head(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Rdy(o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Tail(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_Vld(i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Data(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Head(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Data(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Head(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Rdy(o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Tail(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_Vld(i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Data(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Head(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Data(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Head(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Rdy(o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Tail(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_Vld(i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Data(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Head(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Data(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Head(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Rdy(o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Tail(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_Vld(i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Data(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Head(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Data(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Head(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Rdy(o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Tail(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_Vld(i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Data(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Head(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Data(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Head(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Rdy(o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Tail(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_Vld(i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Data(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Head(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Data(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Head(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Rdy(o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Tail(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_Vld(i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Data(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Head(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Data(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Head(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Rdy(o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Tail(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_Vld(i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Data(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Head(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Data(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Head(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Rdy(o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Tail(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_Vld(i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Data(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Head(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Data(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Head(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Rdy(o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Tail(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail),
    .dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_Vld(i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Data(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Head(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Data(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Head(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Rdy(o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Tail(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail),
    .dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_Vld(i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Data(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Head(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Rdy(i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Tail(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail),
    .dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_Vld(o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Data(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Head(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Rdy(o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Tail(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail),
    .dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_Vld(i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Data(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Head(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Rdy(i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Tail(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail),
    .dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_Vld(o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld),
    .l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .noc_clk(i_noc_clk),
    .noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en),
    .sdma_0_aon_clk(i_sdma_0_aon_clk),
    .sdma_0_aon_rst_n(i_sdma_0_aon_rst_n),
    .sdma_0_clk(i_sdma_0_clk),
    .sdma_0_clken(i_sdma_0_clken),
    .sdma_0_init_ht_0_rd_Ar_Addr(sdma_0_init_ht_0_axi_s_araddr_msb_fixed),
    .sdma_0_init_ht_0_rd_Ar_Burst(i_sdma_0_init_ht_0_axi_s_arburst),
    .sdma_0_init_ht_0_rd_Ar_Cache(i_sdma_0_init_ht_0_axi_s_arcache),
    .sdma_0_init_ht_0_rd_Ar_Id(i_sdma_0_init_ht_0_axi_s_arid),
    .sdma_0_init_ht_0_rd_Ar_Len(i_sdma_0_init_ht_0_axi_s_arlen),
    .sdma_0_init_ht_0_rd_Ar_Lock(i_sdma_0_init_ht_0_axi_s_arlock),
    .sdma_0_init_ht_0_rd_Ar_Prot(i_sdma_0_init_ht_0_axi_s_arprot),
    .sdma_0_init_ht_0_rd_Ar_Ready(o_sdma_0_init_ht_0_axi_s_arready),
    .sdma_0_init_ht_0_rd_Ar_Size(i_sdma_0_init_ht_0_axi_s_arsize),
    .sdma_0_init_ht_0_rd_Ar_Valid(i_sdma_0_init_ht_0_axi_s_arvalid),
    .sdma_0_init_ht_0_rd_R_Data(o_sdma_0_init_ht_0_axi_s_rdata),
    .sdma_0_init_ht_0_rd_R_Id(o_sdma_0_init_ht_0_axi_s_rid),
    .sdma_0_init_ht_0_rd_R_Last(o_sdma_0_init_ht_0_axi_s_rlast),
    .sdma_0_init_ht_0_rd_R_Ready(i_sdma_0_init_ht_0_axi_s_rready),
    .sdma_0_init_ht_0_rd_R_Resp(o_sdma_0_init_ht_0_axi_s_rresp),
    .sdma_0_init_ht_0_rd_R_Valid(o_sdma_0_init_ht_0_axi_s_rvalid),
    .sdma_0_init_ht_0_wr_Aw_Addr(sdma_0_init_ht_0_axi_s_awaddr_msb_fixed),
    .sdma_0_init_ht_0_wr_Aw_Burst(i_sdma_0_init_ht_0_axi_s_awburst),
    .sdma_0_init_ht_0_wr_Aw_Cache(i_sdma_0_init_ht_0_axi_s_awcache),
    .sdma_0_init_ht_0_wr_Aw_Id(i_sdma_0_init_ht_0_axi_s_awid),
    .sdma_0_init_ht_0_wr_Aw_Len(i_sdma_0_init_ht_0_axi_s_awlen),
    .sdma_0_init_ht_0_wr_Aw_Lock(i_sdma_0_init_ht_0_axi_s_awlock),
    .sdma_0_init_ht_0_wr_Aw_Prot(i_sdma_0_init_ht_0_axi_s_awprot),
    .sdma_0_init_ht_0_wr_Aw_Ready(o_sdma_0_init_ht_0_axi_s_awready),
    .sdma_0_init_ht_0_wr_Aw_Size(i_sdma_0_init_ht_0_axi_s_awsize),
    .sdma_0_init_ht_0_wr_Aw_Valid(i_sdma_0_init_ht_0_axi_s_awvalid),
    .sdma_0_init_ht_0_wr_B_Id(o_sdma_0_init_ht_0_axi_s_bid),
    .sdma_0_init_ht_0_wr_B_Ready(i_sdma_0_init_ht_0_axi_s_bready),
    .sdma_0_init_ht_0_wr_B_Resp(o_sdma_0_init_ht_0_axi_s_bresp),
    .sdma_0_init_ht_0_wr_B_Valid(o_sdma_0_init_ht_0_axi_s_bvalid),
    .sdma_0_init_ht_0_wr_W_Data(i_sdma_0_init_ht_0_axi_s_wdata),
    .sdma_0_init_ht_0_wr_W_Last(i_sdma_0_init_ht_0_axi_s_wlast),
    .sdma_0_init_ht_0_wr_W_Ready(o_sdma_0_init_ht_0_axi_s_wready),
    .sdma_0_init_ht_0_wr_W_Strb(i_sdma_0_init_ht_0_axi_s_wstrb),
    .sdma_0_init_ht_0_wr_W_Valid(i_sdma_0_init_ht_0_axi_s_wvalid),
    .sdma_0_init_ht_1_rd_Ar_Addr(sdma_0_init_ht_1_axi_s_araddr_msb_fixed),
    .sdma_0_init_ht_1_rd_Ar_Burst(i_sdma_0_init_ht_1_axi_s_arburst),
    .sdma_0_init_ht_1_rd_Ar_Cache(i_sdma_0_init_ht_1_axi_s_arcache),
    .sdma_0_init_ht_1_rd_Ar_Id(i_sdma_0_init_ht_1_axi_s_arid),
    .sdma_0_init_ht_1_rd_Ar_Len(i_sdma_0_init_ht_1_axi_s_arlen),
    .sdma_0_init_ht_1_rd_Ar_Lock(i_sdma_0_init_ht_1_axi_s_arlock),
    .sdma_0_init_ht_1_rd_Ar_Prot(i_sdma_0_init_ht_1_axi_s_arprot),
    .sdma_0_init_ht_1_rd_Ar_Ready(o_sdma_0_init_ht_1_axi_s_arready),
    .sdma_0_init_ht_1_rd_Ar_Size(i_sdma_0_init_ht_1_axi_s_arsize),
    .sdma_0_init_ht_1_rd_Ar_Valid(i_sdma_0_init_ht_1_axi_s_arvalid),
    .sdma_0_init_ht_1_rd_R_Data(o_sdma_0_init_ht_1_axi_s_rdata),
    .sdma_0_init_ht_1_rd_R_Id(o_sdma_0_init_ht_1_axi_s_rid),
    .sdma_0_init_ht_1_rd_R_Last(o_sdma_0_init_ht_1_axi_s_rlast),
    .sdma_0_init_ht_1_rd_R_Ready(i_sdma_0_init_ht_1_axi_s_rready),
    .sdma_0_init_ht_1_rd_R_Resp(o_sdma_0_init_ht_1_axi_s_rresp),
    .sdma_0_init_ht_1_rd_R_Valid(o_sdma_0_init_ht_1_axi_s_rvalid),
    .sdma_0_init_ht_1_wr_Aw_Addr(sdma_0_init_ht_1_axi_s_awaddr_msb_fixed),
    .sdma_0_init_ht_1_wr_Aw_Burst(i_sdma_0_init_ht_1_axi_s_awburst),
    .sdma_0_init_ht_1_wr_Aw_Cache(i_sdma_0_init_ht_1_axi_s_awcache),
    .sdma_0_init_ht_1_wr_Aw_Id(i_sdma_0_init_ht_1_axi_s_awid),
    .sdma_0_init_ht_1_wr_Aw_Len(i_sdma_0_init_ht_1_axi_s_awlen),
    .sdma_0_init_ht_1_wr_Aw_Lock(i_sdma_0_init_ht_1_axi_s_awlock),
    .sdma_0_init_ht_1_wr_Aw_Prot(i_sdma_0_init_ht_1_axi_s_awprot),
    .sdma_0_init_ht_1_wr_Aw_Ready(o_sdma_0_init_ht_1_axi_s_awready),
    .sdma_0_init_ht_1_wr_Aw_Size(i_sdma_0_init_ht_1_axi_s_awsize),
    .sdma_0_init_ht_1_wr_Aw_Valid(i_sdma_0_init_ht_1_axi_s_awvalid),
    .sdma_0_init_ht_1_wr_B_Id(o_sdma_0_init_ht_1_axi_s_bid),
    .sdma_0_init_ht_1_wr_B_Ready(i_sdma_0_init_ht_1_axi_s_bready),
    .sdma_0_init_ht_1_wr_B_Resp(o_sdma_0_init_ht_1_axi_s_bresp),
    .sdma_0_init_ht_1_wr_B_Valid(o_sdma_0_init_ht_1_axi_s_bvalid),
    .sdma_0_init_ht_1_wr_W_Data(i_sdma_0_init_ht_1_axi_s_wdata),
    .sdma_0_init_ht_1_wr_W_Last(i_sdma_0_init_ht_1_axi_s_wlast),
    .sdma_0_init_ht_1_wr_W_Ready(o_sdma_0_init_ht_1_axi_s_wready),
    .sdma_0_init_ht_1_wr_W_Strb(i_sdma_0_init_ht_1_axi_s_wstrb),
    .sdma_0_init_ht_1_wr_W_Valid(i_sdma_0_init_ht_1_axi_s_wvalid),
    .sdma_0_init_lt_Ar_Addr(sdma_0_init_lt_axi_s_araddr_msb_fixed),
    .sdma_0_init_lt_Ar_Burst(i_sdma_0_init_lt_axi_s_arburst),
    .sdma_0_init_lt_Ar_Cache(i_sdma_0_init_lt_axi_s_arcache),
    .sdma_0_init_lt_Ar_Id(i_sdma_0_init_lt_axi_s_arid),
    .sdma_0_init_lt_Ar_Len(i_sdma_0_init_lt_axi_s_arlen),
    .sdma_0_init_lt_Ar_Lock(i_sdma_0_init_lt_axi_s_arlock),
    .sdma_0_init_lt_Ar_Prot(i_sdma_0_init_lt_axi_s_arprot),
    .sdma_0_init_lt_Ar_Qos(i_sdma_0_init_lt_axi_s_arqos),
    .sdma_0_init_lt_Ar_Ready(o_sdma_0_init_lt_axi_s_arready),
    .sdma_0_init_lt_Ar_Size(i_sdma_0_init_lt_axi_s_arsize),
    .sdma_0_init_lt_Ar_Valid(i_sdma_0_init_lt_axi_s_arvalid),
    .sdma_0_init_lt_Aw_Addr(sdma_0_init_lt_axi_s_awaddr_msb_fixed),
    .sdma_0_init_lt_Aw_Burst(i_sdma_0_init_lt_axi_s_awburst),
    .sdma_0_init_lt_Aw_Cache(i_sdma_0_init_lt_axi_s_awcache),
    .sdma_0_init_lt_Aw_Id(i_sdma_0_init_lt_axi_s_awid),
    .sdma_0_init_lt_Aw_Len(i_sdma_0_init_lt_axi_s_awlen),
    .sdma_0_init_lt_Aw_Lock(i_sdma_0_init_lt_axi_s_awlock),
    .sdma_0_init_lt_Aw_Prot(i_sdma_0_init_lt_axi_s_awprot),
    .sdma_0_init_lt_Aw_Qos(i_sdma_0_init_lt_axi_s_awqos),
    .sdma_0_init_lt_Aw_Ready(o_sdma_0_init_lt_axi_s_awready),
    .sdma_0_init_lt_Aw_Size(i_sdma_0_init_lt_axi_s_awsize),
    .sdma_0_init_lt_Aw_Valid(i_sdma_0_init_lt_axi_s_awvalid),
    .sdma_0_init_lt_B_Id(o_sdma_0_init_lt_axi_s_bid),
    .sdma_0_init_lt_B_Ready(i_sdma_0_init_lt_axi_s_bready),
    .sdma_0_init_lt_B_Resp(o_sdma_0_init_lt_axi_s_bresp),
    .sdma_0_init_lt_B_Valid(o_sdma_0_init_lt_axi_s_bvalid),
    .sdma_0_init_lt_R_Data(o_sdma_0_init_lt_axi_s_rdata),
    .sdma_0_init_lt_R_Id(o_sdma_0_init_lt_axi_s_rid),
    .sdma_0_init_lt_R_Last(o_sdma_0_init_lt_axi_s_rlast),
    .sdma_0_init_lt_R_Ready(i_sdma_0_init_lt_axi_s_rready),
    .sdma_0_init_lt_R_Resp(o_sdma_0_init_lt_axi_s_rresp),
    .sdma_0_init_lt_R_Valid(o_sdma_0_init_lt_axi_s_rvalid),
    .sdma_0_init_lt_W_Data(i_sdma_0_init_lt_axi_s_wdata),
    .sdma_0_init_lt_W_Last(i_sdma_0_init_lt_axi_s_wlast),
    .sdma_0_init_lt_W_Ready(o_sdma_0_init_lt_axi_s_wready),
    .sdma_0_init_lt_W_Strb(i_sdma_0_init_lt_axi_s_wstrb),
    .sdma_0_init_lt_W_Valid(i_sdma_0_init_lt_axi_s_wvalid),
    .sdma_0_pwr_Idle(o_sdma_0_pwr_idle_val),
    .sdma_0_pwr_IdleAck(o_sdma_0_pwr_idle_ack),
    .sdma_0_pwr_IdleReq(i_sdma_0_pwr_idle_req),
    .sdma_0_rst_n(i_sdma_0_rst_n),
    .sdma_0_targ_lt_Ar_Addr(sdma_0_targ_lt_axi_m_araddr_msb_fixed),
    .sdma_0_targ_lt_Ar_Burst(o_sdma_0_targ_lt_axi_m_arburst),
    .sdma_0_targ_lt_Ar_Cache(o_sdma_0_targ_lt_axi_m_arcache),
    .sdma_0_targ_lt_Ar_Id(o_sdma_0_targ_lt_axi_m_arid),
    .sdma_0_targ_lt_Ar_Len(o_sdma_0_targ_lt_axi_m_arlen),
    .sdma_0_targ_lt_Ar_Lock(o_sdma_0_targ_lt_axi_m_arlock),
    .sdma_0_targ_lt_Ar_Prot(o_sdma_0_targ_lt_axi_m_arprot),
    .sdma_0_targ_lt_Ar_Qos(o_sdma_0_targ_lt_axi_m_arqos),
    .sdma_0_targ_lt_Ar_Ready(i_sdma_0_targ_lt_axi_m_arready),
    .sdma_0_targ_lt_Ar_Size(o_sdma_0_targ_lt_axi_m_arsize),
    .sdma_0_targ_lt_Ar_Valid(o_sdma_0_targ_lt_axi_m_arvalid),
    .sdma_0_targ_lt_Aw_Addr(sdma_0_targ_lt_axi_m_awaddr_msb_fixed),
    .sdma_0_targ_lt_Aw_Burst(o_sdma_0_targ_lt_axi_m_awburst),
    .sdma_0_targ_lt_Aw_Cache(o_sdma_0_targ_lt_axi_m_awcache),
    .sdma_0_targ_lt_Aw_Id(o_sdma_0_targ_lt_axi_m_awid),
    .sdma_0_targ_lt_Aw_Len(o_sdma_0_targ_lt_axi_m_awlen),
    .sdma_0_targ_lt_Aw_Lock(o_sdma_0_targ_lt_axi_m_awlock),
    .sdma_0_targ_lt_Aw_Prot(o_sdma_0_targ_lt_axi_m_awprot),
    .sdma_0_targ_lt_Aw_Qos(o_sdma_0_targ_lt_axi_m_awqos),
    .sdma_0_targ_lt_Aw_Ready(i_sdma_0_targ_lt_axi_m_awready),
    .sdma_0_targ_lt_Aw_Size(o_sdma_0_targ_lt_axi_m_awsize),
    .sdma_0_targ_lt_Aw_Valid(o_sdma_0_targ_lt_axi_m_awvalid),
    .sdma_0_targ_lt_B_Id(i_sdma_0_targ_lt_axi_m_bid),
    .sdma_0_targ_lt_B_Ready(o_sdma_0_targ_lt_axi_m_bready),
    .sdma_0_targ_lt_B_Resp(i_sdma_0_targ_lt_axi_m_bresp),
    .sdma_0_targ_lt_B_Valid(i_sdma_0_targ_lt_axi_m_bvalid),
    .sdma_0_targ_lt_R_Data(i_sdma_0_targ_lt_axi_m_rdata),
    .sdma_0_targ_lt_R_Id(i_sdma_0_targ_lt_axi_m_rid),
    .sdma_0_targ_lt_R_Last(i_sdma_0_targ_lt_axi_m_rlast),
    .sdma_0_targ_lt_R_Ready(o_sdma_0_targ_lt_axi_m_rready),
    .sdma_0_targ_lt_R_Resp(i_sdma_0_targ_lt_axi_m_rresp),
    .sdma_0_targ_lt_R_Valid(i_sdma_0_targ_lt_axi_m_rvalid),
    .sdma_0_targ_lt_W_Data(o_sdma_0_targ_lt_axi_m_wdata),
    .sdma_0_targ_lt_W_Last(o_sdma_0_targ_lt_axi_m_wlast),
    .sdma_0_targ_lt_W_Ready(i_sdma_0_targ_lt_axi_m_wready),
    .sdma_0_targ_lt_W_Strb(o_sdma_0_targ_lt_axi_m_wstrb),
    .sdma_0_targ_lt_W_Valid(o_sdma_0_targ_lt_axi_m_wvalid),
    .sdma_0_targ_syscfg_PAddr(o_sdma_0_targ_syscfg_apb_m_paddr),
    .sdma_0_targ_syscfg_PEnable(o_sdma_0_targ_syscfg_apb_m_penable),
    .sdma_0_targ_syscfg_PProt(o_sdma_0_targ_syscfg_apb_m_pprot),
    .sdma_0_targ_syscfg_PRData(i_sdma_0_targ_syscfg_apb_m_prdata),
    .sdma_0_targ_syscfg_PReady(i_sdma_0_targ_syscfg_apb_m_pready),
    .sdma_0_targ_syscfg_PSel(o_sdma_0_targ_syscfg_apb_m_psel),
    .sdma_0_targ_syscfg_PSlvErr(i_sdma_0_targ_syscfg_apb_m_pslverr),
    .sdma_0_targ_syscfg_PStrb(o_sdma_0_targ_syscfg_apb_m_pstrb),
    .sdma_0_targ_syscfg_PWData(o_sdma_0_targ_syscfg_apb_m_pwdata),
    .sdma_0_targ_syscfg_PWrite(o_sdma_0_targ_syscfg_apb_m_pwrite),
    .sdma_1_aon_clk(i_sdma_1_aon_clk),
    .sdma_1_aon_rst_n(i_sdma_1_aon_rst_n),
    .sdma_1_clk(i_sdma_1_clk),
    .sdma_1_clken(i_sdma_1_clken),
    .sdma_1_init_ht_0_rd_Ar_Addr(sdma_1_init_ht_0_axi_s_araddr_msb_fixed),
    .sdma_1_init_ht_0_rd_Ar_Burst(i_sdma_1_init_ht_0_axi_s_arburst),
    .sdma_1_init_ht_0_rd_Ar_Cache(i_sdma_1_init_ht_0_axi_s_arcache),
    .sdma_1_init_ht_0_rd_Ar_Id(i_sdma_1_init_ht_0_axi_s_arid),
    .sdma_1_init_ht_0_rd_Ar_Len(i_sdma_1_init_ht_0_axi_s_arlen),
    .sdma_1_init_ht_0_rd_Ar_Lock(i_sdma_1_init_ht_0_axi_s_arlock),
    .sdma_1_init_ht_0_rd_Ar_Prot(i_sdma_1_init_ht_0_axi_s_arprot),
    .sdma_1_init_ht_0_rd_Ar_Ready(o_sdma_1_init_ht_0_axi_s_arready),
    .sdma_1_init_ht_0_rd_Ar_Size(i_sdma_1_init_ht_0_axi_s_arsize),
    .sdma_1_init_ht_0_rd_Ar_Valid(i_sdma_1_init_ht_0_axi_s_arvalid),
    .sdma_1_init_ht_0_rd_R_Data(o_sdma_1_init_ht_0_axi_s_rdata),
    .sdma_1_init_ht_0_rd_R_Id(o_sdma_1_init_ht_0_axi_s_rid),
    .sdma_1_init_ht_0_rd_R_Last(o_sdma_1_init_ht_0_axi_s_rlast),
    .sdma_1_init_ht_0_rd_R_Ready(i_sdma_1_init_ht_0_axi_s_rready),
    .sdma_1_init_ht_0_rd_R_Resp(o_sdma_1_init_ht_0_axi_s_rresp),
    .sdma_1_init_ht_0_rd_R_Valid(o_sdma_1_init_ht_0_axi_s_rvalid),
    .sdma_1_init_ht_0_wr_Aw_Addr(sdma_1_init_ht_0_axi_s_awaddr_msb_fixed),
    .sdma_1_init_ht_0_wr_Aw_Burst(i_sdma_1_init_ht_0_axi_s_awburst),
    .sdma_1_init_ht_0_wr_Aw_Cache(i_sdma_1_init_ht_0_axi_s_awcache),
    .sdma_1_init_ht_0_wr_Aw_Id(i_sdma_1_init_ht_0_axi_s_awid),
    .sdma_1_init_ht_0_wr_Aw_Len(i_sdma_1_init_ht_0_axi_s_awlen),
    .sdma_1_init_ht_0_wr_Aw_Lock(i_sdma_1_init_ht_0_axi_s_awlock),
    .sdma_1_init_ht_0_wr_Aw_Prot(i_sdma_1_init_ht_0_axi_s_awprot),
    .sdma_1_init_ht_0_wr_Aw_Ready(o_sdma_1_init_ht_0_axi_s_awready),
    .sdma_1_init_ht_0_wr_Aw_Size(i_sdma_1_init_ht_0_axi_s_awsize),
    .sdma_1_init_ht_0_wr_Aw_Valid(i_sdma_1_init_ht_0_axi_s_awvalid),
    .sdma_1_init_ht_0_wr_B_Id(o_sdma_1_init_ht_0_axi_s_bid),
    .sdma_1_init_ht_0_wr_B_Ready(i_sdma_1_init_ht_0_axi_s_bready),
    .sdma_1_init_ht_0_wr_B_Resp(o_sdma_1_init_ht_0_axi_s_bresp),
    .sdma_1_init_ht_0_wr_B_Valid(o_sdma_1_init_ht_0_axi_s_bvalid),
    .sdma_1_init_ht_0_wr_W_Data(i_sdma_1_init_ht_0_axi_s_wdata),
    .sdma_1_init_ht_0_wr_W_Last(i_sdma_1_init_ht_0_axi_s_wlast),
    .sdma_1_init_ht_0_wr_W_Ready(o_sdma_1_init_ht_0_axi_s_wready),
    .sdma_1_init_ht_0_wr_W_Strb(i_sdma_1_init_ht_0_axi_s_wstrb),
    .sdma_1_init_ht_0_wr_W_Valid(i_sdma_1_init_ht_0_axi_s_wvalid),
    .sdma_1_init_ht_1_rd_Ar_Addr(sdma_1_init_ht_1_axi_s_araddr_msb_fixed),
    .sdma_1_init_ht_1_rd_Ar_Burst(i_sdma_1_init_ht_1_axi_s_arburst),
    .sdma_1_init_ht_1_rd_Ar_Cache(i_sdma_1_init_ht_1_axi_s_arcache),
    .sdma_1_init_ht_1_rd_Ar_Id(i_sdma_1_init_ht_1_axi_s_arid),
    .sdma_1_init_ht_1_rd_Ar_Len(i_sdma_1_init_ht_1_axi_s_arlen),
    .sdma_1_init_ht_1_rd_Ar_Lock(i_sdma_1_init_ht_1_axi_s_arlock),
    .sdma_1_init_ht_1_rd_Ar_Prot(i_sdma_1_init_ht_1_axi_s_arprot),
    .sdma_1_init_ht_1_rd_Ar_Ready(o_sdma_1_init_ht_1_axi_s_arready),
    .sdma_1_init_ht_1_rd_Ar_Size(i_sdma_1_init_ht_1_axi_s_arsize),
    .sdma_1_init_ht_1_rd_Ar_Valid(i_sdma_1_init_ht_1_axi_s_arvalid),
    .sdma_1_init_ht_1_rd_R_Data(o_sdma_1_init_ht_1_axi_s_rdata),
    .sdma_1_init_ht_1_rd_R_Id(o_sdma_1_init_ht_1_axi_s_rid),
    .sdma_1_init_ht_1_rd_R_Last(o_sdma_1_init_ht_1_axi_s_rlast),
    .sdma_1_init_ht_1_rd_R_Ready(i_sdma_1_init_ht_1_axi_s_rready),
    .sdma_1_init_ht_1_rd_R_Resp(o_sdma_1_init_ht_1_axi_s_rresp),
    .sdma_1_init_ht_1_rd_R_Valid(o_sdma_1_init_ht_1_axi_s_rvalid),
    .sdma_1_init_ht_1_wr_Aw_Addr(sdma_1_init_ht_1_axi_s_awaddr_msb_fixed),
    .sdma_1_init_ht_1_wr_Aw_Burst(i_sdma_1_init_ht_1_axi_s_awburst),
    .sdma_1_init_ht_1_wr_Aw_Cache(i_sdma_1_init_ht_1_axi_s_awcache),
    .sdma_1_init_ht_1_wr_Aw_Id(i_sdma_1_init_ht_1_axi_s_awid),
    .sdma_1_init_ht_1_wr_Aw_Len(i_sdma_1_init_ht_1_axi_s_awlen),
    .sdma_1_init_ht_1_wr_Aw_Lock(i_sdma_1_init_ht_1_axi_s_awlock),
    .sdma_1_init_ht_1_wr_Aw_Prot(i_sdma_1_init_ht_1_axi_s_awprot),
    .sdma_1_init_ht_1_wr_Aw_Ready(o_sdma_1_init_ht_1_axi_s_awready),
    .sdma_1_init_ht_1_wr_Aw_Size(i_sdma_1_init_ht_1_axi_s_awsize),
    .sdma_1_init_ht_1_wr_Aw_Valid(i_sdma_1_init_ht_1_axi_s_awvalid),
    .sdma_1_init_ht_1_wr_B_Id(o_sdma_1_init_ht_1_axi_s_bid),
    .sdma_1_init_ht_1_wr_B_Ready(i_sdma_1_init_ht_1_axi_s_bready),
    .sdma_1_init_ht_1_wr_B_Resp(o_sdma_1_init_ht_1_axi_s_bresp),
    .sdma_1_init_ht_1_wr_B_Valid(o_sdma_1_init_ht_1_axi_s_bvalid),
    .sdma_1_init_ht_1_wr_W_Data(i_sdma_1_init_ht_1_axi_s_wdata),
    .sdma_1_init_ht_1_wr_W_Last(i_sdma_1_init_ht_1_axi_s_wlast),
    .sdma_1_init_ht_1_wr_W_Ready(o_sdma_1_init_ht_1_axi_s_wready),
    .sdma_1_init_ht_1_wr_W_Strb(i_sdma_1_init_ht_1_axi_s_wstrb),
    .sdma_1_init_ht_1_wr_W_Valid(i_sdma_1_init_ht_1_axi_s_wvalid),
    .sdma_1_init_lt_Ar_Addr(sdma_1_init_lt_axi_s_araddr_msb_fixed),
    .sdma_1_init_lt_Ar_Burst(i_sdma_1_init_lt_axi_s_arburst),
    .sdma_1_init_lt_Ar_Cache(i_sdma_1_init_lt_axi_s_arcache),
    .sdma_1_init_lt_Ar_Id(i_sdma_1_init_lt_axi_s_arid),
    .sdma_1_init_lt_Ar_Len(i_sdma_1_init_lt_axi_s_arlen),
    .sdma_1_init_lt_Ar_Lock(i_sdma_1_init_lt_axi_s_arlock),
    .sdma_1_init_lt_Ar_Prot(i_sdma_1_init_lt_axi_s_arprot),
    .sdma_1_init_lt_Ar_Qos(i_sdma_1_init_lt_axi_s_arqos),
    .sdma_1_init_lt_Ar_Ready(o_sdma_1_init_lt_axi_s_arready),
    .sdma_1_init_lt_Ar_Size(i_sdma_1_init_lt_axi_s_arsize),
    .sdma_1_init_lt_Ar_Valid(i_sdma_1_init_lt_axi_s_arvalid),
    .sdma_1_init_lt_Aw_Addr(sdma_1_init_lt_axi_s_awaddr_msb_fixed),
    .sdma_1_init_lt_Aw_Burst(i_sdma_1_init_lt_axi_s_awburst),
    .sdma_1_init_lt_Aw_Cache(i_sdma_1_init_lt_axi_s_awcache),
    .sdma_1_init_lt_Aw_Id(i_sdma_1_init_lt_axi_s_awid),
    .sdma_1_init_lt_Aw_Len(i_sdma_1_init_lt_axi_s_awlen),
    .sdma_1_init_lt_Aw_Lock(i_sdma_1_init_lt_axi_s_awlock),
    .sdma_1_init_lt_Aw_Prot(i_sdma_1_init_lt_axi_s_awprot),
    .sdma_1_init_lt_Aw_Qos(i_sdma_1_init_lt_axi_s_awqos),
    .sdma_1_init_lt_Aw_Ready(o_sdma_1_init_lt_axi_s_awready),
    .sdma_1_init_lt_Aw_Size(i_sdma_1_init_lt_axi_s_awsize),
    .sdma_1_init_lt_Aw_Valid(i_sdma_1_init_lt_axi_s_awvalid),
    .sdma_1_init_lt_B_Id(o_sdma_1_init_lt_axi_s_bid),
    .sdma_1_init_lt_B_Ready(i_sdma_1_init_lt_axi_s_bready),
    .sdma_1_init_lt_B_Resp(o_sdma_1_init_lt_axi_s_bresp),
    .sdma_1_init_lt_B_Valid(o_sdma_1_init_lt_axi_s_bvalid),
    .sdma_1_init_lt_R_Data(o_sdma_1_init_lt_axi_s_rdata),
    .sdma_1_init_lt_R_Id(o_sdma_1_init_lt_axi_s_rid),
    .sdma_1_init_lt_R_Last(o_sdma_1_init_lt_axi_s_rlast),
    .sdma_1_init_lt_R_Ready(i_sdma_1_init_lt_axi_s_rready),
    .sdma_1_init_lt_R_Resp(o_sdma_1_init_lt_axi_s_rresp),
    .sdma_1_init_lt_R_Valid(o_sdma_1_init_lt_axi_s_rvalid),
    .sdma_1_init_lt_W_Data(i_sdma_1_init_lt_axi_s_wdata),
    .sdma_1_init_lt_W_Last(i_sdma_1_init_lt_axi_s_wlast),
    .sdma_1_init_lt_W_Ready(o_sdma_1_init_lt_axi_s_wready),
    .sdma_1_init_lt_W_Strb(i_sdma_1_init_lt_axi_s_wstrb),
    .sdma_1_init_lt_W_Valid(i_sdma_1_init_lt_axi_s_wvalid),
    .sdma_1_pwr_Idle(o_sdma_1_pwr_idle_val),
    .sdma_1_pwr_IdleAck(o_sdma_1_pwr_idle_ack),
    .sdma_1_pwr_IdleReq(i_sdma_1_pwr_idle_req),
    .sdma_1_rst_n(i_sdma_1_rst_n),
    .sdma_1_targ_lt_Ar_Addr(sdma_1_targ_lt_axi_m_araddr_msb_fixed),
    .sdma_1_targ_lt_Ar_Burst(o_sdma_1_targ_lt_axi_m_arburst),
    .sdma_1_targ_lt_Ar_Cache(o_sdma_1_targ_lt_axi_m_arcache),
    .sdma_1_targ_lt_Ar_Id(o_sdma_1_targ_lt_axi_m_arid),
    .sdma_1_targ_lt_Ar_Len(o_sdma_1_targ_lt_axi_m_arlen),
    .sdma_1_targ_lt_Ar_Lock(o_sdma_1_targ_lt_axi_m_arlock),
    .sdma_1_targ_lt_Ar_Prot(o_sdma_1_targ_lt_axi_m_arprot),
    .sdma_1_targ_lt_Ar_Qos(o_sdma_1_targ_lt_axi_m_arqos),
    .sdma_1_targ_lt_Ar_Ready(i_sdma_1_targ_lt_axi_m_arready),
    .sdma_1_targ_lt_Ar_Size(o_sdma_1_targ_lt_axi_m_arsize),
    .sdma_1_targ_lt_Ar_Valid(o_sdma_1_targ_lt_axi_m_arvalid),
    .sdma_1_targ_lt_Aw_Addr(sdma_1_targ_lt_axi_m_awaddr_msb_fixed),
    .sdma_1_targ_lt_Aw_Burst(o_sdma_1_targ_lt_axi_m_awburst),
    .sdma_1_targ_lt_Aw_Cache(o_sdma_1_targ_lt_axi_m_awcache),
    .sdma_1_targ_lt_Aw_Id(o_sdma_1_targ_lt_axi_m_awid),
    .sdma_1_targ_lt_Aw_Len(o_sdma_1_targ_lt_axi_m_awlen),
    .sdma_1_targ_lt_Aw_Lock(o_sdma_1_targ_lt_axi_m_awlock),
    .sdma_1_targ_lt_Aw_Prot(o_sdma_1_targ_lt_axi_m_awprot),
    .sdma_1_targ_lt_Aw_Qos(o_sdma_1_targ_lt_axi_m_awqos),
    .sdma_1_targ_lt_Aw_Ready(i_sdma_1_targ_lt_axi_m_awready),
    .sdma_1_targ_lt_Aw_Size(o_sdma_1_targ_lt_axi_m_awsize),
    .sdma_1_targ_lt_Aw_Valid(o_sdma_1_targ_lt_axi_m_awvalid),
    .sdma_1_targ_lt_B_Id(i_sdma_1_targ_lt_axi_m_bid),
    .sdma_1_targ_lt_B_Ready(o_sdma_1_targ_lt_axi_m_bready),
    .sdma_1_targ_lt_B_Resp(i_sdma_1_targ_lt_axi_m_bresp),
    .sdma_1_targ_lt_B_Valid(i_sdma_1_targ_lt_axi_m_bvalid),
    .sdma_1_targ_lt_R_Data(i_sdma_1_targ_lt_axi_m_rdata),
    .sdma_1_targ_lt_R_Id(i_sdma_1_targ_lt_axi_m_rid),
    .sdma_1_targ_lt_R_Last(i_sdma_1_targ_lt_axi_m_rlast),
    .sdma_1_targ_lt_R_Ready(o_sdma_1_targ_lt_axi_m_rready),
    .sdma_1_targ_lt_R_Resp(i_sdma_1_targ_lt_axi_m_rresp),
    .sdma_1_targ_lt_R_Valid(i_sdma_1_targ_lt_axi_m_rvalid),
    .sdma_1_targ_lt_W_Data(o_sdma_1_targ_lt_axi_m_wdata),
    .sdma_1_targ_lt_W_Last(o_sdma_1_targ_lt_axi_m_wlast),
    .sdma_1_targ_lt_W_Ready(i_sdma_1_targ_lt_axi_m_wready),
    .sdma_1_targ_lt_W_Strb(o_sdma_1_targ_lt_axi_m_wstrb),
    .sdma_1_targ_lt_W_Valid(o_sdma_1_targ_lt_axi_m_wvalid),
    .sdma_1_targ_syscfg_PAddr(o_sdma_1_targ_syscfg_apb_m_paddr),
    .sdma_1_targ_syscfg_PEnable(o_sdma_1_targ_syscfg_apb_m_penable),
    .sdma_1_targ_syscfg_PProt(o_sdma_1_targ_syscfg_apb_m_pprot),
    .sdma_1_targ_syscfg_PRData(i_sdma_1_targ_syscfg_apb_m_prdata),
    .sdma_1_targ_syscfg_PReady(i_sdma_1_targ_syscfg_apb_m_pready),
    .sdma_1_targ_syscfg_PSel(o_sdma_1_targ_syscfg_apb_m_psel),
    .sdma_1_targ_syscfg_PSlvErr(i_sdma_1_targ_syscfg_apb_m_pslverr),
    .sdma_1_targ_syscfg_PStrb(o_sdma_1_targ_syscfg_apb_m_pstrb),
    .sdma_1_targ_syscfg_PWData(o_sdma_1_targ_syscfg_apb_m_pwdata),
    .sdma_1_targ_syscfg_PWrite(o_sdma_1_targ_syscfg_apb_m_pwrite)
);

endmodule
