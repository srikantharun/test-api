
// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
module ai_core
  import chip_pkg::*;
  import axi_pkg::*;
  import ai_core_pkg::*;


(

  input wire    i_clk,
  input wire    i_ref_clk,
  input wire    i_pvt_clk,
  input wire    i_rst_n,

  output  chip_axi_addr_t o_ht_axi_m_awaddr,
  output  ai_core_init_ht_axi_id_t o_ht_axi_m_awid,
  output  axi_len_t o_ht_axi_m_awlen,
  output  axi_size_t o_ht_axi_m_awsize,
  output  axi_burst_t o_ht_axi_m_awburst,
  output  axi_cache_t o_ht_axi_m_awcache,
  output  axi_prot_t o_ht_axi_m_awprot,
   output logic  o_ht_axi_m_awlock,
  output  axi_qos_t o_ht_axi_m_awqos,
  output  axi_region_t o_ht_axi_m_awregion,
  output  chip_axi_ht_awuser_t o_ht_axi_m_awuser,
   output logic  o_ht_axi_m_awvalid,
   input logic  i_ht_axi_m_awready,
  output  chip_axi_ht_data_t o_ht_axi_m_wdata,
  output  chip_axi_ht_wstrb_t o_ht_axi_m_wstrb,
   output logic  o_ht_axi_m_wlast,
  output  chip_axi_ht_wuser_t o_ht_axi_m_wuser,
   output logic  o_ht_axi_m_wvalid,
   input logic  i_ht_axi_m_wready,
   input logic  i_ht_axi_m_bvalid,
  input  ai_core_init_ht_axi_id_t i_ht_axi_m_bid,
  input  chip_axi_ht_buser_t i_ht_axi_m_buser,
  input  axi_resp_t i_ht_axi_m_bresp,
   output logic  o_ht_axi_m_bready,
  output  chip_axi_addr_t o_ht_axi_m_araddr,
  output  ai_core_init_ht_axi_id_t o_ht_axi_m_arid,
  output  axi_len_t o_ht_axi_m_arlen,
  output  axi_size_t o_ht_axi_m_arsize,
  output  axi_burst_t o_ht_axi_m_arburst,
  output  axi_cache_t o_ht_axi_m_arcache,
  output  axi_prot_t o_ht_axi_m_arprot,
  output  axi_qos_t o_ht_axi_m_arqos,
  output  axi_region_t o_ht_axi_m_arregion,
  output  chip_axi_ht_aruser_t o_ht_axi_m_aruser,
   output logic  o_ht_axi_m_arlock,
   output logic  o_ht_axi_m_arvalid,
   input logic  i_ht_axi_m_arready,
   input logic  i_ht_axi_m_rvalid,
   input logic  i_ht_axi_m_rlast,
  input  ai_core_init_ht_axi_id_t i_ht_axi_m_rid,
  input  chip_axi_ht_data_t i_ht_axi_m_rdata,
  input  chip_axi_ht_ruser_t i_ht_axi_m_ruser,
  input  axi_resp_t i_ht_axi_m_rresp,
   output logic  o_ht_axi_m_rready,
  output  chip_axi_addr_t o_lt_axi_m_awaddr,
  output  ai_core_init_lt_axi_id_t o_lt_axi_m_awid,
  output  axi_len_t o_lt_axi_m_awlen,
  output  axi_size_t o_lt_axi_m_awsize,
  output  axi_burst_t o_lt_axi_m_awburst,
  output  axi_cache_t o_lt_axi_m_awcache,
  output  axi_prot_t o_lt_axi_m_awprot,
   output logic  o_lt_axi_m_awlock,
  output  axi_qos_t o_lt_axi_m_awqos,
  output  axi_region_t o_lt_axi_m_awregion,
  output  chip_axi_lt_awuser_t o_lt_axi_m_awuser,
   output logic  o_lt_axi_m_awvalid,
   input logic  i_lt_axi_m_awready,
  output  chip_axi_lt_data_t o_lt_axi_m_wdata,
  output  chip_axi_lt_wstrb_t o_lt_axi_m_wstrb,
   output logic  o_lt_axi_m_wlast,
  output  chip_axi_lt_wuser_t o_lt_axi_m_wuser,
   output logic  o_lt_axi_m_wvalid,
   input logic  i_lt_axi_m_wready,
   input logic  i_lt_axi_m_bvalid,
  input  ai_core_init_lt_axi_id_t i_lt_axi_m_bid,
  input  chip_axi_lt_buser_t i_lt_axi_m_buser,
  input  axi_resp_t i_lt_axi_m_bresp,
   output logic  o_lt_axi_m_bready,
  output  chip_axi_addr_t o_lt_axi_m_araddr,
  output  ai_core_init_lt_axi_id_t o_lt_axi_m_arid,
  output  axi_len_t o_lt_axi_m_arlen,
  output  axi_size_t o_lt_axi_m_arsize,
  output  axi_burst_t o_lt_axi_m_arburst,
  output  axi_cache_t o_lt_axi_m_arcache,
  output  axi_prot_t o_lt_axi_m_arprot,
  output  axi_qos_t o_lt_axi_m_arqos,
  output  axi_region_t o_lt_axi_m_arregion,
  output  chip_axi_lt_aruser_t o_lt_axi_m_aruser,
   output logic  o_lt_axi_m_arlock,
   output logic  o_lt_axi_m_arvalid,
   input logic  i_lt_axi_m_arready,
   input logic  i_lt_axi_m_rvalid,
   input logic  i_lt_axi_m_rlast,
  input  ai_core_init_lt_axi_id_t i_lt_axi_m_rid,
  input  chip_axi_lt_data_t i_lt_axi_m_rdata,
  input  chip_axi_lt_ruser_t i_lt_axi_m_ruser,
  input  axi_resp_t i_lt_axi_m_rresp,
   output logic  o_lt_axi_m_rready,
  input  chip_axi_addr_t i_lt_axi_s_awaddr,
  input  ai_core_targ_lt_axi_id_t i_lt_axi_s_awid,
  input  axi_len_t i_lt_axi_s_awlen,
  input  axi_size_t i_lt_axi_s_awsize,
  input  axi_burst_t i_lt_axi_s_awburst,
  input  axi_cache_t i_lt_axi_s_awcache,
  input  axi_prot_t i_lt_axi_s_awprot,
   input logic  i_lt_axi_s_awlock,
  input  axi_qos_t i_lt_axi_s_awqos,
  input  axi_region_t i_lt_axi_s_awregion,
  input  chip_axi_lt_awuser_t i_lt_axi_s_awuser,
   input logic  i_lt_axi_s_awvalid,
   output logic  o_lt_axi_s_awready,
  input  chip_axi_lt_data_t i_lt_axi_s_wdata,
  input  chip_axi_lt_wstrb_t i_lt_axi_s_wstrb,
   input logic  i_lt_axi_s_wlast,
  input  chip_axi_lt_wuser_t i_lt_axi_s_wuser,
   input logic  i_lt_axi_s_wvalid,
   output logic  o_lt_axi_s_wready,
   output logic  o_lt_axi_s_bvalid,
  output  ai_core_targ_lt_axi_id_t o_lt_axi_s_bid,
  output  chip_axi_lt_buser_t o_lt_axi_s_buser,
  output  axi_resp_t o_lt_axi_s_bresp,
   input logic  i_lt_axi_s_bready,
  input  chip_axi_addr_t i_lt_axi_s_araddr,
  input  ai_core_targ_lt_axi_id_t i_lt_axi_s_arid,
  input  axi_len_t i_lt_axi_s_arlen,
  input  axi_size_t i_lt_axi_s_arsize,
  input  axi_burst_t i_lt_axi_s_arburst,
  input  axi_cache_t i_lt_axi_s_arcache,
  input  axi_prot_t i_lt_axi_s_arprot,
  input  axi_qos_t i_lt_axi_s_arqos,
  input  axi_region_t i_lt_axi_s_arregion,
  input  chip_axi_lt_aruser_t i_lt_axi_s_aruser,
   input logic  i_lt_axi_s_arlock,
   input logic  i_lt_axi_s_arvalid,
   output logic  o_lt_axi_s_arready,
   output logic  o_lt_axi_s_rvalid,
   output logic  o_lt_axi_s_rlast,
  output  ai_core_targ_lt_axi_id_t o_lt_axi_s_rid,
  output  chip_axi_lt_data_t o_lt_axi_s_rdata,
  output  chip_axi_lt_ruser_t o_lt_axi_s_ruser,
  output  axi_resp_t o_lt_axi_s_rresp,
   input logic  i_lt_axi_s_rready,
  input  chip_syscfg_addr_t i_cfg_apb4_s_paddr,
  input  chip_apb_syscfg_data_t i_cfg_apb4_s_pwdata,
   input logic  i_cfg_apb4_s_pwrite,
   input logic  i_cfg_apb4_s_psel,
   input logic  i_cfg_apb4_s_penable,
  input  chip_apb_syscfg_strb_t i_cfg_apb4_s_pstrb,
   input logic [3-1:0]  i_cfg_apb4_s_pprot,
   output logic  o_cfg_apb4_s_pready,
  output  chip_apb_syscfg_data_t o_cfg_apb4_s_prdata,
   output logic  o_cfg_apb4_s_pslverr,

  // DFT signals stay here temparally, they belongs to the _p wrapper file.
  // should not be in the real ai_core.sv file
  input wire    ijtag_tck,
  input wire    ssn_bus_clk,
  input wire    bisr_clk,
  input wire    ijtag_resetn,
  input wire    bisr_resetn,
  input logic    ijtag_sel,
  input logic    ijtag_ue,
  input logic    ijtag_se,
  input logic    ijtag_ce,
  input logic    ijtag_si,
  input logic    bisr_shift_en,
  input logic    bisr_si,
  input logic  [24:0] ssn_bus_data_in,
  output logic    ijtag_so,
  output logic    bisr_so,
  output logic  [24:0] ssn_bus_data_out

);

endmodule

