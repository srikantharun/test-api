
// (C) Copyright 2025 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_noc_tok_h_south
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_tok_h_south (
  input wire  i_aic_0_clk,
  input wire  i_aic_0_clken,
  input logic [7:0] i_aic_0_init_tok_ocpl_s_maddr,
  input logic [2:0] i_aic_0_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_0_init_tok_ocpl_s_mdata,
  output logic  o_aic_0_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_0_pwr_tok_idle_val,
  output logic  o_aic_0_pwr_tok_idle_ack,
  input logic  i_aic_0_pwr_tok_idle_req,
  input wire  i_aic_0_rst_n,
  output logic [7:0] o_aic_0_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_aic_0_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_0_targ_tok_ocpl_m_mdata,
  input logic  i_aic_0_targ_tok_ocpl_m_scmdaccept,
  input wire  i_aic_1_clk,
  input wire  i_aic_1_clken,
  input logic [7:0] i_aic_1_init_tok_ocpl_s_maddr,
  input logic [2:0] i_aic_1_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_1_init_tok_ocpl_s_mdata,
  output logic  o_aic_1_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_1_pwr_tok_idle_val,
  output logic  o_aic_1_pwr_tok_idle_ack,
  input logic  i_aic_1_pwr_tok_idle_req,
  input wire  i_aic_1_rst_n,
  output logic [7:0] o_aic_1_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_aic_1_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_1_targ_tok_ocpl_m_mdata,
  input logic  i_aic_1_targ_tok_ocpl_m_scmdaccept,
  input wire  i_aic_2_clk,
  input wire  i_aic_2_clken,
  input logic [7:0] i_aic_2_init_tok_ocpl_s_maddr,
  input logic [2:0] i_aic_2_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_2_init_tok_ocpl_s_mdata,
  output logic  o_aic_2_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_2_pwr_tok_idle_val,
  output logic  o_aic_2_pwr_tok_idle_ack,
  input logic  i_aic_2_pwr_tok_idle_req,
  input wire  i_aic_2_rst_n,
  output logic [7:0] o_aic_2_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_aic_2_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_2_targ_tok_ocpl_m_mdata,
  input logic  i_aic_2_targ_tok_ocpl_m_scmdaccept,
  input wire  i_aic_3_clk,
  input wire  i_aic_3_clken,
  input logic [7:0] i_aic_3_init_tok_ocpl_s_maddr,
  input logic [2:0] i_aic_3_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_3_init_tok_ocpl_s_mdata,
  output logic  o_aic_3_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_3_pwr_tok_idle_val,
  output logic  o_aic_3_pwr_tok_idle_ack,
  input logic  i_aic_3_pwr_tok_idle_req,
  input wire  i_aic_3_rst_n,
  output logic [7:0] o_aic_3_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_aic_3_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_3_targ_tok_ocpl_m_mdata,
  input logic  i_aic_3_targ_tok_ocpl_m_scmdaccept,
  input logic [31:0] i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld,
  input wire  i_noc_clk,
  input wire  i_noc_rst_n,
  input logic  scan_en
);

noc_tok_art_h_south u_noc_tok_art_h_south (
  .aic_0_clk(i_aic_0_clk),
  .aic_0_clken(i_aic_0_clken),
  .aic_0_init_tok_MAddr(i_aic_0_init_tok_ocpl_s_maddr),
  .aic_0_init_tok_MCmd(i_aic_0_init_tok_ocpl_s_mcmd),
  .aic_0_init_tok_MData(i_aic_0_init_tok_ocpl_s_mdata),
  .aic_0_init_tok_SCmdAccept(o_aic_0_init_tok_ocpl_s_scmdaccept),
  .aic_0_pwr_tok_Idle(o_aic_0_pwr_tok_idle_val),
  .aic_0_pwr_tok_IdleAck(o_aic_0_pwr_tok_idle_ack),
  .aic_0_pwr_tok_IdleReq(i_aic_0_pwr_tok_idle_req),
  .aic_0_rst_n(i_aic_0_rst_n),
  .aic_0_targ_tok_MAddr(o_aic_0_targ_tok_ocpl_m_maddr),
  .aic_0_targ_tok_MCmd(o_aic_0_targ_tok_ocpl_m_mcmd),
  .aic_0_targ_tok_MData(o_aic_0_targ_tok_ocpl_m_mdata),
  .aic_0_targ_tok_SCmdAccept(i_aic_0_targ_tok_ocpl_m_scmdaccept),
  .aic_1_clk(i_aic_1_clk),
  .aic_1_clken(i_aic_1_clken),
  .aic_1_init_tok_MAddr(i_aic_1_init_tok_ocpl_s_maddr),
  .aic_1_init_tok_MCmd(i_aic_1_init_tok_ocpl_s_mcmd),
  .aic_1_init_tok_MData(i_aic_1_init_tok_ocpl_s_mdata),
  .aic_1_init_tok_SCmdAccept(o_aic_1_init_tok_ocpl_s_scmdaccept),
  .aic_1_pwr_tok_Idle(o_aic_1_pwr_tok_idle_val),
  .aic_1_pwr_tok_IdleAck(o_aic_1_pwr_tok_idle_ack),
  .aic_1_pwr_tok_IdleReq(i_aic_1_pwr_tok_idle_req),
  .aic_1_rst_n(i_aic_1_rst_n),
  .aic_1_targ_tok_MAddr(o_aic_1_targ_tok_ocpl_m_maddr),
  .aic_1_targ_tok_MCmd(o_aic_1_targ_tok_ocpl_m_mcmd),
  .aic_1_targ_tok_MData(o_aic_1_targ_tok_ocpl_m_mdata),
  .aic_1_targ_tok_SCmdAccept(i_aic_1_targ_tok_ocpl_m_scmdaccept),
  .aic_2_clk(i_aic_2_clk),
  .aic_2_clken(i_aic_2_clken),
  .aic_2_init_tok_MAddr(i_aic_2_init_tok_ocpl_s_maddr),
  .aic_2_init_tok_MCmd(i_aic_2_init_tok_ocpl_s_mcmd),
  .aic_2_init_tok_MData(i_aic_2_init_tok_ocpl_s_mdata),
  .aic_2_init_tok_SCmdAccept(o_aic_2_init_tok_ocpl_s_scmdaccept),
  .aic_2_pwr_tok_Idle(o_aic_2_pwr_tok_idle_val),
  .aic_2_pwr_tok_IdleAck(o_aic_2_pwr_tok_idle_ack),
  .aic_2_pwr_tok_IdleReq(i_aic_2_pwr_tok_idle_req),
  .aic_2_rst_n(i_aic_2_rst_n),
  .aic_2_targ_tok_MAddr(o_aic_2_targ_tok_ocpl_m_maddr),
  .aic_2_targ_tok_MCmd(o_aic_2_targ_tok_ocpl_m_mcmd),
  .aic_2_targ_tok_MData(o_aic_2_targ_tok_ocpl_m_mdata),
  .aic_2_targ_tok_SCmdAccept(i_aic_2_targ_tok_ocpl_m_scmdaccept),
  .aic_3_clk(i_aic_3_clk),
  .aic_3_clken(i_aic_3_clken),
  .aic_3_init_tok_MAddr(i_aic_3_init_tok_ocpl_s_maddr),
  .aic_3_init_tok_MCmd(i_aic_3_init_tok_ocpl_s_mcmd),
  .aic_3_init_tok_MData(i_aic_3_init_tok_ocpl_s_mdata),
  .aic_3_init_tok_SCmdAccept(o_aic_3_init_tok_ocpl_s_scmdaccept),
  .aic_3_pwr_tok_Idle(o_aic_3_pwr_tok_idle_val),
  .aic_3_pwr_tok_IdleAck(o_aic_3_pwr_tok_idle_ack),
  .aic_3_pwr_tok_IdleReq(i_aic_3_pwr_tok_idle_req),
  .aic_3_rst_n(i_aic_3_rst_n),
  .aic_3_targ_tok_MAddr(o_aic_3_targ_tok_ocpl_m_maddr),
  .aic_3_targ_tok_MCmd(o_aic_3_targ_tok_ocpl_m_mcmd),
  .aic_3_targ_tok_MData(o_aic_3_targ_tok_ocpl_m_mdata),
  .aic_3_targ_tok_SCmdAccept(i_aic_3_targ_tok_ocpl_m_scmdaccept),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Data(i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Head(i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Rdy(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Tail(i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Vld(i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Data(i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Head(i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Rdy(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Tail(i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Vld(i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Data(o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Head(o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Rdy(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Tail(o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Vld(o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Data(o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Head(o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Rdy(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Tail(o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Vld(o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld),
  .noc_clk(i_noc_clk),
  .noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en)
);
endmodule
