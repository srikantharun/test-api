// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: Luyi <yi.lu@axelera.ai>


/// TODO:__one_line_summary_of_asic_pkg__
///
package asic_pkg;

endpackage
