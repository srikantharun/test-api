bind sys_ctrl_p Axi4PC # (
				.DATA_WIDTH(SYS_CTRL_LP_AXI_DATA_WIDTH),
                .ADDR_WIDTH(SYS_CTRL_LP_AXI_ADDR_WIDTH),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (SYS_CTRL_LP_AXI_S_ID_WIDTH),
				.WID_WIDTH  (SYS_CTRL_LP_AXI_S_ID_WIDTH),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
	      .AWREADY_MAXWAITS ( 50 ),
        .ARREADY_MAXWAITS ( 50 ),
        .WREADY_MAXWAITS ( 50 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_AIP_SYS_CTRL_LP_s_protocol_checker
				(
				.ACLK(sys_ctrl_clk_ctrl_i),
				.ARESETn(sys_ctrl_rst_no),
				.ARVALID(axi_lp_s_arvalid),
				.ARADDR(axi_lp_s_araddr ),
				.ARLEN(axi_lp_s_arlen),
				.ARSIZE( axi_lp_s_arsize),
				.ARBURST( axi_lp_s_arburst ),
				.ARLOCK( axi_lp_s_arlock),
				.ARCACHE( axi_lp_s_arcache ),
				.ARPROT( axi_lp_s_arprot ),
				.ARID( axi_lp_s_arid ),
				.ARREADY( axi_lp_s_arready ),
				.RREADY( axi_lp_s_rready ),
				.RVALID( axi_lp_s_rvalid ),
				.RLAST( axi_lp_s_rlast ),
				.RDATA(   axi_lp_s_rdata ),
				.RRESP( axi_lp_s_rresp ),
				.RID( axi_lp_s_rid ),
				.AWVALID( axi_lp_s_awvalid ),
				.AWADDR( axi_lp_s_awaddr ),
				.AWLEN( axi_lp_s_awlen),
				.AWSIZE( axi_lp_s_awsize ),
				.AWBURST( axi_lp_s_awburst ),
				.AWLOCK( axi_lp_s_awlock ),
				.AWCACHE( axi_lp_s_awcache ),
				.AWPROT( axi_lp_s_awprot ),
				.AWID( axi_lp_s_awid ),
				.AWREADY( axi_lp_s_awready ),
				.WVALID( axi_lp_s_wvalid ),
				.WLAST( axi_lp_s_wlast ),
				.WDATA(  axi_lp_s_wdata ),
				.WSTRB( axi_lp_s_wstrb ),
				.WREADY( axi_lp_s_wready),
				.BREADY( axi_lp_s_bready ),
				.BVALID( axi_lp_s_bvalid ),
				.BRESP( axi_lp_s_bresp ),
				.BID( axi_lp_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);





bind sys_ctrl_p Axi4PC # (
				.DATA_WIDTH(SYS_CTRL_LP_AXI_DATA_WIDTH),
                .ADDR_WIDTH(SYS_CTRL_LP_AXI_ADDR_WIDTH),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (SYS_CTRL_LP_AXI_M_ID_WIDTH),
				.WID_WIDTH  (SYS_CTRL_LP_AXI_M_ID_WIDTH),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
	      .AWREADY_MAXWAITS ( 50 ),
        .ARREADY_MAXWAITS ( 50 ),
        .WREADY_MAXWAITS ( 50 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_AIP_SYS_CTRL_LP_m_protocol_checker
				(
				.ACLK(sys_ctrl_clk_ctrl_i),
				.ARESETn(sys_ctrl_rst_no),
				.ARVALID(axi_lp_m_arvalid),
				.ARADDR(axi_lp_m_araddr ),
				.ARLEN(axi_lp_m_arlen),
				.ARSIZE( axi_lp_m_arsize),
				.ARBURST( axi_lp_m_arburst ),
				.ARLOCK( axi_lp_m_arlock),
				.ARCACHE( axi_lp_m_arcache ),
				.ARPROT( axi_lp_m_arprot ),
				.ARID( axi_lp_m_arid ),
				.ARREADY( axi_lp_m_arready ),
				.RREADY( axi_lp_m_rready ),
				.RVALID( axi_lp_m_rvalid ),
				.RLAST( axi_lp_m_rlast ),
				.RDATA(  axi_lp_m_rdata ),
				.RRESP( axi_lp_m_rresp ),
				.RID( axi_lp_m_rid ),
				.AWVALID( axi_lp_m_awvalid ),
				.AWADDR( axi_lp_m_awaddr ),
				.AWLEN( axi_lp_m_awlen),
				.AWSIZE( axi_lp_m_awsize ),
				.AWBURST( axi_lp_m_awburst ),
				.AWLOCK( axi_lp_m_awlock ),
				.AWCACHE( axi_lp_m_awcache ),
				.AWPROT( axi_lp_m_awprot ),
				.AWID( axi_lp_m_awid ),
				.AWREADY( axi_lp_m_awready ),
				.WVALID( axi_lp_m_wvalid ),
				.WLAST( axi_lp_m_wlast ),
				.WDATA(  axi_lp_m_wdata ),
				.WSTRB( axi_lp_m_wstrb ),
				.WREADY( axi_lp_m_wready),
				.BREADY( axi_lp_m_bready ),
				.BVALID( axi_lp_m_bvalid ),
				.BRESP( axi_lp_m_bresp ),
				.BID( axi_lp_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);


bind sys_ctrl_p Axi4PC # (
				.DATA_WIDTH(SYS_DMA_HP_AXI_DATA_WIDTH),
                .ADDR_WIDTH(SYS_DMA_HP_AXI_ADDR_WIDTH),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (SYS_DMA_HP_AXI_ID_WIDTH),
				.WID_WIDTH  (SYS_DMA_HP_AXI_ID_WIDTH),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
      	.AWREADY_MAXWAITS ( 50 ),
        .ARREADY_MAXWAITS ( 50 ),
        .WREADY_MAXWAITS ( 50 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_AIP_SYS_CTRL_hp_dma_0_protocol_checker
				(
				.ACLK(sys_ctrl_clk_ctrl_i),
				.ARESETn(dma_rst_no),
				.ARVALID(sys_dma_0_axi_hp_m_arvalid),
				.ARADDR(sys_dma_0_axi_hp_m_araddr ),
				.ARLEN(sys_dma_0_axi_hp_m_arlen),
				.ARSIZE( sys_dma_0_axi_hp_m_arsize),
				.ARBURST( sys_dma_0_axi_hp_m_arburst ),
				.ARLOCK( sys_dma_0_axi_hp_m_arlock),
				.ARCACHE( sys_dma_0_axi_hp_m_arcache ),
				.ARPROT( sys_dma_0_axi_hp_m_arprot ),
				.ARID( sys_dma_0_axi_hp_m_arid ),
				.ARREADY( sys_dma_0_axi_hp_m_arready ),
				.RREADY( sys_dma_0_axi_hp_m_rready ),
				.RVALID( sys_dma_0_axi_hp_m_rvalid ),
				.RLAST( sys_dma_0_axi_hp_m_rlast ),
				.RDATA(  sys_dma_0_axi_hp_m_rdata ),
				.RRESP( sys_dma_0_axi_hp_m_rresp ),
				.RID( sys_dma_0_axi_hp_m_rid ),
				.AWVALID( sys_dma_0_axi_hp_m_awvalid ),
				.AWADDR( sys_dma_0_axi_hp_m_awaddr ),
				.AWLEN( sys_dma_0_axi_hp_m_awlen),
				.AWSIZE( sys_dma_0_axi_hp_m_awsize ),
				.AWBURST( sys_dma_0_axi_hp_m_awburst ),
				.AWLOCK( sys_dma_0_axi_hp_m_awlock ),
				.AWCACHE( sys_dma_0_axi_hp_m_awcache ),
				.AWPROT( sys_dma_0_axi_hp_m_awprot ),
				.AWID( sys_dma_0_axi_hp_m_awid ),
				.AWREADY( sys_dma_0_axi_hp_m_awready ),
				.WVALID( sys_dma_0_axi_hp_m_wvalid ),
				.WLAST( sys_dma_0_axi_hp_m_wlast ),
				.WDATA(  sys_dma_0_axi_hp_m_wdata ),
				.WSTRB( sys_dma_0_axi_hp_m_wstrb ),
				.WREADY( sys_dma_0_axi_hp_m_wready),
				.BREADY( sys_dma_0_axi_hp_m_bready ),
				.BVALID( sys_dma_0_axi_hp_m_bvalid ),
				.BRESP( sys_dma_0_axi_hp_m_bresp ),
				.BID( sys_dma_0_axi_hp_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);



bind sys_ctrl_p Axi4PC # (
				.DATA_WIDTH(SYS_DMA_HP_AXI_DATA_WIDTH),
                .ADDR_WIDTH(SYS_DMA_HP_AXI_ADDR_WIDTH),
				//.ID_WIDTH  (`DW_VIP_AXI_AID_PORT_WIDTH),
				.RID_WIDTH  (SYS_DMA_HP_AXI_ID_WIDTH),
				.WID_WIDTH  (SYS_DMA_HP_AXI_ID_WIDTH),
                .MAXWBURSTS(20),
                .MAXRBURSTS(20),
                .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
	      .AWREADY_MAXWAITS ( 50 ),
        .ARREADY_MAXWAITS ( 50 ),
        .WREADY_MAXWAITS ( 50 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_AIP_SYS_CTRL_hp_dma_1_protocol_checker
				(
				.ACLK(sys_ctrl_clk_ctrl_i),
				.ARESETn(dma_rst_no),
				.ARVALID(sys_dma_1_axi_hp_m_arvalid),
				.ARADDR(sys_dma_1_axi_hp_m_araddr ),
				.ARLEN(sys_dma_1_axi_hp_m_arlen),
				.ARSIZE( sys_dma_1_axi_hp_m_arsize),
				.ARBURST( sys_dma_1_axi_hp_m_arburst ),
				.ARLOCK( sys_dma_1_axi_hp_m_arlock),
				.ARCACHE( sys_dma_1_axi_hp_m_arcache ),
				.ARPROT( sys_dma_1_axi_hp_m_arprot ),
				.ARID( sys_dma_1_axi_hp_m_arid ),
				.ARREADY( sys_dma_1_axi_hp_m_arready ),
				.RREADY( sys_dma_1_axi_hp_m_rready ),
				.RVALID( sys_dma_1_axi_hp_m_rvalid ),
				.RLAST( sys_dma_1_axi_hp_m_rlast ),
				.RDATA(  sys_dma_1_axi_hp_m_rdata ),
				.RRESP( sys_dma_1_axi_hp_m_rresp ),
				.RID( sys_dma_1_axi_hp_m_rid ),
				.AWVALID( sys_dma_1_axi_hp_m_awvalid ),
				.AWADDR( sys_dma_1_axi_hp_m_awaddr ),
				.AWLEN( sys_dma_1_axi_hp_m_awlen),
				.AWSIZE( sys_dma_1_axi_hp_m_awsize ),
				.AWBURST( sys_dma_1_axi_hp_m_awburst ),
				.AWLOCK( sys_dma_1_axi_hp_m_awlock ),
				.AWCACHE( sys_dma_1_axi_hp_m_awcache ),
				.AWPROT( sys_dma_1_axi_hp_m_awprot ),
				.AWID( sys_dma_1_axi_hp_m_awid ),
				.AWREADY( sys_dma_1_axi_hp_m_awready ),
				.WVALID( sys_dma_1_axi_hp_m_wvalid ),
				.WLAST( sys_dma_1_axi_hp_m_wlast ),
				.WDATA(  sys_dma_1_axi_hp_m_wdata ),
				.WSTRB( sys_dma_1_axi_hp_m_wstrb ),
				.WREADY( sys_dma_1_axi_hp_m_wready),
				.BREADY( sys_dma_1_axi_hp_m_bready ),
				.BVALID( sys_dma_1_axi_hp_m_bvalid ),
				.BRESP( sys_dma_1_axi_hp_m_bresp ),
				.BID( sys_dma_1_axi_hp_m_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER(32'h0),  .AWREGION(4'b0) , .AWQOS(4'b0) , .ARQOS(4'b0), .ARREGION(4'b0),.CACTIVE(1'b0),.CSYSREQ(1'b0),.CSYSACK(1'b0)
				);

