
package allegro_tb_uvm_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import decoder_uvm_pkg::*;

  `include "allegro_tb_demoter.svh"
  `include "allegro_tb_test.svh"

endpackage : allegro_tb_uvm_pkg
