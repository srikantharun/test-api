
// (C) Copyright 2025 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_noc_tok_soc
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_tok_soc (
  input logic [7:0] i_apu_init_tok_ocpl_s_maddr,
  input logic [2:0] i_apu_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_apu_init_tok_ocpl_s_mdata,
  output logic  o_apu_init_tok_ocpl_s_scmdaccept,
  output logic  o_apu_pwr_tok_idle_val,
  output logic  o_apu_pwr_tok_idle_ack,
  input logic  i_apu_pwr_tok_idle_req,
  output logic [7:0] o_apu_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_apu_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_apu_targ_tok_ocpl_m_mdata,
  input logic  i_apu_targ_tok_ocpl_m_scmdaccept,
  input wire  i_apu_x_clk,
  input wire  i_apu_x_clken,
  input wire  i_apu_x_rst_n,
  input logic [41:0] i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld,
  input wire  i_noc_clk,
  input wire  i_noc_rst_n,
  input logic  scan_en
);

noc_tok_art_soc u_noc_tok_art_soc (
  .apu_init_tok_MAddr(i_apu_init_tok_ocpl_s_maddr),
  .apu_init_tok_MCmd(i_apu_init_tok_ocpl_s_mcmd),
  .apu_init_tok_MData(i_apu_init_tok_ocpl_s_mdata),
  .apu_init_tok_SCmdAccept(o_apu_init_tok_ocpl_s_scmdaccept),
  .apu_pwr_tok_Idle(o_apu_pwr_tok_idle_val),
  .apu_pwr_tok_IdleAck(o_apu_pwr_tok_idle_ack),
  .apu_pwr_tok_IdleReq(i_apu_pwr_tok_idle_req),
  .apu_targ_tok_MAddr(o_apu_targ_tok_ocpl_m_maddr),
  .apu_targ_tok_MCmd(o_apu_targ_tok_ocpl_m_mcmd),
  .apu_targ_tok_MData(o_apu_targ_tok_ocpl_m_mdata),
  .apu_targ_tok_SCmdAccept(i_apu_targ_tok_ocpl_m_scmdaccept),
  .apu_x_clk(i_apu_x_clk),
  .apu_x_clken(i_apu_x_clken),
  .apu_x_rst_n(i_apu_x_rst_n),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Data(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Head(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Rdy(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Tail(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Vld(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Data(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Head(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Rdy(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Tail(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Vld(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Data(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Head(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Rdy(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Tail(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Vld(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Data(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Head(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Rdy(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Tail(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Vld(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld),
  .noc_clk(i_noc_clk),
  .noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en)
);
endmodule
