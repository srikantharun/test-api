// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Derived address map for AI Core with local addresses that can be used by IPs
// Owner: Sander Geursen <sander.geursen@axelera.ai>

`ifndef AIC_ADDR_MAP_PKG_SV
`define AIC_ADDR_MAP_PKG_SV

package aic_addr_map_pkg;
  import aipu_addr_map_pkg::*;

  parameter int unsigned AIC_AXI_LT_LOCAL_ADDR_WIDTH = 28;

  typedef logic [chip_pkg::CHIP_AXI_ADDR_W-1:0]   ext_addr_t;
  typedef logic [AIC_AXI_LT_LOCAL_ADDR_WIDTH-1:0] loc_addr_t;

  ////////////////////////
  ///  Datapath regions:
  parameter ext_addr_t AIC_DP_CSR_ST_ADDR   = AICORE_0_DATAPATH_CSR_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_DP_CSR_END_ADDR  = AICORE_0_DATAPATH_CSR_DID_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_DP_CMD_ST_ADDR   = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_DP_CMD_END_ADDR  = AICORE_0_DATAPATH_COMMAND_DID_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_DP_PRG_ST_ADDR   = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_DP_PRG_END_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_DID_RESERVED_END_ADDR;

  parameter ext_addr_t AIC_DP_ALL_ST_ADDR   = AIC_DP_CSR_ST_ADDR;
  parameter ext_addr_t AIC_DP_ALL_END_ADDR  = AIC_DP_PRG_END_ADDR;


  ///////////////////////////////////////////////////////////
  // external addresses for specific devices:
  parameter ext_addr_t AIC_CFG_CSR_INFRA_PART_ST_ADDR  = AICORE_0_CONFIGURATION_PERIPHERALS_CSR_INFRA_ST_ADDR;
  parameter ext_addr_t AIC_CFG_CSR_INFRA_PART_END_ADDR = AICORE_0_CONFIGURATION_PERIPHERALS_CSR_INFRA_END_ADDR;
  parameter ext_addr_t AIC_CFG_CSR_MID_PART_ST_ADDR    = AICORE_0_CONFIGURATION_PERIPHERALS_CSR_MID_ST_ADDR;
  parameter ext_addr_t AIC_CFG_CSR_MID_PART_END_ADDR   = AICORE_0_CONFIGURATION_PERIPHERALS_CSR_MID_END_ADDR;
  parameter ext_addr_t AIC_CFG_MAILBOX_ST_ADDR         = AICORE_0_CONFIGURATION_PERIPHERALS_MAILBOX_ST_ADDR;
  parameter ext_addr_t AIC_CFG_MAILBOX_END_ADDR        = AICORE_0_CONFIGURATION_PERIPHERALS_MAILBOX_END_ADDR;
  parameter ext_addr_t AIC_CFG_TOK_MGR_ST_ADDR         = AICORE_0_CONFIGURATION_PERIPHERALS_TOKEN_MANAGER_ST_ADDR;
  parameter ext_addr_t AIC_CFG_TOK_MGR_END_ADDR        = AICORE_0_CONFIGURATION_PERIPHERALS_TOKEN_MANAGER_END_ADDR;
  parameter ext_addr_t AIC_CFG_PLIC_ST_ADDR            = AICORE_0_CONFIGURATION_PERIPHERALS_PLIC_ST_ADDR;
  parameter ext_addr_t AIC_CFG_PLIC_END_ADDR           = AICORE_0_CONFIGURATION_PERIPHERALS_PLIC_END_ADDR;
  parameter ext_addr_t AIC_CFG_TIMESTAMP_CSR_ST_ADDR   = AICORE_0_CONFIGURATION_PERIPHERALS_TIMESTAMP_UNIT_CSR_ST_ADDR;
  parameter ext_addr_t AIC_CFG_TIMESTAMP_CSR_END_ADDR  = AICORE_0_CONFIGURATION_PERIPHERALS_TIMESTAMP_UNIT_CSR_END_ADDR;
  parameter ext_addr_t AIC_CFG_TIMESTAMP_MEM_ST_ADDR   = AICORE_0_CONFIGURATION_PERIPHERALS_TIMESTAMP_UNIT_MEM_ST_ADDR;
  parameter ext_addr_t AIC_CFG_TIMESTAMP_MEM_END_ADDR  = AICORE_0_CONFIGURATION_PERIPHERALS_TIMESTAMP_UNIT_MEM_END_ADDR;
  parameter ext_addr_t AIC_CFG_TIMESTAMP_ST_ADDR       = AIC_CFG_TIMESTAMP_CSR_ST_ADDR;
  parameter ext_addr_t AIC_CFG_TIMESTAMP_END_ADDR      = AIC_CFG_TIMESTAMP_MEM_END_ADDR;

  parameter ext_addr_t AIC_CFG_ACD_CSR_ST_ADDR         = AICORE_0_CONFIGURATION_CONTROL_ACD_CSR_ST_ADDR;
  parameter ext_addr_t AIC_CFG_ACD_CSR_END_ADDR        = AICORE_0_CONFIGURATION_CONTROL_ACD_CSR_END_ADDR;
  parameter ext_addr_t AIC_CFG_ACD_CMD_ST_ADDR         = AICORE_0_CONFIGURATION_CONTROL_ACD_COMMAND_ST_ADDR;
  parameter ext_addr_t AIC_CFG_ACD_CMD_END_ADDR        = AICORE_0_CONFIGURATION_CONTROL_ACD_COMMAND_END_ADDR;
  parameter ext_addr_t AIC_CFG_ACD_ST_ADDR             = AIC_CFG_ACD_CSR_ST_ADDR;
  parameter ext_addr_t AIC_CFG_ACD_END_ADDR            = AIC_CFG_ACD_CMD_END_ADDR;
  parameter ext_addr_t AIC_CFG_LP_DMA_ST_ADDR          = AICORE_0_CONFIGURATION_CONTROL_LP_DMA_ST_ADDR;
  parameter ext_addr_t AIC_CFG_LP_DMA_END_ADDR         = AICORE_0_CONFIGURATION_CONTROL_LP_DMA_END_ADDR;

  parameter ext_addr_t AIC_SPM_ST_ADDR                 = AICORE_0_SPM_ST_ADDR;
  parameter ext_addr_t AIC_SPM_END_ADDR                = AICORE_0_SPM_END_ADDR;
  parameter ext_addr_t AIC_L1_ST_ADDR                  = AICORE_0_L1_ST_ADDR;
  parameter ext_addr_t AIC_L1_END_ADDR                 = AICORE_0_L1_END_ADDR;

  parameter ext_addr_t AIC_CFG_PERIPH_ST_ADDR          = AICORE_0_CONFIGURATION_PERIPHERALS_MAILBOX_ST_ADDR;
  parameter ext_addr_t AIC_CFG_PERIPH_END_ADDR         = AICORE_0_CONFIGURATION_PERIPHERALS_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_CFG_CTRL_ST_ADDR            = AICORE_0_CONFIGURATION_CONTROL_ACD_CSR_ST_ADDR;
  parameter ext_addr_t AIC_CFG_CTRL_END_ADDR           = AICORE_0_CONFIGURATION_CONTROL_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_CFG_ST_ADDR                 = AIC_CFG_PERIPH_ST_ADDR;
  parameter ext_addr_t AIC_CFG_END_ADDR                = AICORE_0_CONFIGURATION_CONTROL_RESERVED_END_ADDR;

  // local addresses for specific devices, that need a local version:
  parameter loc_addr_t AIC_LOC_CFG_CSR_INFRA_PART_ST_ADDR  = AIC_CFG_CSR_INFRA_PART_ST_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_CSR_INFRA_PART_END_ADDR = AIC_CFG_CSR_INFRA_PART_END_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_CSR_MID_PART_ST_ADDR    = AIC_CFG_CSR_MID_PART_ST_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_CSR_MID_PART_END_ADDR   = AIC_CFG_CSR_MID_PART_END_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_TIMESTAMP_CSR_ST_ADDR   = AIC_CFG_TIMESTAMP_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_TIMESTAMP_CSR_END_ADDR  = AIC_CFG_TIMESTAMP_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_TIMESTAMP_MEM_ST_ADDR   = AIC_CFG_TIMESTAMP_MEM_ST_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_TIMESTAMP_MEM_END_ADDR  = AIC_CFG_TIMESTAMP_MEM_END_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_ACD_CSR_ST_ADDR         = AIC_CFG_ACD_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_ACD_CSR_END_ADDR        = AIC_CFG_ACD_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_ACD_CMD_ST_ADDR         = AIC_CFG_ACD_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_CFG_ACD_CMD_END_ADDR        = AIC_CFG_ACD_CMD_END_ADDR;


  // external addresses for datapath devices:
    // Devices:
    // M_IFD0
  parameter ext_addr_t AIC_M_IFD_0_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_0_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_M_IFD_0_END_ADDR;
  parameter ext_addr_t AIC_M_IFD_0_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_0_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_0_END_ADDR;
  parameter ext_addr_t AIC_M_IFD_0_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_0_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_0_END_ADDR;
    // M_IFD1
  parameter ext_addr_t AIC_M_IFD_1_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_M_IFD_1_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_1_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_M_IFD_1_END_ADDR;
  parameter ext_addr_t AIC_M_IFD_1_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_1_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_1_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_1_END_ADDR;
  parameter ext_addr_t AIC_M_IFD_1_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_1_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_1_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_1_END_ADDR;
    // M_IFD2
  parameter ext_addr_t AIC_M_IFD_2_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_M_IFD_2_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_2_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_M_IFD_2_END_ADDR;
  parameter ext_addr_t AIC_M_IFD_2_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_2_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_2_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_2_END_ADDR;
  parameter ext_addr_t AIC_M_IFD_2_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_2_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_2_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_2_END_ADDR;
    // M_IFDW
  parameter ext_addr_t AIC_M_IFD_W_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_M_IFD_W_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_W_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_M_IFD_W_END_ADDR;
  parameter ext_addr_t AIC_M_IFD_W_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_W_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_W_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_W_END_ADDR;
  parameter ext_addr_t AIC_M_IFD_W_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_W_ST_ADDR;
  parameter ext_addr_t AIC_M_IFD_W_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_W_END_ADDR;
    // M_ODR
  parameter ext_addr_t AIC_M_ODR_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_M_ODR_ST_ADDR;
  parameter ext_addr_t AIC_M_ODR_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_M_ODR_END_ADDR;
  parameter ext_addr_t AIC_M_ODR_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_M_ODR_ST_ADDR;
  parameter ext_addr_t AIC_M_ODR_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_M_ODR_END_ADDR;
  parameter ext_addr_t AIC_M_ODR_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_ODR_ST_ADDR;
  parameter ext_addr_t AIC_M_ODR_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_ODR_END_ADDR;
    // D_IFD0
  parameter ext_addr_t AIC_D_IFD_0_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_D_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_D_IFD_0_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_D_IFD_0_END_ADDR;
  parameter ext_addr_t AIC_D_IFD_0_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_D_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_D_IFD_0_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_D_IFD_0_END_ADDR;
  parameter ext_addr_t AIC_D_IFD_0_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_D_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_D_IFD_0_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_D_IFD_0_END_ADDR;
    // D_IFD1
  parameter ext_addr_t AIC_D_IFD_1_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_D_IFD_1_ST_ADDR;
  parameter ext_addr_t AIC_D_IFD_1_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_D_IFD_1_END_ADDR;
  parameter ext_addr_t AIC_D_IFD_1_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_D_IFD_1_ST_ADDR;
  parameter ext_addr_t AIC_D_IFD_1_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_D_IFD_1_END_ADDR;
  parameter ext_addr_t AIC_D_IFD_1_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_D_IFD_1_ST_ADDR;
  parameter ext_addr_t AIC_D_IFD_1_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_D_IFD_1_END_ADDR;
    // D_ODR
  parameter ext_addr_t AIC_D_ODR_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_D_ODR_ST_ADDR;
  parameter ext_addr_t AIC_D_ODR_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_D_ODR_END_ADDR;
  parameter ext_addr_t AIC_D_ODR_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_D_ODR_ST_ADDR;
  parameter ext_addr_t AIC_D_ODR_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_D_ODR_END_ADDR;
  parameter ext_addr_t AIC_D_ODR_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_D_ODR_ST_ADDR;
  parameter ext_addr_t AIC_D_ODR_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_D_ODR_END_ADDR;

    // M_MVM_EXE
  parameter ext_addr_t AIC_M_MVM_EXE_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_MID_M_MVMEXE_ST_ADDR;
  parameter ext_addr_t AIC_M_MVM_EXE_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_MID_M_MVMEXE_END_ADDR;
  parameter ext_addr_t AIC_M_MVM_EXE_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_MID_M_MVMEXE_ST_ADDR;
  parameter ext_addr_t AIC_M_MVM_EXE_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_MID_M_MVMEXE_END_ADDR;
  parameter ext_addr_t AIC_M_MVM_EXE_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_MVMEXE_ST_ADDR;
  parameter ext_addr_t AIC_M_MVM_EXE_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_MVMEXE_END_ADDR;
    // M_MVM_PRG
  parameter ext_addr_t AIC_M_MVM_PRG_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_MID_M_MVMPRG_ST_ADDR;
  parameter ext_addr_t AIC_M_MVM_PRG_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_MID_M_MVMPRG_END_ADDR;
  parameter ext_addr_t AIC_M_MVM_PRG_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_MID_M_MVMPRG_ST_ADDR;
  parameter ext_addr_t AIC_M_MVM_PRG_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_MID_M_MVMPRG_END_ADDR;
  parameter ext_addr_t AIC_M_MVM_PRG_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_MVMPRG_ST_ADDR;
  parameter ext_addr_t AIC_M_MVM_PRG_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_MVMPRG_END_ADDR;
    // M_IAU
  parameter ext_addr_t AIC_M_IAU_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_MID_M_IAU_ST_ADDR;
  parameter ext_addr_t AIC_M_IAU_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_MID_M_IAU_END_ADDR;
  parameter ext_addr_t AIC_M_IAU_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_MID_M_IAU_ST_ADDR;
  parameter ext_addr_t AIC_M_IAU_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_MID_M_IAU_END_ADDR;
  parameter ext_addr_t AIC_M_IAU_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_IAU_ST_ADDR;
  parameter ext_addr_t AIC_M_IAU_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_IAU_END_ADDR;
    // M_DPU
  parameter ext_addr_t AIC_M_DPU_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_MID_M_DPU_ST_ADDR;
  parameter ext_addr_t AIC_M_DPU_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_MID_M_DPU_END_ADDR;
  parameter ext_addr_t AIC_M_DPU_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_MID_M_DPU_ST_ADDR;
  parameter ext_addr_t AIC_M_DPU_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_MID_M_DPU_END_ADDR;
  parameter ext_addr_t AIC_M_DPU_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_DPU_ST_ADDR;
  parameter ext_addr_t AIC_M_DPU_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_DPU_END_ADDR;
    // D_DWPU
  parameter ext_addr_t AIC_D_DWPU_CSR_ST_ADDR  =AICORE_0_DATAPATH_CSR_DID_D_DWPU_ST_ADDR;
  parameter ext_addr_t AIC_D_DWPU_CSR_END_ADDR =AICORE_0_DATAPATH_CSR_DID_D_DWPU_END_ADDR;
  parameter ext_addr_t AIC_D_DWPU_CMD_ST_ADDR  =AICORE_0_DATAPATH_COMMAND_DID_D_DWPU_ST_ADDR;
  parameter ext_addr_t AIC_D_DWPU_CMD_END_ADDR =AICORE_0_DATAPATH_COMMAND_DID_D_DWPU_END_ADDR;
  parameter ext_addr_t AIC_D_DWPU_PRG_ST_ADDR  =AICORE_0_DATAPATH_INSTRUCTIONS_DID_D_DWPU_ST_ADDR;
  parameter ext_addr_t AIC_D_DWPU_PRG_END_ADDR =AICORE_0_DATAPATH_INSTRUCTIONS_DID_D_DWPU_END_ADDR;
    // D_IAU
  parameter ext_addr_t AIC_D_IAU_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_DID_D_IAU_ST_ADDR;
  parameter ext_addr_t AIC_D_IAU_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_DID_D_IAU_END_ADDR;
  parameter ext_addr_t AIC_D_IAU_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_DID_D_IAU_ST_ADDR;
  parameter ext_addr_t AIC_D_IAU_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_DID_D_IAU_END_ADDR;
  parameter ext_addr_t AIC_D_IAU_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_DID_D_IAU_ST_ADDR;
  parameter ext_addr_t AIC_D_IAU_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_DID_D_IAU_END_ADDR;
    // D_DPU
  parameter ext_addr_t AIC_D_DPU_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_DID_D_DPU_ST_ADDR;
  parameter ext_addr_t AIC_D_DPU_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_DID_D_DPU_END_ADDR;
  parameter ext_addr_t AIC_D_DPU_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_DID_D_DPU_ST_ADDR;
  parameter ext_addr_t AIC_D_DPU_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_DID_D_DPU_END_ADDR;
  parameter ext_addr_t AIC_D_DPU_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_DID_D_DPU_ST_ADDR;
  parameter ext_addr_t AIC_D_DPU_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_DID_D_DPU_END_ADDR;

    // HP_DMA common parts
  parameter ext_addr_t AIC_HP_DMA_MMU_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_DMA_MMU_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_MMU_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_DMA_MMU_END_ADDR;
  parameter ext_addr_t AIC_HP_DMA_COMMON_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_DMA_COMMON_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_COMMON_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_DMA_COMMON_END_ADDR;

    // HP_DMA_0
  parameter ext_addr_t AIC_HP_DMA_0_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_DMA_HP_DMA_0_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_0_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_DMA_HP_DMA_0_END_ADDR;
  parameter ext_addr_t AIC_HP_DMA_0_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_DMA_HP_DMA_0_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_0_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_DMA_HP_DMA_0_END_ADDR;
  parameter ext_addr_t AIC_HP_DMA_0_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_DMA_HP_DMA_0_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_0_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_DMA_HP_DMA_0_END_ADDR;
    // HP_DMA_1
  parameter ext_addr_t AIC_HP_DMA_1_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_DMA_HP_DMA_1_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_1_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_DMA_HP_DMA_1_END_ADDR;
  parameter ext_addr_t AIC_HP_DMA_1_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_DMA_HP_DMA_1_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_1_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_DMA_HP_DMA_1_END_ADDR;
  parameter ext_addr_t AIC_HP_DMA_1_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_DMA_HP_DMA_1_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_1_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_DMA_HP_DMA_1_END_ADDR;

  ///////////////////////////////////////////////////////////
  // local addresses for datapath devices:
    // Devices:
    // M_IFD0
  parameter loc_addr_t AIC_LOC_M_IFD_0_CSR_ST_ADDR  = AIC_M_IFD_0_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_0_CSR_END_ADDR = AIC_M_IFD_0_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_0_CMD_ST_ADDR  = AIC_M_IFD_0_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_0_CMD_END_ADDR = AIC_M_IFD_0_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_0_PRG_ST_ADDR  = AIC_M_IFD_0_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_0_PRG_END_ADDR = AIC_M_IFD_0_PRG_END_ADDR;
    // M_IFD1
  parameter loc_addr_t AIC_LOC_M_IFD_1_CSR_ST_ADDR  = AIC_M_IFD_1_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_1_CSR_END_ADDR = AIC_M_IFD_1_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_1_CMD_ST_ADDR  = AIC_M_IFD_1_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_1_CMD_END_ADDR = AIC_M_IFD_1_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_1_PRG_ST_ADDR  = AIC_M_IFD_1_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_1_PRG_END_ADDR = AIC_M_IFD_1_PRG_END_ADDR;
    // M_IFD2
  parameter loc_addr_t AIC_LOC_M_IFD_2_CSR_ST_ADDR  = AIC_M_IFD_2_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_2_CSR_END_ADDR = AIC_M_IFD_2_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_2_CMD_ST_ADDR  = AIC_M_IFD_2_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_2_CMD_END_ADDR = AIC_M_IFD_2_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_2_PRG_ST_ADDR  = AIC_M_IFD_2_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_2_PRG_END_ADDR = AIC_M_IFD_2_PRG_END_ADDR;
    // M_IFDW
  parameter loc_addr_t AIC_LOC_M_IFD_W_CSR_ST_ADDR  = AIC_M_IFD_W_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_W_CSR_END_ADDR = AIC_M_IFD_W_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_W_CMD_ST_ADDR  = AIC_M_IFD_W_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_W_CMD_END_ADDR = AIC_M_IFD_W_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_W_PRG_ST_ADDR  = AIC_M_IFD_W_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IFD_W_PRG_END_ADDR = AIC_M_IFD_W_PRG_END_ADDR;
    // M_ODR
  parameter loc_addr_t AIC_LOC_M_ODR_CSR_ST_ADDR  = AIC_M_ODR_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_ODR_CSR_END_ADDR = AIC_M_ODR_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_ODR_CMD_ST_ADDR  = AIC_M_ODR_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_ODR_CMD_END_ADDR = AIC_M_ODR_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_ODR_PRG_ST_ADDR  = AIC_M_ODR_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_ODR_PRG_END_ADDR = AIC_M_ODR_PRG_END_ADDR;
    // D_IFD0
  parameter loc_addr_t AIC_LOC_D_IFD_0_CSR_ST_ADDR  = AIC_D_IFD_0_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_0_CSR_END_ADDR = AIC_D_IFD_0_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_0_CMD_ST_ADDR  = AIC_D_IFD_0_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_0_CMD_END_ADDR = AIC_D_IFD_0_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_0_PRG_ST_ADDR  = AIC_D_IFD_0_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_0_PRG_END_ADDR = AIC_D_IFD_0_PRG_END_ADDR;
    // D_IFD1
  parameter loc_addr_t AIC_LOC_D_IFD_1_CSR_ST_ADDR  = AIC_D_IFD_1_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_1_CSR_END_ADDR = AIC_D_IFD_1_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_1_CMD_ST_ADDR  = AIC_D_IFD_1_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_1_CMD_END_ADDR = AIC_D_IFD_1_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_1_PRG_ST_ADDR  = AIC_D_IFD_1_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IFD_1_PRG_END_ADDR = AIC_D_IFD_1_PRG_END_ADDR;
    // D_ODR
  parameter loc_addr_t AIC_LOC_D_ODR_CSR_ST_ADDR  = AIC_D_ODR_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_ODR_CSR_END_ADDR = AIC_D_ODR_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_ODR_CMD_ST_ADDR  = AIC_D_ODR_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_ODR_CMD_END_ADDR = AIC_D_ODR_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_ODR_PRG_ST_ADDR  = AIC_D_ODR_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_ODR_PRG_END_ADDR = AIC_D_ODR_PRG_END_ADDR;
    // M_MVM_EXE
  parameter loc_addr_t AIC_LOC_M_MVM_EXE_CSR_ST_ADDR  = AIC_M_MVM_EXE_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_EXE_CSR_END_ADDR = AIC_M_MVM_EXE_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_EXE_CMD_ST_ADDR  = AIC_M_MVM_EXE_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_EXE_CMD_END_ADDR = AIC_M_MVM_EXE_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_EXE_PRG_ST_ADDR  = AIC_M_MVM_EXE_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_EXE_PRG_END_ADDR = AIC_M_MVM_EXE_PRG_END_ADDR;
    // M_MVM_PRG
  parameter loc_addr_t AIC_LOC_M_MVM_PRG_CSR_ST_ADDR  = AIC_M_MVM_PRG_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_PRG_CSR_END_ADDR = AIC_M_MVM_PRG_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_PRG_CMD_ST_ADDR  = AIC_M_MVM_PRG_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_PRG_CMD_END_ADDR = AIC_M_MVM_PRG_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_PRG_PRG_ST_ADDR  = AIC_M_MVM_PRG_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_MVM_PRG_PRG_END_ADDR = AIC_M_MVM_PRG_PRG_END_ADDR;
    // M_IAU
  parameter loc_addr_t AIC_LOC_M_IAU_CSR_ST_ADDR  = AIC_M_IAU_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IAU_CSR_END_ADDR = AIC_M_IAU_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IAU_CMD_ST_ADDR  = AIC_M_IAU_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IAU_CMD_END_ADDR = AIC_M_IAU_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_IAU_PRG_ST_ADDR  = AIC_M_IAU_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_IAU_PRG_END_ADDR = AIC_M_IAU_PRG_END_ADDR;
    // M_DPU
  parameter loc_addr_t AIC_LOC_M_DPU_CSR_ST_ADDR  = AIC_M_DPU_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_DPU_CSR_END_ADDR = AIC_M_DPU_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_DPU_CMD_ST_ADDR  = AIC_M_DPU_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_DPU_CMD_END_ADDR = AIC_M_DPU_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_M_DPU_PRG_ST_ADDR  = AIC_M_DPU_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_M_DPU_PRG_END_ADDR = AIC_M_DPU_PRG_END_ADDR;
    // D_DWPU
  parameter loc_addr_t AIC_LOC_D_DWPU_CSR_ST_ADDR  = AIC_D_DWPU_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_DWPU_CSR_END_ADDR = AIC_D_DWPU_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_DWPU_CMD_ST_ADDR  = AIC_D_DWPU_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_DWPU_CMD_END_ADDR = AIC_D_DWPU_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_DWPU_PRG_ST_ADDR  = AIC_D_DWPU_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_DWPU_PRG_END_ADDR = AIC_D_DWPU_PRG_END_ADDR;
    // D_IAU
  parameter loc_addr_t AIC_LOC_D_IAU_CSR_ST_ADDR  = AIC_D_IAU_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IAU_CSR_END_ADDR = AIC_D_IAU_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_IAU_CMD_ST_ADDR  = AIC_D_IAU_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IAU_CMD_END_ADDR = AIC_D_IAU_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_IAU_PRG_ST_ADDR  = AIC_D_IAU_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_IAU_PRG_END_ADDR = AIC_D_IAU_PRG_END_ADDR;
    // D_DPU
  parameter loc_addr_t AIC_LOC_D_DPU_CSR_ST_ADDR  = AIC_D_DPU_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_DPU_CSR_END_ADDR = AIC_D_DPU_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_DPU_CMD_ST_ADDR  = AIC_D_DPU_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_DPU_CMD_END_ADDR = AIC_D_DPU_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_D_DPU_PRG_ST_ADDR  = AIC_D_DPU_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_D_DPU_PRG_END_ADDR = AIC_D_DPU_PRG_END_ADDR;

    // HP_DMA common parts
  parameter loc_addr_t AIC_LOC_HP_DMA_MMU_CSR_ST_ADDR  = AIC_HP_DMA_MMU_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_MMU_CSR_END_ADDR = AIC_HP_DMA_MMU_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_COMMON_CSR_ST_ADDR  = AIC_HP_DMA_COMMON_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_COMMON_CSR_END_ADDR = AIC_HP_DMA_COMMON_CSR_END_ADDR;
    // HP_DMA_0
  parameter loc_addr_t AIC_LOC_HP_DMA_0_CSR_ST_ADDR  = AIC_HP_DMA_0_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_0_CSR_END_ADDR = AIC_HP_DMA_0_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_0_CMD_ST_ADDR  = AIC_HP_DMA_0_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_0_CMD_END_ADDR = AIC_HP_DMA_0_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_0_PRG_ST_ADDR  = AIC_HP_DMA_0_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_0_PRG_END_ADDR = AIC_HP_DMA_0_PRG_END_ADDR;
    // HP_DMA_1
  parameter loc_addr_t AIC_LOC_HP_DMA_1_CSR_ST_ADDR  = AIC_HP_DMA_1_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_1_CSR_END_ADDR = AIC_HP_DMA_1_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_1_CMD_ST_ADDR  = AIC_HP_DMA_1_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_1_CMD_END_ADDR = AIC_HP_DMA_1_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_1_PRG_ST_ADDR  = AIC_HP_DMA_1_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_1_PRG_END_ADDR = AIC_HP_DMA_1_PRG_END_ADDR;

  ///////////////////////////
    // IP's
  parameter ext_addr_t AIC_DMC_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_DMC_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_LS_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_DMC_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_DMC_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_LS_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_DMC_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_LS_M_IFD_0_ST_ADDR;
  parameter ext_addr_t AIC_DMC_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_LS_RESERVED_END_ADDR;

  parameter ext_addr_t AIC_MID_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_MID_M_MVMEXE_ST_ADDR;
  parameter ext_addr_t AIC_MID_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_MID_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_MID_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_MID_M_MVMEXE_ST_ADDR;
  parameter ext_addr_t AIC_MID_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_MID_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_MID_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_MID_M_MVMEXE_ST_ADDR;
  parameter ext_addr_t AIC_MID_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_MID_RESERVED_END_ADDR;

  parameter ext_addr_t AIC_DID_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_DID_D_DWPU_ST_ADDR;
  parameter ext_addr_t AIC_DID_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_DID_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_DID_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_DID_D_DWPU_ST_ADDR;
  parameter ext_addr_t AIC_DID_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_DID_RESERVED_END_ADDR;
  parameter ext_addr_t AIC_DID_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_DID_D_DWPU_ST_ADDR;
  parameter ext_addr_t AIC_DID_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_DID_RESERVED_END_ADDR;
    // HP_DMA
  parameter ext_addr_t AIC_HP_DMA_CSR_ST_ADDR  = AICORE_0_DATAPATH_CSR_DMA_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_CSR_END_ADDR = AICORE_0_DATAPATH_CSR_DMA_END_ADDR;
  parameter ext_addr_t AIC_HP_DMA_CMD_ST_ADDR  = AICORE_0_DATAPATH_COMMAND_DMA_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_CMD_END_ADDR = AICORE_0_DATAPATH_COMMAND_DMA_END_ADDR;
  parameter ext_addr_t AIC_HP_DMA_PRG_ST_ADDR  = AICORE_0_DATAPATH_INSTRUCTIONS_DMA_ST_ADDR;
  parameter ext_addr_t AIC_HP_DMA_PRG_END_ADDR = AICORE_0_DATAPATH_INSTRUCTIONS_DMA_END_ADDR;

    // local address IP's
  parameter loc_addr_t AIC_LOC_DMC_CSR_ST_ADDR  = AIC_DMC_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_DMC_CSR_END_ADDR = AIC_DMC_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_DMC_CMD_ST_ADDR  = AIC_DMC_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_DMC_CMD_END_ADDR = AIC_DMC_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_DMC_PRG_ST_ADDR  = AIC_DMC_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_DMC_PRG_END_ADDR = AIC_DMC_PRG_END_ADDR;

  parameter loc_addr_t AIC_LOC_MID_CSR_ST_ADDR  = AIC_MID_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_MID_CSR_END_ADDR = AIC_MID_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_MID_CMD_ST_ADDR  = AIC_MID_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_MID_CMD_END_ADDR = AIC_MID_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_MID_PRG_ST_ADDR  = AIC_MID_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_MID_PRG_END_ADDR = AIC_MID_PRG_END_ADDR;

  parameter loc_addr_t AIC_LOC_DID_CSR_ST_ADDR  = AIC_DID_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_DID_CSR_END_ADDR = AIC_DID_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_DID_CMD_ST_ADDR  = AIC_DID_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_DID_CMD_END_ADDR = AIC_DID_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_DID_PRG_ST_ADDR  = AIC_DID_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_DID_PRG_END_ADDR = AIC_DID_PRG_END_ADDR;
    // HP_DMA
  parameter loc_addr_t AIC_LOC_HP_DMA_CSR_ST_ADDR  = AIC_HP_DMA_CSR_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_CSR_END_ADDR = AIC_HP_DMA_CSR_END_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_CMD_ST_ADDR  = AIC_HP_DMA_CMD_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_CMD_END_ADDR = AIC_HP_DMA_CMD_END_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_PRG_ST_ADDR  = AIC_HP_DMA_PRG_ST_ADDR;
  parameter loc_addr_t AIC_LOC_HP_DMA_PRG_END_ADDR = AIC_HP_DMA_PRG_END_ADDR;

  //////////////////////////////
  ///// Regions
  typedef longint aic_region_t[3];
    //////////////////// IPs:
    // DMC:
  parameter longint AIC_LOC_DMC_REGION_ST_ADDR[3] = {
    AIC_LOC_DMC_CSR_ST_ADDR, AIC_LOC_DMC_CMD_ST_ADDR, AIC_LOC_DMC_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_MID_REGION_ST_ADDR[4] = {
    AIC_LOC_MID_CSR_ST_ADDR, AIC_LOC_MID_CMD_ST_ADDR, AIC_LOC_MID_PRG_ST_ADDR, AIC_LOC_CFG_CSR_MID_PART_ST_ADDR
  };
  parameter longint AIC_LOC_DID_REGION_ST_ADDR[3] = {
    AIC_LOC_DID_CSR_ST_ADDR, AIC_LOC_DID_CMD_ST_ADDR, AIC_LOC_DID_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_DMC_REGION_END_ADDR[3] = {
    AIC_LOC_DMC_CSR_END_ADDR, AIC_LOC_DMC_CMD_END_ADDR, AIC_LOC_DMC_PRG_END_ADDR
  };
  parameter longint AIC_LOC_MID_REGION_END_ADDR[4] = {
    AIC_LOC_MID_CSR_END_ADDR, AIC_LOC_MID_CMD_END_ADDR, AIC_LOC_MID_PRG_END_ADDR, AIC_LOC_CFG_CSR_MID_PART_END_ADDR
  };
  parameter longint AIC_LOC_DID_REGION_END_ADDR[3] = {
    AIC_LOC_DID_CSR_END_ADDR, AIC_LOC_DID_CMD_END_ADDR, AIC_LOC_DID_PRG_END_ADDR
  };

    // DMC devs:
  parameter longint AIC_LOC_M_IFD_0_REGION_ST_ADDR[3] = {
    AIC_LOC_M_IFD_0_CSR_ST_ADDR, AIC_LOC_M_IFD_0_CMD_ST_ADDR, AIC_LOC_M_IFD_0_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_M_IFD_1_REGION_ST_ADDR[3] = {
    AIC_LOC_M_IFD_1_CSR_ST_ADDR, AIC_LOC_M_IFD_1_CMD_ST_ADDR, AIC_LOC_M_IFD_1_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_M_IFD_2_REGION_ST_ADDR[3] = {
    AIC_LOC_M_IFD_2_CSR_ST_ADDR, AIC_LOC_M_IFD_2_CMD_ST_ADDR, AIC_LOC_M_IFD_2_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_M_IFD_W_REGION_ST_ADDR[3] = {
    AIC_LOC_M_IFD_W_CSR_ST_ADDR, AIC_LOC_M_IFD_W_CMD_ST_ADDR, AIC_LOC_M_IFD_W_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_M_ODR_REGION_ST_ADDR[3] = {
    AIC_LOC_M_ODR_CSR_ST_ADDR, AIC_LOC_M_ODR_CMD_ST_ADDR, AIC_LOC_M_ODR_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_D_IFD_0_REGION_ST_ADDR[3] = {
    AIC_LOC_D_IFD_0_CSR_ST_ADDR, AIC_LOC_D_IFD_0_CMD_ST_ADDR, AIC_LOC_D_IFD_0_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_D_IFD_1_REGION_ST_ADDR[3] = {
    AIC_LOC_D_IFD_1_CSR_ST_ADDR, AIC_LOC_D_IFD_1_CMD_ST_ADDR, AIC_LOC_D_IFD_1_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_D_ODR_REGION_ST_ADDR[3] = {
    AIC_LOC_D_ODR_CSR_ST_ADDR, AIC_LOC_D_ODR_CMD_ST_ADDR, AIC_LOC_D_ODR_PRG_ST_ADDR
  };

  parameter longint AIC_LOC_M_IFD_0_REGION_END_ADDR[3] = {
    AIC_LOC_M_IFD_0_CSR_END_ADDR, AIC_LOC_M_IFD_0_CMD_END_ADDR, AIC_LOC_M_IFD_0_PRG_END_ADDR
  };
  parameter longint AIC_LOC_M_IFD_1_REGION_END_ADDR[3] = {
    AIC_LOC_M_IFD_1_CSR_END_ADDR, AIC_LOC_M_IFD_1_CMD_END_ADDR, AIC_LOC_M_IFD_1_PRG_END_ADDR
  };
  parameter longint AIC_LOC_M_IFD_2_REGION_END_ADDR[3] = {
    AIC_LOC_M_IFD_2_CSR_END_ADDR, AIC_LOC_M_IFD_2_CMD_END_ADDR, AIC_LOC_M_IFD_2_PRG_END_ADDR
  };
  parameter longint AIC_LOC_M_IFD_W_REGION_END_ADDR[3] = {
    AIC_LOC_M_IFD_W_CSR_END_ADDR, AIC_LOC_M_IFD_W_CMD_END_ADDR, AIC_LOC_M_IFD_W_PRG_END_ADDR
  };
  parameter longint AIC_LOC_M_ODR_REGION_END_ADDR[3] = {
    AIC_LOC_M_ODR_CSR_END_ADDR, AIC_LOC_M_ODR_CMD_END_ADDR, AIC_LOC_M_ODR_PRG_END_ADDR
  };
  parameter longint AIC_LOC_D_IFD_0_REGION_END_ADDR[3] = {
    AIC_LOC_D_IFD_0_CSR_END_ADDR, AIC_LOC_D_IFD_0_CMD_END_ADDR, AIC_LOC_D_IFD_0_PRG_END_ADDR
  };
  parameter longint AIC_LOC_D_IFD_1_REGION_END_ADDR[3] = {
    AIC_LOC_D_IFD_1_CSR_END_ADDR, AIC_LOC_D_IFD_1_CMD_END_ADDR, AIC_LOC_D_IFD_1_PRG_END_ADDR
  };
  parameter longint AIC_LOC_D_ODR_REGION_END_ADDR[3] = {
    AIC_LOC_D_ODR_CSR_END_ADDR, AIC_LOC_D_ODR_CMD_END_ADDR, AIC_LOC_D_ODR_PRG_END_ADDR
  };

    // MID devs:
  parameter longint AIC_LOC_M_MVM_REGION_ST_ADDR[6] = {
    AIC_LOC_M_MVM_EXE_CSR_ST_ADDR, AIC_LOC_M_MVM_EXE_CMD_ST_ADDR, AIC_LOC_M_MVM_EXE_PRG_ST_ADDR,
    AIC_LOC_M_MVM_PRG_CSR_ST_ADDR, AIC_LOC_M_MVM_PRG_CMD_ST_ADDR, AIC_LOC_M_MVM_PRG_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_M_IAU_REGION_ST_ADDR[3] = {
    AIC_LOC_M_IAU_CSR_ST_ADDR, AIC_LOC_M_IAU_CMD_ST_ADDR, AIC_LOC_M_IAU_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_M_DPU_REGION_ST_ADDR[3] = {
    AIC_LOC_M_DPU_CSR_ST_ADDR, AIC_LOC_M_DPU_CMD_ST_ADDR, AIC_LOC_M_DPU_PRG_ST_ADDR
  };

  parameter longint AIC_LOC_M_MVM_REGION_END_ADDR[6] = {
    AIC_LOC_M_MVM_EXE_CSR_END_ADDR, AIC_LOC_M_MVM_EXE_CMD_END_ADDR, AIC_LOC_M_MVM_EXE_PRG_END_ADDR,
    AIC_LOC_M_MVM_PRG_CSR_END_ADDR, AIC_LOC_M_MVM_PRG_CMD_END_ADDR, AIC_LOC_M_MVM_PRG_PRG_END_ADDR
  };
  parameter longint AIC_LOC_M_IAU_REGION_END_ADDR[3] = {
    AIC_LOC_M_IAU_CSR_END_ADDR, AIC_LOC_M_IAU_CMD_END_ADDR, AIC_LOC_M_IAU_PRG_END_ADDR
  };
  parameter longint AIC_LOC_M_DPU_REGION_END_ADDR[3] = {
    AIC_LOC_M_DPU_CSR_END_ADDR, AIC_LOC_M_DPU_CMD_END_ADDR, AIC_LOC_M_DPU_PRG_END_ADDR
  };

    // DID devs:
  parameter longint AIC_LOC_D_DWPU_REGION_ST_ADDR[3] = {
    AIC_LOC_D_DWPU_CSR_ST_ADDR, AIC_LOC_D_DWPU_CMD_ST_ADDR, AIC_LOC_D_DWPU_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_D_IAU_REGION_ST_ADDR[3] = {
    AIC_LOC_D_IAU_CSR_ST_ADDR, AIC_LOC_D_IAU_CMD_ST_ADDR, AIC_LOC_D_IAU_PRG_ST_ADDR
  };
  parameter longint AIC_LOC_D_DPU_REGION_ST_ADDR[3] = {
    AIC_LOC_D_DPU_CSR_ST_ADDR, AIC_LOC_D_DPU_CMD_ST_ADDR, AIC_LOC_D_DPU_PRG_ST_ADDR
  };

  parameter longint AIC_LOC_D_DWPU_REGION_END_ADDR[3] = {
    AIC_LOC_D_DWPU_CSR_END_ADDR, AIC_LOC_D_DWPU_CMD_END_ADDR, AIC_LOC_D_DWPU_PRG_END_ADDR
  };
  parameter longint AIC_LOC_D_IAU_REGION_END_ADDR[3] = {
    AIC_LOC_D_IAU_CSR_END_ADDR, AIC_LOC_D_IAU_CMD_END_ADDR, AIC_LOC_D_IAU_PRG_END_ADDR
  };
  parameter longint AIC_LOC_D_DPU_REGION_END_ADDR[3] = {
    AIC_LOC_D_DPU_CSR_END_ADDR, AIC_LOC_D_DPU_CMD_END_ADDR, AIC_LOC_D_DPU_PRG_END_ADDR
  };
endpackage
`endif // AIC_ADDR_MAP_PKG_SV
