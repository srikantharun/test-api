// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024



// maximum number of BITS passed within vector fields
`ifndef TREK_MAX_IO_VECTOR_VALUE_SIZE
 `define TREK_MAX_IO_VECTOR_VALUE_SIZE 1024
`endif // TREK_MAX_IO_VECTOR_VALUE_SIZE

///@defgroup dpi_g DPI Functions
///
/// These methods define the SV Application Programming Interface to TrekSoC. They are used
/// to pull data in and out of TrekSoC at runtime, to a Verilog simulator or emulator, etc.
///
/// The methods can be loosely arranged into four groups...
///
///@{

///@defgroup dpi_1_se_g  DPI: Starting and Ending TrekSoc
///
/// Starting and Ending TrekSoC
/// ---------------------------
///
/// TrekSoC always thinks it is *in charge* of a test. Once TrekSoC believes that all *events* have
/// been observed, the value returned by `trek_done()` will change from `false` to `true`.
///
/// All method calls are non-blocking.
///
///@{

///@brief Check to see if the test has finished
///@return 1 if the test has completed, 0 otherwise.
import "DPI-C" context function int               trek_done                      ( );

///@} // end of dpi_1_se_g

///@defgroup dpi_2_c2t_g  DPI: C2T Messages
///
/// C2T interface
/// -------------
/// When the PSS/graph model (aka. "C") wants to send messages to the testbench (aka. "T"), it uses methods in this category.
/// All method calls are non-blocking.
///
///@{

///@brief Issue a message from the PSS/Graph model to the testbench using UVM messaging.
///@param[in] timestamp  TBD
///@param[in] cpu_id     TBD
///@param[in] message    TBD
///@return               TBD
///@todo
import "DPI-C" context function int       trek_c2t_message               ( input longint unsigned timestamp, input int cpu_id, input longint unsigned message );

///@} // end of dpi_2_c2t_g

///@defgroup dpi_3_get_g  DPI: TLM "Get" Interface
///
/// TLM "Get" interface
/// -------------------
///
/// Methods in this category allow a testbench to *pull* TLM transactions from the PSS/Graph model into the
/// testbench. All method calls are non-blocking.
///
/// Each thread through the graph that interacts with the testbench maintains at least one *port*, identified
/// by a unique `tb_path` identifier/name. Ports used with the *Get* interface will be of type `hsi::get_port`
/// or `hsi::master_port`.
///
/// The general flow for the testbench side is for each thread to poll `trek_can_get()` until it returns `true`.
/// Then it will call the various `trek_get_...()`  methods to retrieve the values of each field. Note that you
/// can retrieve only the fields that you need. When you are *done* retrieving fields, you call `trek_get_done()`.
/// On a `pss::get_port`, this indicates that you are *done* with the transaction and on a `pss::master_port` it
/// indicates that you are ready for another transaction. (A `pss::master_port` indicates *done* by sending a
/// response back through its *put* interface.
///
/// Note that the numeric fields are all stored as 64-bit integers or 64-bit unsigned integers. The return
/// value is checked for the app
///
///@{

///@brief Is a transaction available on this port?
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_can_get                   ( input string tb_path );

///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects an integer field within the available transaction.
///@return  8-bit signed field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function byte              trek_get_byte                  ( input string tb_path, input string field_name );
///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects an integer field within the available transaction.
///@return  16-bit signed field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function shortint          trek_get_shortint              ( input string tb_path, input string field_name );
///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects an integer field within the available transaction.
///@return  32-bit signed field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function int               trek_get_int                   ( input string tb_path, input string field_name );
///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects an integer field within the available transaction.
///@return  64-bit signed field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function longint           trek_get_longint               ( input string tb_path, input string field_name );

///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects an integer field within the available transaction.
///@return  8-bit unsigned field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function byte unsigned     trek_get_byte_unsigned         ( input string tb_path, input string field_name );
///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects an integer field within the available transaction.
///@return  16-bit unsigned field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function shortint unsigned trek_get_shortint_unsigned     ( input string tb_path, input string field_name );
///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects an integer field within the available transaction.
///@return  32-bit unsigned field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function int unsigned      trek_get_int_unsigned          ( input string tb_path, input string field_name );
///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects an integer field within the available transaction.
///@return  64-bit unsigned field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function longint unsigned  trek_get_longint_unsigned      ( input string tb_path, input string field_name );

///@brief From the transaction available on this port, return the contents of the given field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects a `pss::bit` field within the available transaction.
///@return  String field value. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function string            trek_get_string                ( input string tb_path, input string field_name );

///@brief From the transaction available on this port, return the number of bytes in the given bitvector field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects a pss::bytes field within the available transaction.
///@return  32-bit unsigned number of bytes. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function int unsigned      trek_get_bitvector_size        ( input string tb_path, input string field_name );
///@brief From the transaction available on this port, return the contents of the given bitvector field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects a pss::bytes field within the available transaction.
///@param[out] value  Two-state bitvector value in the field. Typically, only the low-order bytes of the vector are valid. Maximum width is from the Verilog macro `TREK_MAX_IO_VECTOR_VALUE_SIZE`.
///@return  `true` if the contents of `value` are valid, `false` if the value is not valid
import "DPI-C" context function int               trek_get_bitvector             ( input string tb_path, input string field_name, output bit[`TREK_MAX_IO_VECTOR_VALUE_SIZE-1:0] value );

///@brief From the transaction available on this port, return the number of bytes in the given byte array field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects a pss::bytes field within the available transaction.
///@return  32-bit unsigned number of bytes. If trek_can_get() is `false` the returned value is undefined.
import "DPI-C" context function int unsigned      trek_get_bytearray_size        ( input string tb_path, input string field_name );
///@brief From the transaction available on this port, return the contents of the given byte array field.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that selects a pss::bytes field within the available transaction.
///@param[out] value  Two-state bitvector value in the field. Typically, only the low-order bytes of the vector are valid. Maximum width is from the Verilog macro `TREK_MAX_IO_VECTOR_VALUE_SIZE`.
///@return  `true` if the contents of `value` are valid, `false` if the value is not valid
import "DPI-C" context function int               trek_get_bytearray             ( input string tb_path, input string field_name, output byte unsigned value[] );

///@brief  From the transaction available on this port, return the value of the transaction_id.
///        Note that UINT64_MAX (-1) is the "default"/"sentinal" for an unset value and generally means we must operate in-order.
///        Note also that we will return zero on failure, so we suggest that you do not use that value in your modeling.
///@note   Trek uses 64-bit transaction_ids, while UVM uses 32-bit transaction_ids
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and the test bench.
///@return  zero on failure, otherwise the transaction_id
import "DPI-C" context function longint unsigned  trek_get_transaction_id        ( input string tb_path );


///@brief The testbench uses this method to indicate to the PSS/Graph model that no more fields will be retrieved from the current transaction. TrekSoC will *pop* it from the outgoing port.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@return  `true` if the transaction was *popped* successfully, `false` otherwise
import "DPI-C" context function int               trek_get_done                  ( input string tb_path );

///@} // end of dpi_3_get_g

///@defgroup dpi_4_put_g  DPI: TLM "Put" Interface
///
/// TLM "Put" interface
/// -------------------
///
/// Methods in this category allow a testbench to *push* TLM transactions to the PSS/Graph model from the
/// testbench. All method calls are non-blocking.
///
/// Each thread through the graph that interacts with the testbench maintains at least one *port*, identified
/// by a unique `tb_path` identifier/name. Ports used with the *Put* interface will be of type `hsi::put_port`,
/// `hsi::master_port` or `hsi::check_port`.
///
/// The general flow for the testbench side is for each thread to poll `trek_can_get()` until it returns `true`.
/// The first call to a `trek_put_...()` method will create an empty transaction in the port. Subsequent calls
/// to each of the various `trek_put_...()` will create fields in that transaction and set their values. When
/// you are *done* sending fields, you call `trek_put_done()`, to finalize creation of the transaction and
/// *push* the transaction into the port.
///
/// Note that the numeric fields are all stored as 64-bit integers or 64-bit unsigned integers. The *value*
/// argument is checked for the appropriate range/size when you call the `trek_put_...()` method.
/// 
///@{

///@brief Is there space to push a TLM transaction on this port?
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_can_put                   ( input string tb_path );

///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names an integer field within the available transaction.
///@param[in] value  8-bit signed number to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_byte                  ( input string tb_path, input string field_name, input byte              value );
///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names an integer field within the available transaction.
///@param[in] value  16-bit signed number to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_shortint              ( input string tb_path, input string field_name, input shortint          value );
///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names an integer field within the available transaction.
///@param[in] value  32-bit signed number to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_int                   ( input string tb_path, input string field_name, input int               value );
///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names an integer field within the available transaction.
///@param[in] value  64-bit signed number to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_longint               ( input string tb_path, input string field_name, input longint           value );

///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names a `pss::bit` field within the available transaction.
///@param[in] value  8-bit unsigned number to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_byte_unsigned         ( input string tb_path, input string field_name, input byte unsigned     value );
///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names a `pss::bit` field within the available transaction.
///@param[in] value  16-bit unsigned number to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_shortint_unsigned     ( input string tb_path, input string field_name, input shortint unsigned value );
///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names a `pss::bit` field within the available transaction.
///@param[in] value  32-bit unsigned number to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_int_unsigned          ( input string tb_path, input string field_name, input int unsigned      value );
///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names a `pss::bit` field within the available transaction.
///@param[in] value 64-bit unsigned number to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_longint_unsigned      ( input string tb_path, input string field_name, input longint unsigned  value );

///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names a `std::string` field within the available transaction.
///@param[in] value  string value to store in the field contents.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_string                ( input string tb_path, input string field_name, input string            value );

///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names a `pss::bytes` field within the available transaction.
///@param[in] size_in_bytes  Number of bytes that are valid in the vector. If you need to send a bitvector that does not fit evenly into bytes (for example, 125 bits), then you should use another field to capture the "extra" bits.
///@param[in] value  Two-state bitvector. Typically, only the low-order bytes of the vector are valid. Maximum width is from the Verilog macro `TREK_MAX_IO_VECTOR_VALUE_SIZE`.
///@return  `true` if the contents of `value` are valid, `false` if the value is not valid
import "DPI-C" context function int               trek_put_bitvector             ( input string tb_path, input string field_name, input int unsigned size_in_bytes, input bit[`TREK_MAX_IO_VECTOR_VALUE_SIZE-1:0] value );

///@brief Create or replace a field in the incoming transaction.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@param[in] field_name  String that names a `pss::bytes` field within the available transaction.
///@param[in] value  Array of two-state bytes.
///@return  `true` if the contents of `value` are valid, `false` if the value is not valid
import "DPI-C" context function int               trek_put_bytearray             ( input string tb_path, input string field_name, input byte unsigned value[] );

///@brief  Store the transaction_id for the incoming transaction. This is
///        important for tracking out-of-order request completion.
///@note   Trek uses 64-bit transaction_ids, while UVM uses 32-bit transaction_ids
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph
///                    model and the test bench.
///@param[in] transaction_id  Value to store as the ID.
///@return  zero on success, non-zero error code otherwise.
import "DPI-C" context function int               trek_put_transaction_id        ( input string tb_path, input longint unsigned transaction_id = 64'hffffffff_ffffffff);


///@brief The testbench uses this method to indicate to the PSS/Graph model that no more fields will be added to the current transaction. TrekSoC will *push* the transaction into the incoming port.
///@param[in] tb_path  Unique port identifier/name; identical in the PSS/Graph model and in the testbench.
///@return  `true` if the transaction was *popped* successfully, `false` otherwise
import "DPI-C" context function int               trek_put_done                  ( input string tb_path );

///@} // end of  dpi_4_put_g

///@} // end of dpi_g
