// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024



`ifndef GUARD__TREK_DELAY_REQ_DELAY_REQ_ADAPTER__SV
`define GUARD__TREK_DELAY_REQ_DELAY_REQ_ADAPTER__SV

virtual class trek_delay_req_delay_req_adapter#(
    type VIP_REQ = `TREK_TLM_ADAPTER_VIP_BASE_TYPE,
    type VIP_RSP = VIP_REQ)
        extends trek_tlm_adapter#(
            .TREK_REQ(trek_delay_req),
            .TREK_RSP(trek_delay_req),
            .VIP_REQ(VIP_REQ),
            .VIP_RSP(VIP_RSP));

  function new(string name = "trek_delay_req_delay_req_adapter");
    super.new(name);
  endfunction
endclass: trek_delay_req_delay_req_adapter

`endif  // GUARD__TREK_DELAY_REQ_DELAY_REQ_ADAPTER__SV
