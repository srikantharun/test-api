//
// Copyright (c) 2005-2024 Imperas Software Ltd. All Rights Reserved.
//
// THIS SOFTWARE CONTAINS CONFIDENTIAL INFORMATION AND TRADE SECRETS
// OF IMPERAS SOFTWARE LTD. USE, DISCLOSURE, OR REPRODUCTION IS PROHIBITED
// EXCEPT AS MAY BE PROVIDED FOR IN A WRITTEN AGREEMENT WITH IMPERAS SOFTWARE LTD.
//
//

package RISCV_coverage_pkg_cva6v;

import idvPkg::*;
import rvviApiPkg::*;

import idvApiPkg::*;

//`include "coverage/RISCV_coverage_global.svh"
`include "RISCV_coverage_common_cva6v.svh"
`include "coverage/RISCV_trace_data.svh"
`include "coverage/RISCV_config_checks.svh"
`include "RISCV_instruction_base_cva6v.svh"

`include "RISCV_coverage_base_cva6v.svh"

endpackage

