// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: Leonidas Katselas <leonidas.katselas@axelera.ai>

/// Dual core AVC HEVC JPEG DECODER with RISC-V IP
///
module codec
  import allegro_codec_pkg::*;
(
  /// Clock, positive edge triggered
  input  wire i_clk,
  input  wire i_mclk,
  /// Asynchronous reset, active low
  input  wire i_rst_n,
  input  wire i_mrst_n,
  /// AXI master 0 write address signals
  output logic [        CODEC_AXI_ID_WIDTH-1:0] o_dec_0_axi_m_awid,
  output logic [      CODEC_AXI_ADDR_WIDTH-1:0] o_dec_0_axi_m_awaddr,
  output logic [       CODEC_AXI_LEN_WIDTH-1:0] o_dec_0_axi_m_awlen,
  output logic [      CODEC_AXI_SIZE_WIDTH-1:0] o_dec_0_axi_m_awsize,
  output logic [      CODEC_AXI_PROT_WIDTH-1:0] o_dec_0_axi_m_awprot,
  output logic [CODEC_AXI_BURST_TYPE_WIDTH-1:0] o_dec_0_axi_m_awburst,
  output logic                                  o_dec_0_axi_m_awvalid,
  input  logic                                  i_dec_0_axi_m_awready,
  /// AXI master 0 write data signals
  output logic [      CODEC_AXI_DATA_WIDTH-1:0] o_dec_0_axi_m_wdata,
  output logic [     CODEC_AXI_WSTRB_WIDTH-1:0] o_dec_0_axi_m_wstrb,
  output logic                                  o_dec_0_axi_m_wlast,
  output logic                                  o_dec_0_axi_m_wvalid,
  input  logic                                  i_dec_0_axi_m_wready,
  /// AXI master 0 write response signals
  input  logic [      CODEC_AXI_RESP_WIDTH-1:0] i_dec_0_axi_m_bresp,
  input  logic [        CODEC_AXI_ID_WIDTH-1:0] i_dec_0_axi_m_bid,
  input  logic                                  i_dec_0_axi_m_bvalid,
  output logic                                  o_dec_0_axi_m_bready,
  /// AXI master 0 read address signals
  output logic [        CODEC_AXI_ID_WIDTH-1:0] o_dec_0_axi_m_arid,
  output logic [      CODEC_AXI_ADDR_WIDTH-1:0] o_dec_0_axi_m_araddr,
  output logic [       CODEC_AXI_LEN_WIDTH-1:0] o_dec_0_axi_m_arlen,
  output logic [      CODEC_AXI_SIZE_WIDTH-1:0] o_dec_0_axi_m_arsize,
  output logic [      CODEC_AXI_PROT_WIDTH-1:0] o_dec_0_axi_m_arprot,
  output logic [CODEC_AXI_BURST_TYPE_WIDTH-1:0] o_dec_0_axi_m_arburst,
  output logic                                  o_dec_0_axi_m_arvalid,
  input  logic                                  i_dec_0_axi_m_arready,
  /// AXI master 0 read data signals
  input  logic [        CODEC_AXI_ID_WIDTH-1:0] i_dec_0_axi_m_rid,
  input  logic [      CODEC_AXI_DATA_WIDTH-1:0] i_dec_0_axi_m_rdata,
  input  logic                                  i_dec_0_axi_m_rlast,
  input  logic [      CODEC_AXI_RESP_WIDTH-1:0] i_dec_0_axi_m_rresp,
  input  logic                                  i_dec_0_axi_m_rvalid,
  output logic                                  o_dec_0_axi_m_rready,
  /// AXI master 1 write address signals
  output logic [        CODEC_AXI_ID_WIDTH-1:0] o_dec_1_axi_m_awid,
  output logic [      CODEC_AXI_ADDR_WIDTH-1:0] o_dec_1_axi_m_awaddr,
  output logic [       CODEC_AXI_LEN_WIDTH-1:0] o_dec_1_axi_m_awlen,
  output logic [      CODEC_AXI_SIZE_WIDTH-1:0] o_dec_1_axi_m_awsize,
  output logic [      CODEC_AXI_PROT_WIDTH-1:0] o_dec_1_axi_m_awprot,
  output logic [CODEC_AXI_BURST_TYPE_WIDTH-1:0] o_dec_1_axi_m_awburst,
  output logic                                  o_dec_1_axi_m_awvalid,
  input  logic                                  i_dec_1_axi_m_awready,
  /// AXI master 1 write data signals
  output logic [      CODEC_AXI_DATA_WIDTH-1:0] o_dec_1_axi_m_wdata,
  output logic [     CODEC_AXI_WSTRB_WIDTH-1:0] o_dec_1_axi_m_wstrb,
  output logic                                  o_dec_1_axi_m_wlast,
  output logic                                  o_dec_1_axi_m_wvalid,
  input  logic                                  i_dec_1_axi_m_wready,
  /// AXI master 1 write response signals
  input  logic [      CODEC_AXI_RESP_WIDTH-1:0] i_dec_1_axi_m_bresp,
  input  logic [        CODEC_AXI_ID_WIDTH-1:0] i_dec_1_axi_m_bid,
  input  logic                                  i_dec_1_axi_m_bvalid,
  output logic                                  o_dec_1_axi_m_bready,
  /// AXI master 1 read address signals
  output logic [        CODEC_AXI_ID_WIDTH-1:0] o_dec_1_axi_m_arid,
  output logic [      CODEC_AXI_ADDR_WIDTH-1:0] o_dec_1_axi_m_araddr,
  output logic [       CODEC_AXI_LEN_WIDTH-1:0] o_dec_1_axi_m_arlen,
  output logic [      CODEC_AXI_SIZE_WIDTH-1:0] o_dec_1_axi_m_arsize,
  output logic [      CODEC_AXI_PROT_WIDTH-1:0] o_dec_1_axi_m_arprot,
  output logic [CODEC_AXI_BURST_TYPE_WIDTH-1:0] o_dec_1_axi_m_arburst,
  output logic                                  o_dec_1_axi_m_arvalid,
  input  logic                                  i_dec_1_axi_m_arready,
  /// AXI master 1 read data signals
  input  logic [        CODEC_AXI_ID_WIDTH-1:0] i_dec_1_axi_m_rid,
  input  logic [      CODEC_AXI_DATA_WIDTH-1:0] i_dec_1_axi_m_rdata,
  input  logic                                  i_dec_1_axi_m_rlast,
  input  logic                                  i_dec_1_axi_m_rvalid,
  input  logic [      CODEC_AXI_RESP_WIDTH-1:0] i_dec_1_axi_m_rresp,
  output logic                                  o_dec_1_axi_m_rready,
  /// AXI master 2 write address signals
  output logic [        CODEC_AXI_ID_WIDTH-1:0] o_dec_2_axi_m_awid,
  output logic [      CODEC_AXI_ADDR_WIDTH-1:0] o_dec_2_axi_m_awaddr,
  output logic [       CODEC_AXI_LEN_WIDTH-1:0] o_dec_2_axi_m_awlen,
  output logic [      CODEC_AXI_SIZE_WIDTH-1:0] o_dec_2_axi_m_awsize,
  output logic [      CODEC_AXI_PROT_WIDTH-1:0] o_dec_2_axi_m_awprot,
  output logic [CODEC_AXI_BURST_TYPE_WIDTH-1:0] o_dec_2_axi_m_awburst,
  output logic                                  o_dec_2_axi_m_awvalid,
  input  logic                                  i_dec_2_axi_m_awready,
  /// AXI master 2 write data signals
  output logic [      CODEC_AXI_DATA_WIDTH-1:0] o_dec_2_axi_m_wdata,
  output logic [     CODEC_AXI_WSTRB_WIDTH-1:0] o_dec_2_axi_m_wstrb,
  output logic                                  o_dec_2_axi_m_wlast,
  output logic                                  o_dec_2_axi_m_wvalid,
  input  logic                                  i_dec_2_axi_m_wready,
  /// AXI master 2 write response signals
  input  logic [      CODEC_AXI_RESP_WIDTH-1:0] i_dec_2_axi_m_bresp,
  input  logic [        CODEC_AXI_ID_WIDTH-1:0] i_dec_2_axi_m_bid,
  input  logic                                  i_dec_2_axi_m_bvalid,
  output logic                                  o_dec_2_axi_m_bready,
  /// AXI master 2 read address signals
  output logic [        CODEC_AXI_ID_WIDTH-1:0] o_dec_2_axi_m_arid,
  output logic [      CODEC_AXI_ADDR_WIDTH-1:0] o_dec_2_axi_m_araddr,
  output logic [       CODEC_AXI_LEN_WIDTH-1:0] o_dec_2_axi_m_arlen,
  output logic [      CODEC_AXI_SIZE_WIDTH-1:0] o_dec_2_axi_m_arsize,
  output logic [      CODEC_AXI_PROT_WIDTH-1:0] o_dec_2_axi_m_arprot,
  output logic [CODEC_AXI_BURST_TYPE_WIDTH-1:0] o_dec_2_axi_m_arburst,
  output logic                                  o_dec_2_axi_m_arvalid,
  input  logic                                  i_dec_2_axi_m_arready,
  /// AXI master 2 read data signals
  input  logic [        CODEC_AXI_ID_WIDTH-1:0] i_dec_2_axi_m_rid,
  input  logic [      CODEC_AXI_DATA_WIDTH-1:0] i_dec_2_axi_m_rdata,
  input  logic                                  i_dec_2_axi_m_rlast,
  input  logic [      CODEC_AXI_RESP_WIDTH-1:0] i_dec_2_axi_m_rresp,
  input  logic                                  i_dec_2_axi_m_rvalid,
  output logic                                  o_dec_2_axi_m_rready,
  /// RISC-V interrupt signals
  output logic                                  o_mcu_int_next,
  input  logic                                  i_mcu_ack_next,
  input  logic                                  i_mcu_int_prev,
  output logic                                  o_mcu_ack_prev,
  /// RISC-V JTAG signals
  /// TODO:fix the naming convention
  input  wire                                   i_jtag_clk,
  input  logic                                  i_jtag_ms,
  input  logic                                  i_jtag_di,
  output logic                                  o_jtag_do,
  /// RISC-V AXI master write address signals
  output logic [        CODEC_AXI_ID_WIDTH-1:0] o_mcu_axi_m_awid,
  output logic [      CODEC_AXI_ADDR_WIDTH-1:0] o_mcu_axi_m_awaddr,
  output logic [       CODEC_AXI_LEN_WIDTH-1:0] o_mcu_axi_m_awlen,
  output logic [      CODEC_AXI_SIZE_WIDTH-1:0] o_mcu_axi_m_awsize,
  output logic [      CODEC_AXI_PROT_WIDTH-1:0] o_mcu_axi_m_awprot,
  output logic [CODEC_AXI_BURST_TYPE_WIDTH-1:0] o_mcu_axi_m_awburst,
  output logic                                  o_mcu_axi_m_awvalid,
  input  logic                                  i_mcu_axi_m_awready,
  /// RISC-V AXI master write data signals
  output logic [      CODEC_AXI_DATA_WIDTH-1:0] o_mcu_axi_m_wdata,
  output logic [     CODEC_AXI_WSTRB_WIDTH-1:0] o_mcu_axi_m_wstrb,
  output logic                                  o_mcu_axi_m_wlast,
  output logic                                  o_mcu_axi_m_wvalid,
  input  logic                                  i_mcu_axi_m_wready,
  /// RISC-V AXI master write response signals
  input  logic [      CODEC_AXI_RESP_WIDTH-1:0] i_mcu_axi_m_bresp,
  input  logic [        CODEC_AXI_ID_WIDTH-1:0] i_mcu_axi_m_bid,
  input  logic                                  i_mcu_axi_m_bvalid,
  output logic                                  o_mcu_axi_m_bready,
  /// RISC-V AXI master read address signals
  output logic [        CODEC_AXI_ID_WIDTH-1:0] o_mcu_axi_m_arid,
  output logic [      CODEC_AXI_ADDR_WIDTH-1:0] o_mcu_axi_m_araddr,
  output logic [       CODEC_AXI_LEN_WIDTH-1:0] o_mcu_axi_m_arlen,
  output logic [      CODEC_AXI_SIZE_WIDTH-1:0] o_mcu_axi_m_arsize,
  output logic [      CODEC_AXI_PROT_WIDTH-1:0] o_mcu_axi_m_arprot,
  output logic [CODEC_AXI_BURST_TYPE_WIDTH-1:0] o_mcu_axi_m_arburst,
  output logic                                  o_mcu_axi_m_arvalid,
  input  logic                                  i_mcu_axi_m_arready,
  /// RISC-V AXI master read data signals
  input  logic [        CODEC_AXI_ID_WIDTH-1:0] i_mcu_axi_m_rid,
  input  logic [      CODEC_AXI_DATA_WIDTH-1:0] i_mcu_axi_m_rdata,
  input  logic                                  i_mcu_axi_m_rlast,
  input  logic [      CODEC_AXI_RESP_WIDTH-1:0] i_mcu_axi_m_rresp,
  input  logic                                  i_mcu_axi_m_rvalid,
  output logic                                  o_mcu_axi_m_rready,
  /// APB slave signals,
  input  dcd_targ_cfg_apb_addr_t            i_cfg_apb4_s_paddr,
  input  dcd_targ_cfg_apb_data_t            i_cfg_apb4_s_pwdata,
  input  logic                                  i_cfg_apb4_s_pwrite,
  input  logic                                  i_cfg_apb4_s_psel,
  input  logic                                  i_cfg_apb4_s_penable,
  input  dcd_targ_cfg_apb_strb_t            i_cfg_apb4_s_pstrb,
  input  logic [                           2:0] i_cfg_apb4_s_pprot,
  output logic                                  o_cfg_apb4_s_pready,
  output dcd_targ_cfg_apb_data_t            o_cfg_apb4_s_prdata,
  output logic                                  o_cfg_apb4_s_pslverr,
  /// decoder global signals
  output logic                                  o_pintreq,
  output logic [                          31:0] o_pintbus,
  // DfT
  input  logic                                  i_test_mode,
  input  logic                                  i_scan_en,

  // SRAM configuration
  input  axe_tcl_sram_pkg::impl_inp_t     [3:0] i_impl,
  output axe_tcl_sram_pkg::impl_oup_t     [3:0] o_impl
);

assign o_cfg_apb4_s_pslverr = '0;

alg_vcu_dec_top u_alg_vcu_dec_top (
  .clk          (i_clk),
  .rstn         (i_rst_n),
  .awid0        (o_dec_0_axi_m_awid),
  .awaddr0      (o_dec_0_axi_m_awaddr),
  .awlen0       (o_dec_0_axi_m_awlen),
  .awsize0      (o_dec_0_axi_m_awsize),
  .awprot0      (o_dec_0_axi_m_awprot),
  .awburst0     (o_dec_0_axi_m_awburst),
  .awvalid0     (o_dec_0_axi_m_awvalid),
  .awready0     (i_dec_0_axi_m_awready),
  .wdata0       (o_dec_0_axi_m_wdata),
  .wstrb0       (o_dec_0_axi_m_wstrb),
  .wlast0       (o_dec_0_axi_m_wlast),
  .wvalid0      (o_dec_0_axi_m_wvalid),
  .wready0      (i_dec_0_axi_m_wready),
  .bready0      (o_dec_0_axi_m_bready),
  .bvalid0      (i_dec_0_axi_m_bvalid),
  .bresp0       (i_dec_0_axi_m_bresp),
  .bid0         (i_dec_0_axi_m_bid),
  .arid0        (o_dec_0_axi_m_arid),
  .araddr0      (o_dec_0_axi_m_araddr),
  .arlen0       (o_dec_0_axi_m_arlen),
  .arsize0      (o_dec_0_axi_m_arsize),
  .arprot0      (o_dec_0_axi_m_arprot),
  .arburst0     (o_dec_0_axi_m_arburst),
  .arvalid0     (o_dec_0_axi_m_arvalid),
  .arready0     (i_dec_0_axi_m_arready),
  .rid0         (i_dec_0_axi_m_rid),
  .rdata0       (i_dec_0_axi_m_rdata),
  .rlast0       (i_dec_0_axi_m_rlast),
  .rvalid0      (i_dec_0_axi_m_rvalid),
  .rresp0       (i_dec_0_axi_m_rresp),
  .rready0      (o_dec_0_axi_m_rready),
  .awid1        (o_dec_1_axi_m_awid),
  .awaddr1      (o_dec_1_axi_m_awaddr),
  .awlen1       (o_dec_1_axi_m_awlen),
  .awsize1      (o_dec_1_axi_m_awsize),
  .awprot1      (o_dec_1_axi_m_awprot),
  .awburst1     (o_dec_1_axi_m_awburst),
  .awvalid1     (o_dec_1_axi_m_awvalid),
  .awready1     (i_dec_1_axi_m_awready),
  .wdata1       (o_dec_1_axi_m_wdata),
  .wstrb1       (o_dec_1_axi_m_wstrb),
  .wlast1       (o_dec_1_axi_m_wlast),
  .wvalid1      (o_dec_1_axi_m_wvalid),
  .wready1      (i_dec_1_axi_m_wready),
  .bready1      (o_dec_1_axi_m_bready),
  .bvalid1      (i_dec_1_axi_m_bvalid),
  .bresp1       (i_dec_1_axi_m_bresp),
  .bid1         (i_dec_1_axi_m_bid),
  .arid1        (o_dec_1_axi_m_arid),
  .araddr1      (o_dec_1_axi_m_araddr),
  .arlen1       (o_dec_1_axi_m_arlen),
  .arsize1      (o_dec_1_axi_m_arsize),
  .arprot1      (o_dec_1_axi_m_arprot),
  .arburst1     (o_dec_1_axi_m_arburst),
  .arvalid1     (o_dec_1_axi_m_arvalid),
  .arready1     (i_dec_1_axi_m_arready),
  .rid1         (i_dec_1_axi_m_rid),
  .rdata1       (i_dec_1_axi_m_rdata),
  .rlast1       (i_dec_1_axi_m_rlast),
  .rvalid1      (i_dec_1_axi_m_rvalid),
  .rresp1       (i_dec_1_axi_m_rresp),
  .rready1      (o_dec_1_axi_m_rready),
  .awid2        (o_dec_2_axi_m_awid),
  .awaddr2      (o_dec_2_axi_m_awaddr),
  .awlen2       (o_dec_2_axi_m_awlen),
  .awsize2      (o_dec_2_axi_m_awsize),
  .awprot2      (o_dec_2_axi_m_awprot),
  .awburst2     (o_dec_2_axi_m_awburst),
  .awvalid2     (o_dec_2_axi_m_awvalid),
  .awready2     (i_dec_2_axi_m_awready),
  .wdata2       (o_dec_2_axi_m_wdata),
  .wstrb2       (o_dec_2_axi_m_wstrb),
  .wlast2       (o_dec_2_axi_m_wlast),
  .wvalid2      (o_dec_2_axi_m_wvalid),
  .wready2      (i_dec_2_axi_m_wready),
  .bready2      (o_dec_2_axi_m_bready),
  .bvalid2      (i_dec_2_axi_m_bvalid),
  .bresp2       (i_dec_2_axi_m_bresp),
  .bid2         (i_dec_2_axi_m_bid),
  .arid2        (o_dec_2_axi_m_arid),
  .araddr2      (o_dec_2_axi_m_araddr),
  .arlen2       (o_dec_2_axi_m_arlen),
  .arsize2      (o_dec_2_axi_m_arsize),
  .arprot2      (o_dec_2_axi_m_arprot),
  .arburst2     (o_dec_2_axi_m_arburst),
  .arvalid2     (o_dec_2_axi_m_arvalid),
  .arready2     (i_dec_2_axi_m_arready),
  .rid2         (i_dec_2_axi_m_rid),
  .rdata2       (i_dec_2_axi_m_rdata),
  .rlast2       (i_dec_2_axi_m_rlast),
  .rvalid2      (i_dec_2_axi_m_rvalid),
  .rresp2       (i_dec_2_axi_m_rresp),
  .rready2      (o_dec_2_axi_m_rready),
  .mclk         (i_mclk),
  .mrstn        (i_mrst_n),
  .mcu_int_next (o_mcu_int_next),
  .mcu_ack_next (i_mcu_ack_next),
  .mcu_int_prev (i_mcu_int_prev),
  .mcu_ack_prev (o_mcu_ack_prev),
  .jtag_clk     (i_jtag_clk),
  .jtag_ms      (i_jtag_ms),
  .jtag_di      (i_jtag_di),
  .jtag_do      (o_jtag_do),
  .awid_mcu     (o_mcu_axi_m_awid),
  .awaddr_mcu   (o_mcu_axi_m_awaddr),
  .awlen_mcu    (o_mcu_axi_m_awlen),
  .awsize_mcu   (o_mcu_axi_m_awsize),
  .awprot_mcu   (o_mcu_axi_m_awprot),
  .awburst_mcu  (o_mcu_axi_m_awburst),
  .awvalid_mcu  (o_mcu_axi_m_awvalid),
  .awready_mcu  (i_mcu_axi_m_awready),
  .wdata_mcu    (o_mcu_axi_m_wdata),
  .wstrb_mcu    (o_mcu_axi_m_wstrb),
  .wlast_mcu    (o_mcu_axi_m_wlast),
  .wvalid_mcu   (o_mcu_axi_m_wvalid),
  .wready_mcu   (i_mcu_axi_m_wready),
  .bready_mcu   (o_mcu_axi_m_bready),
  .bvalid_mcu   (i_mcu_axi_m_bvalid),
  .bresp_mcu    (i_mcu_axi_m_bresp),
  .bid_mcu      (i_mcu_axi_m_bid),
  .arid_mcu     (o_mcu_axi_m_arid),
  .araddr_mcu   (o_mcu_axi_m_araddr),
  .arlen_mcu    (o_mcu_axi_m_arlen),
  .arsize_mcu   (o_mcu_axi_m_arsize),
  .arprot_mcu   (o_mcu_axi_m_arprot),
  .arburst_mcu  (o_mcu_axi_m_arburst),
  .arvalid_mcu  (o_mcu_axi_m_arvalid),
  .arready_mcu  (i_mcu_axi_m_arready),
  .rid_mcu      (i_mcu_axi_m_rid),
  .rdata_mcu    (i_mcu_axi_m_rdata),
  .rlast_mcu    (i_mcu_axi_m_rlast),
  .rvalid_mcu   (i_mcu_axi_m_rvalid),
  .rresp_mcu    (i_mcu_axi_m_rresp),
  .rready_mcu   (o_mcu_axi_m_rready),
  .psel         (i_cfg_apb4_s_psel),
  .penable      (i_cfg_apb4_s_penable),
  .pwrite       (i_cfg_apb4_s_pwrite),
  .pwdata       (i_cfg_apb4_s_pwdata),
  .paddr        (i_cfg_apb4_s_paddr),
  .prdata       (o_cfg_apb4_s_prdata),
  .pready       (o_cfg_apb4_s_pready),
  .pintreq      (o_pintreq),
  .pintbus      (o_pintbus),
  .i_test_mode  (i_test_mode),
  .dft_clk_en   (i_scan_en),
  // Memory configutation pins
  .i_impl       (i_impl),
  .o_impl       (o_impl)
);


endmodule
