// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_h_north
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_h_north (
    input  wire                                    i_aic_4_aon_clk,
    input  wire                                    i_aic_4_aon_rst_n,
    input  wire                                    i_aic_4_clk,
    input  wire                                    i_aic_4_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_4_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_4_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_4_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_4_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_4_init_ht_axi_s_arlen,
    input  logic                                   i_aic_4_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_4_init_ht_axi_s_arprot,
    output logic                                   o_aic_4_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_4_init_ht_axi_s_arsize,
    input  logic                                   i_aic_4_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_4_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_4_init_ht_axi_s_rid,
    output logic                                   o_aic_4_init_ht_axi_s_rlast,
    input  logic                                   i_aic_4_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_4_init_ht_axi_s_rresp,
    output logic                                   o_aic_4_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_4_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_4_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_4_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_4_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_4_init_ht_axi_s_awlen,
    input  logic                                   i_aic_4_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_4_init_ht_axi_s_awprot,
    output logic                                   o_aic_4_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_4_init_ht_axi_s_awsize,
    input  logic                                   i_aic_4_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_4_init_ht_axi_s_bid,
    input  logic                                   i_aic_4_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_4_init_ht_axi_s_bresp,
    output logic                                   o_aic_4_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_4_init_ht_axi_s_wdata,
    input  logic                                   i_aic_4_init_ht_axi_s_wlast,
    output logic                                   o_aic_4_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_4_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_4_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_4_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_4_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_4_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_4_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_4_init_lt_axi_s_arlen,
    input  logic                                   i_aic_4_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_4_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_4_init_lt_axi_s_arqos,
    output logic                                   o_aic_4_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_4_init_lt_axi_s_arsize,
    input  logic                                   i_aic_4_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_4_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_4_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_4_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_4_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_4_init_lt_axi_s_awlen,
    input  logic                                   i_aic_4_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_4_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_4_init_lt_axi_s_awqos,
    output logic                                   o_aic_4_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_4_init_lt_axi_s_awsize,
    input  logic                                   i_aic_4_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_4_init_lt_axi_s_bid,
    input  logic                                   i_aic_4_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_4_init_lt_axi_s_bresp,
    output logic                                   o_aic_4_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_4_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_4_init_lt_axi_s_rid,
    output logic                                   o_aic_4_init_lt_axi_s_rlast,
    input  logic                                   i_aic_4_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_4_init_lt_axi_s_rresp,
    output logic                                   o_aic_4_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_4_init_lt_axi_s_wdata,
    input  logic                                   i_aic_4_init_lt_axi_s_wlast,
    output logic                                   o_aic_4_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_4_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_4_init_lt_axi_s_wvalid,
    output logic                                   o_aic_4_pwr_idle_val,
    output logic                                   o_aic_4_pwr_idle_ack,
    input  logic                                   i_aic_4_pwr_idle_req,
    input  wire                                    i_aic_4_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_4_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_4_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_4_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_4_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_4_targ_lt_axi_m_arlen,
    output logic                                   o_aic_4_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_4_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_4_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_4_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_4_targ_lt_axi_m_arsize,
    output logic                                   o_aic_4_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_4_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_4_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_4_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_4_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_4_targ_lt_axi_m_awlen,
    output logic                                   o_aic_4_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_4_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_4_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_4_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_4_targ_lt_axi_m_awsize,
    output logic                                   o_aic_4_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_4_targ_lt_axi_m_bid,
    output logic                                   o_aic_4_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_4_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_4_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_4_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_4_targ_lt_axi_m_rid,
    input  logic                                   i_aic_4_targ_lt_axi_m_rlast,
    output logic                                   o_aic_4_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_4_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_4_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_4_targ_lt_axi_m_wdata,
    output logic                                   o_aic_4_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_4_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_4_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_4_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_4_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_4_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_4_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_4_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_4_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_4_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_4_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_4_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_4_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_4_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_5_aon_clk,
    input  wire                                    i_aic_5_aon_rst_n,
    input  wire                                    i_aic_5_clk,
    input  wire                                    i_aic_5_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_5_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_5_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_5_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_5_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_5_init_ht_axi_s_arlen,
    input  logic                                   i_aic_5_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_5_init_ht_axi_s_arprot,
    output logic                                   o_aic_5_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_5_init_ht_axi_s_arsize,
    input  logic                                   i_aic_5_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_5_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_5_init_ht_axi_s_rid,
    output logic                                   o_aic_5_init_ht_axi_s_rlast,
    input  logic                                   i_aic_5_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_5_init_ht_axi_s_rresp,
    output logic                                   o_aic_5_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_5_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_5_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_5_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_5_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_5_init_ht_axi_s_awlen,
    input  logic                                   i_aic_5_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_5_init_ht_axi_s_awprot,
    output logic                                   o_aic_5_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_5_init_ht_axi_s_awsize,
    input  logic                                   i_aic_5_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_5_init_ht_axi_s_bid,
    input  logic                                   i_aic_5_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_5_init_ht_axi_s_bresp,
    output logic                                   o_aic_5_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_5_init_ht_axi_s_wdata,
    input  logic                                   i_aic_5_init_ht_axi_s_wlast,
    output logic                                   o_aic_5_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_5_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_5_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_5_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_5_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_5_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_5_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_5_init_lt_axi_s_arlen,
    input  logic                                   i_aic_5_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_5_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_5_init_lt_axi_s_arqos,
    output logic                                   o_aic_5_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_5_init_lt_axi_s_arsize,
    input  logic                                   i_aic_5_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_5_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_5_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_5_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_5_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_5_init_lt_axi_s_awlen,
    input  logic                                   i_aic_5_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_5_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_5_init_lt_axi_s_awqos,
    output logic                                   o_aic_5_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_5_init_lt_axi_s_awsize,
    input  logic                                   i_aic_5_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_5_init_lt_axi_s_bid,
    input  logic                                   i_aic_5_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_5_init_lt_axi_s_bresp,
    output logic                                   o_aic_5_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_5_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_5_init_lt_axi_s_rid,
    output logic                                   o_aic_5_init_lt_axi_s_rlast,
    input  logic                                   i_aic_5_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_5_init_lt_axi_s_rresp,
    output logic                                   o_aic_5_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_5_init_lt_axi_s_wdata,
    input  logic                                   i_aic_5_init_lt_axi_s_wlast,
    output logic                                   o_aic_5_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_5_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_5_init_lt_axi_s_wvalid,
    output logic                                   o_aic_5_pwr_idle_val,
    output logic                                   o_aic_5_pwr_idle_ack,
    input  logic                                   i_aic_5_pwr_idle_req,
    input  wire                                    i_aic_5_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_5_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_5_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_5_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_5_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_5_targ_lt_axi_m_arlen,
    output logic                                   o_aic_5_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_5_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_5_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_5_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_5_targ_lt_axi_m_arsize,
    output logic                                   o_aic_5_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_5_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_5_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_5_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_5_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_5_targ_lt_axi_m_awlen,
    output logic                                   o_aic_5_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_5_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_5_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_5_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_5_targ_lt_axi_m_awsize,
    output logic                                   o_aic_5_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_5_targ_lt_axi_m_bid,
    output logic                                   o_aic_5_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_5_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_5_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_5_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_5_targ_lt_axi_m_rid,
    input  logic                                   i_aic_5_targ_lt_axi_m_rlast,
    output logic                                   o_aic_5_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_5_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_5_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_5_targ_lt_axi_m_wdata,
    output logic                                   o_aic_5_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_5_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_5_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_5_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_5_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_5_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_5_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_5_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_5_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_5_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_5_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_5_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_5_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_5_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_6_aon_clk,
    input  wire                                    i_aic_6_aon_rst_n,
    input  wire                                    i_aic_6_clk,
    input  wire                                    i_aic_6_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_6_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_6_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_6_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_6_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_6_init_ht_axi_s_arlen,
    input  logic                                   i_aic_6_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_6_init_ht_axi_s_arprot,
    output logic                                   o_aic_6_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_6_init_ht_axi_s_arsize,
    input  logic                                   i_aic_6_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_6_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_6_init_ht_axi_s_rid,
    output logic                                   o_aic_6_init_ht_axi_s_rlast,
    input  logic                                   i_aic_6_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_6_init_ht_axi_s_rresp,
    output logic                                   o_aic_6_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_6_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_6_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_6_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_6_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_6_init_ht_axi_s_awlen,
    input  logic                                   i_aic_6_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_6_init_ht_axi_s_awprot,
    output logic                                   o_aic_6_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_6_init_ht_axi_s_awsize,
    input  logic                                   i_aic_6_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_6_init_ht_axi_s_bid,
    input  logic                                   i_aic_6_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_6_init_ht_axi_s_bresp,
    output logic                                   o_aic_6_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_6_init_ht_axi_s_wdata,
    input  logic                                   i_aic_6_init_ht_axi_s_wlast,
    output logic                                   o_aic_6_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_6_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_6_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_6_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_6_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_6_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_6_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_6_init_lt_axi_s_arlen,
    input  logic                                   i_aic_6_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_6_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_6_init_lt_axi_s_arqos,
    output logic                                   o_aic_6_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_6_init_lt_axi_s_arsize,
    input  logic                                   i_aic_6_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_6_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_6_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_6_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_6_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_6_init_lt_axi_s_awlen,
    input  logic                                   i_aic_6_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_6_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_6_init_lt_axi_s_awqos,
    output logic                                   o_aic_6_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_6_init_lt_axi_s_awsize,
    input  logic                                   i_aic_6_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_6_init_lt_axi_s_bid,
    input  logic                                   i_aic_6_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_6_init_lt_axi_s_bresp,
    output logic                                   o_aic_6_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_6_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_6_init_lt_axi_s_rid,
    output logic                                   o_aic_6_init_lt_axi_s_rlast,
    input  logic                                   i_aic_6_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_6_init_lt_axi_s_rresp,
    output logic                                   o_aic_6_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_6_init_lt_axi_s_wdata,
    input  logic                                   i_aic_6_init_lt_axi_s_wlast,
    output logic                                   o_aic_6_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_6_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_6_init_lt_axi_s_wvalid,
    output logic                                   o_aic_6_pwr_idle_val,
    output logic                                   o_aic_6_pwr_idle_ack,
    input  logic                                   i_aic_6_pwr_idle_req,
    input  wire                                    i_aic_6_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_6_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_6_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_6_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_6_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_6_targ_lt_axi_m_arlen,
    output logic                                   o_aic_6_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_6_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_6_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_6_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_6_targ_lt_axi_m_arsize,
    output logic                                   o_aic_6_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_6_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_6_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_6_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_6_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_6_targ_lt_axi_m_awlen,
    output logic                                   o_aic_6_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_6_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_6_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_6_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_6_targ_lt_axi_m_awsize,
    output logic                                   o_aic_6_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_6_targ_lt_axi_m_bid,
    output logic                                   o_aic_6_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_6_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_6_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_6_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_6_targ_lt_axi_m_rid,
    input  logic                                   i_aic_6_targ_lt_axi_m_rlast,
    output logic                                   o_aic_6_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_6_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_6_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_6_targ_lt_axi_m_wdata,
    output logic                                   o_aic_6_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_6_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_6_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_6_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_6_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_6_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_6_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_6_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_6_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_6_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_6_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_6_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_6_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_6_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_7_aon_clk,
    input  wire                                    i_aic_7_aon_rst_n,
    input  wire                                    i_aic_7_clk,
    input  wire                                    i_aic_7_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_7_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_7_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_7_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_7_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_7_init_ht_axi_s_arlen,
    input  logic                                   i_aic_7_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_7_init_ht_axi_s_arprot,
    output logic                                   o_aic_7_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_7_init_ht_axi_s_arsize,
    input  logic                                   i_aic_7_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_7_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_7_init_ht_axi_s_rid,
    output logic                                   o_aic_7_init_ht_axi_s_rlast,
    input  logic                                   i_aic_7_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_7_init_ht_axi_s_rresp,
    output logic                                   o_aic_7_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_7_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_7_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_7_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_7_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_7_init_ht_axi_s_awlen,
    input  logic                                   i_aic_7_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_7_init_ht_axi_s_awprot,
    output logic                                   o_aic_7_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_7_init_ht_axi_s_awsize,
    input  logic                                   i_aic_7_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_7_init_ht_axi_s_bid,
    input  logic                                   i_aic_7_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_7_init_ht_axi_s_bresp,
    output logic                                   o_aic_7_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_7_init_ht_axi_s_wdata,
    input  logic                                   i_aic_7_init_ht_axi_s_wlast,
    output logic                                   o_aic_7_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_7_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_7_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_7_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_7_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_7_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_7_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_7_init_lt_axi_s_arlen,
    input  logic                                   i_aic_7_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_7_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_7_init_lt_axi_s_arqos,
    output logic                                   o_aic_7_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_7_init_lt_axi_s_arsize,
    input  logic                                   i_aic_7_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_7_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_7_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_7_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_7_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_7_init_lt_axi_s_awlen,
    input  logic                                   i_aic_7_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_7_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_7_init_lt_axi_s_awqos,
    output logic                                   o_aic_7_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_7_init_lt_axi_s_awsize,
    input  logic                                   i_aic_7_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_7_init_lt_axi_s_bid,
    input  logic                                   i_aic_7_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_7_init_lt_axi_s_bresp,
    output logic                                   o_aic_7_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_7_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_7_init_lt_axi_s_rid,
    output logic                                   o_aic_7_init_lt_axi_s_rlast,
    input  logic                                   i_aic_7_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_7_init_lt_axi_s_rresp,
    output logic                                   o_aic_7_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_7_init_lt_axi_s_wdata,
    input  logic                                   i_aic_7_init_lt_axi_s_wlast,
    output logic                                   o_aic_7_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_7_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_7_init_lt_axi_s_wvalid,
    output logic                                   o_aic_7_pwr_idle_val,
    output logic                                   o_aic_7_pwr_idle_ack,
    input  logic                                   i_aic_7_pwr_idle_req,
    input  wire                                    i_aic_7_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_7_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_7_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_7_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_7_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_7_targ_lt_axi_m_arlen,
    output logic                                   o_aic_7_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_7_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_7_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_7_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_7_targ_lt_axi_m_arsize,
    output logic                                   o_aic_7_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_7_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_7_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_7_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_7_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_7_targ_lt_axi_m_awlen,
    output logic                                   o_aic_7_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_7_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_7_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_7_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_7_targ_lt_axi_m_awsize,
    output logic                                   o_aic_7_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_7_targ_lt_axi_m_bid,
    output logic                                   o_aic_7_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_7_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_7_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_7_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_7_targ_lt_axi_m_rid,
    input  logic                                   i_aic_7_targ_lt_axi_m_rlast,
    output logic                                   o_aic_7_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_7_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_7_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_7_targ_lt_axi_m_wdata,
    output logic                                   o_aic_7_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_7_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_7_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_7_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_7_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_7_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_7_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_7_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_7_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_7_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_7_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_7_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_7_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_7_targ_syscfg_apb_m_pwrite,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld,
    input  logic [182:0]                           i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld,
    output logic [182:0]                           o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld,
    output logic [182:0]                           o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld,
    input  logic [182:0]                           i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld,
    input  wire                                    i_l2_4_aon_clk,
    input  wire                                    i_l2_4_aon_rst_n,
    input  wire                                    i_l2_4_clk,
    input  wire                                    i_l2_4_clken,
    output logic                                   o_l2_4_pwr_idle_val,
    output logic                                   o_l2_4_pwr_idle_ack,
    input  logic                                   i_l2_4_pwr_idle_req,
    input  wire                                    i_l2_4_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_4_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_4_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_4_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_4_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_4_targ_ht_axi_m_arlen,
    output logic                                   o_l2_4_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_4_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_4_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_4_targ_ht_axi_m_arsize,
    output logic                                   o_l2_4_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_4_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_4_targ_ht_axi_m_rid,
    input  logic                                   i_l2_4_targ_ht_axi_m_rlast,
    output logic                                   o_l2_4_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_4_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_4_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_4_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_4_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_4_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_4_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_4_targ_ht_axi_m_awlen,
    output logic                                   o_l2_4_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_4_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_4_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_4_targ_ht_axi_m_awsize,
    output logic                                   o_l2_4_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_4_targ_ht_axi_m_bid,
    output logic                                   o_l2_4_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_4_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_4_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_4_targ_ht_axi_m_wdata,
    output logic                                   o_l2_4_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_4_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_4_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_4_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_4_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_4_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_4_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_4_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_4_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_4_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_4_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_4_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_4_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_4_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_5_aon_clk,
    input  wire                                    i_l2_5_aon_rst_n,
    input  wire                                    i_l2_5_clk,
    input  wire                                    i_l2_5_clken,
    output logic                                   o_l2_5_pwr_idle_val,
    output logic                                   o_l2_5_pwr_idle_ack,
    input  logic                                   i_l2_5_pwr_idle_req,
    input  wire                                    i_l2_5_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_5_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_5_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_5_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_5_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_5_targ_ht_axi_m_arlen,
    output logic                                   o_l2_5_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_5_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_5_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_5_targ_ht_axi_m_arsize,
    output logic                                   o_l2_5_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_5_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_5_targ_ht_axi_m_rid,
    input  logic                                   i_l2_5_targ_ht_axi_m_rlast,
    output logic                                   o_l2_5_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_5_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_5_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_5_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_5_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_5_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_5_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_5_targ_ht_axi_m_awlen,
    output logic                                   o_l2_5_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_5_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_5_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_5_targ_ht_axi_m_awsize,
    output logic                                   o_l2_5_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_5_targ_ht_axi_m_bid,
    output logic                                   o_l2_5_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_5_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_5_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_5_targ_ht_axi_m_wdata,
    output logic                                   o_l2_5_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_5_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_5_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_5_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_5_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_5_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_5_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_5_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_5_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_5_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_5_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_5_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_5_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_5_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_6_aon_clk,
    input  wire                                    i_l2_6_aon_rst_n,
    input  wire                                    i_l2_6_clk,
    input  wire                                    i_l2_6_clken,
    output logic                                   o_l2_6_pwr_idle_val,
    output logic                                   o_l2_6_pwr_idle_ack,
    input  logic                                   i_l2_6_pwr_idle_req,
    input  wire                                    i_l2_6_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_6_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_6_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_6_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_6_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_6_targ_ht_axi_m_arlen,
    output logic                                   o_l2_6_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_6_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_6_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_6_targ_ht_axi_m_arsize,
    output logic                                   o_l2_6_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_6_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_6_targ_ht_axi_m_rid,
    input  logic                                   i_l2_6_targ_ht_axi_m_rlast,
    output logic                                   o_l2_6_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_6_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_6_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_6_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_6_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_6_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_6_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_6_targ_ht_axi_m_awlen,
    output logic                                   o_l2_6_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_6_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_6_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_6_targ_ht_axi_m_awsize,
    output logic                                   o_l2_6_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_6_targ_ht_axi_m_bid,
    output logic                                   o_l2_6_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_6_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_6_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_6_targ_ht_axi_m_wdata,
    output logic                                   o_l2_6_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_6_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_6_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_6_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_6_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_6_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_6_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_6_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_6_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_6_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_6_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_6_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_6_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_6_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_7_aon_clk,
    input  wire                                    i_l2_7_aon_rst_n,
    input  wire                                    i_l2_7_clk,
    input  wire                                    i_l2_7_clken,
    output logic                                   o_l2_7_pwr_idle_val,
    output logic                                   o_l2_7_pwr_idle_ack,
    input  logic                                   i_l2_7_pwr_idle_req,
    input  wire                                    i_l2_7_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_7_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_7_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_7_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_7_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_7_targ_ht_axi_m_arlen,
    output logic                                   o_l2_7_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_7_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_7_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_7_targ_ht_axi_m_arsize,
    output logic                                   o_l2_7_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_7_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_7_targ_ht_axi_m_rid,
    input  logic                                   i_l2_7_targ_ht_axi_m_rlast,
    output logic                                   o_l2_7_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_7_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_7_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_7_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_7_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_7_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_7_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_7_targ_ht_axi_m_awlen,
    output logic                                   o_l2_7_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_7_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_7_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_7_targ_ht_axi_m_awsize,
    output logic                                   o_l2_7_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_7_targ_ht_axi_m_bid,
    output logic                                   o_l2_7_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_7_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_7_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_7_targ_ht_axi_m_wdata,
    output logic                                   o_l2_7_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_7_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_7_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_7_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_7_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_7_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_7_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_7_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_7_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_7_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_7_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_7_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_7_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_7_targ_syscfg_apb_m_pwrite,
    input  logic                                   i_l2_addr_mode_port_b0,
    input  logic                                   i_l2_addr_mode_port_b1,
    input  logic                                   i_l2_intr_mode_port_b0,
    input  logic                                   i_l2_intr_mode_port_b1,
    input  logic                                   i_lpddr_graph_addr_mode_port_b0,
    input  logic                                   i_lpddr_graph_addr_mode_port_b1,
    input  logic                                   i_lpddr_graph_intr_mode_port_b0,
    input  logic                                   i_lpddr_graph_intr_mode_port_b1,
    input  logic                                   i_lpddr_ppp_addr_mode_port_b0,
    input  logic                                   i_lpddr_ppp_addr_mode_port_b1,
    input  logic                                   i_lpddr_ppp_intr_mode_port_b0,
    input  logic                                   i_lpddr_ppp_intr_mode_port_b1,
    input  wire                                    i_noc_clk,
    input  wire                                    i_noc_rst_n,
    input  logic                                   scan_en
);

    // Automated Address MSB fix: extra nets declaration
    logic[40:0] aic_4_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] aic_4_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_4_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] aic_4_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_4_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] aic_4_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] aic_5_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] aic_5_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_5_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] aic_5_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_5_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] aic_5_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] aic_6_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] aic_6_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_6_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] aic_6_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_6_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] aic_6_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] aic_7_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] aic_7_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_7_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] aic_7_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] aic_7_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] aic_7_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] l2_4_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] l2_4_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] l2_5_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] l2_5_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] l2_6_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] l2_6_targ_ht_axi_m_awaddr_msb_fixed;
    logic[40:0] l2_7_targ_ht_axi_m_araddr_msb_fixed;
    logic[40:0] l2_7_targ_ht_axi_m_awaddr_msb_fixed;

    // Automated Address MSB fix: Initiator-side assignments to extend addresses by 1 bit
    noc_common_addr_msb_setter u_addr_msb_fix_aic_4_init_ht (
        .i_axi_araddr_40b (i_aic_4_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (aic_4_init_ht_axi_s_araddr_msb_fixed)
    );
    assign aic_4_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_aic_4_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_4_init_lt (
        .i_axi_araddr_40b (i_aic_4_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (aic_4_init_lt_axi_s_araddr_msb_fixed)
    );
    assign aic_4_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_aic_4_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_5_init_ht (
        .i_axi_araddr_40b (i_aic_5_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (aic_5_init_ht_axi_s_araddr_msb_fixed)
    );
    assign aic_5_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_aic_5_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_5_init_lt (
        .i_axi_araddr_40b (i_aic_5_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (aic_5_init_lt_axi_s_araddr_msb_fixed)
    );
    assign aic_5_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_aic_5_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_6_init_ht (
        .i_axi_araddr_40b (i_aic_6_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (aic_6_init_ht_axi_s_araddr_msb_fixed)
    );
    assign aic_6_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_aic_6_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_6_init_lt (
        .i_axi_araddr_40b (i_aic_6_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (aic_6_init_lt_axi_s_araddr_msb_fixed)
    );
    assign aic_6_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_aic_6_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_7_init_ht (
        .i_axi_araddr_40b (i_aic_7_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (aic_7_init_ht_axi_s_araddr_msb_fixed)
    );
    assign aic_7_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_aic_7_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_aic_7_init_lt (
        .i_axi_araddr_40b (i_aic_7_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (aic_7_init_lt_axi_s_araddr_msb_fixed)
    );
    assign aic_7_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_aic_7_init_lt_axi_s_awaddr};

    // Automated Address MSB fix: Target-side assignments to drop unused MSB
    assign o_aic_4_targ_lt_axi_m_araddr = aic_4_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_aic_4_targ_lt_axi_m_awaddr = aic_4_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_aic_5_targ_lt_axi_m_araddr = aic_5_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_aic_5_targ_lt_axi_m_awaddr = aic_5_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_aic_6_targ_lt_axi_m_araddr = aic_6_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_aic_6_targ_lt_axi_m_awaddr = aic_6_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_aic_7_targ_lt_axi_m_araddr = aic_7_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_aic_7_targ_lt_axi_m_awaddr = aic_7_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_l2_4_targ_ht_axi_m_araddr = l2_4_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_l2_4_targ_ht_axi_m_awaddr = l2_4_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_l2_5_targ_ht_axi_m_araddr = l2_5_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_l2_5_targ_ht_axi_m_awaddr = l2_5_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_l2_6_targ_ht_axi_m_araddr = l2_6_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_l2_6_targ_ht_axi_m_awaddr = l2_6_targ_ht_axi_m_awaddr_msb_fixed[39:0];
    assign o_l2_7_targ_ht_axi_m_araddr = l2_7_targ_ht_axi_m_araddr_msb_fixed[39:0];
    assign o_l2_7_targ_ht_axi_m_awaddr = l2_7_targ_ht_axi_m_awaddr_msb_fixed[39:0];


    noc_art_h_north u_noc_art_h_north (
    .aic_4_aon_clk(i_aic_4_aon_clk),
    .aic_4_aon_rst_n(i_aic_4_aon_rst_n),
    .aic_4_clk(i_aic_4_clk),
    .aic_4_clken(i_aic_4_clken),
    .aic_4_init_ht_rd_Ar_Addr(aic_4_init_ht_axi_s_araddr_msb_fixed),
    .aic_4_init_ht_rd_Ar_Burst(i_aic_4_init_ht_axi_s_arburst),
    .aic_4_init_ht_rd_Ar_Cache(i_aic_4_init_ht_axi_s_arcache),
    .aic_4_init_ht_rd_Ar_Id(i_aic_4_init_ht_axi_s_arid),
    .aic_4_init_ht_rd_Ar_Len(i_aic_4_init_ht_axi_s_arlen),
    .aic_4_init_ht_rd_Ar_Lock(i_aic_4_init_ht_axi_s_arlock),
    .aic_4_init_ht_rd_Ar_Prot(i_aic_4_init_ht_axi_s_arprot),
    .aic_4_init_ht_rd_Ar_Ready(o_aic_4_init_ht_axi_s_arready),
    .aic_4_init_ht_rd_Ar_Size(i_aic_4_init_ht_axi_s_arsize),
    .aic_4_init_ht_rd_Ar_Valid(i_aic_4_init_ht_axi_s_arvalid),
    .aic_4_init_ht_rd_R_Data(o_aic_4_init_ht_axi_s_rdata),
    .aic_4_init_ht_rd_R_Id(o_aic_4_init_ht_axi_s_rid),
    .aic_4_init_ht_rd_R_Last(o_aic_4_init_ht_axi_s_rlast),
    .aic_4_init_ht_rd_R_Ready(i_aic_4_init_ht_axi_s_rready),
    .aic_4_init_ht_rd_R_Resp(o_aic_4_init_ht_axi_s_rresp),
    .aic_4_init_ht_rd_R_Valid(o_aic_4_init_ht_axi_s_rvalid),
    .aic_4_init_ht_wr_Aw_Addr(aic_4_init_ht_axi_s_awaddr_msb_fixed),
    .aic_4_init_ht_wr_Aw_Burst(i_aic_4_init_ht_axi_s_awburst),
    .aic_4_init_ht_wr_Aw_Cache(i_aic_4_init_ht_axi_s_awcache),
    .aic_4_init_ht_wr_Aw_Id(i_aic_4_init_ht_axi_s_awid),
    .aic_4_init_ht_wr_Aw_Len(i_aic_4_init_ht_axi_s_awlen),
    .aic_4_init_ht_wr_Aw_Lock(i_aic_4_init_ht_axi_s_awlock),
    .aic_4_init_ht_wr_Aw_Prot(i_aic_4_init_ht_axi_s_awprot),
    .aic_4_init_ht_wr_Aw_Ready(o_aic_4_init_ht_axi_s_awready),
    .aic_4_init_ht_wr_Aw_Size(i_aic_4_init_ht_axi_s_awsize),
    .aic_4_init_ht_wr_Aw_Valid(i_aic_4_init_ht_axi_s_awvalid),
    .aic_4_init_ht_wr_B_Id(o_aic_4_init_ht_axi_s_bid),
    .aic_4_init_ht_wr_B_Ready(i_aic_4_init_ht_axi_s_bready),
    .aic_4_init_ht_wr_B_Resp(o_aic_4_init_ht_axi_s_bresp),
    .aic_4_init_ht_wr_B_Valid(o_aic_4_init_ht_axi_s_bvalid),
    .aic_4_init_ht_wr_W_Data(i_aic_4_init_ht_axi_s_wdata),
    .aic_4_init_ht_wr_W_Last(i_aic_4_init_ht_axi_s_wlast),
    .aic_4_init_ht_wr_W_Ready(o_aic_4_init_ht_axi_s_wready),
    .aic_4_init_ht_wr_W_Strb(i_aic_4_init_ht_axi_s_wstrb),
    .aic_4_init_ht_wr_W_Valid(i_aic_4_init_ht_axi_s_wvalid),
    .aic_4_init_lt_Ar_Addr(aic_4_init_lt_axi_s_araddr_msb_fixed),
    .aic_4_init_lt_Ar_Burst(i_aic_4_init_lt_axi_s_arburst),
    .aic_4_init_lt_Ar_Cache(i_aic_4_init_lt_axi_s_arcache),
    .aic_4_init_lt_Ar_Id(i_aic_4_init_lt_axi_s_arid),
    .aic_4_init_lt_Ar_Len(i_aic_4_init_lt_axi_s_arlen),
    .aic_4_init_lt_Ar_Lock(i_aic_4_init_lt_axi_s_arlock),
    .aic_4_init_lt_Ar_Prot(i_aic_4_init_lt_axi_s_arprot),
    .aic_4_init_lt_Ar_Qos(i_aic_4_init_lt_axi_s_arqos),
    .aic_4_init_lt_Ar_Ready(o_aic_4_init_lt_axi_s_arready),
    .aic_4_init_lt_Ar_Size(i_aic_4_init_lt_axi_s_arsize),
    .aic_4_init_lt_Ar_Valid(i_aic_4_init_lt_axi_s_arvalid),
    .aic_4_init_lt_Aw_Addr(aic_4_init_lt_axi_s_awaddr_msb_fixed),
    .aic_4_init_lt_Aw_Burst(i_aic_4_init_lt_axi_s_awburst),
    .aic_4_init_lt_Aw_Cache(i_aic_4_init_lt_axi_s_awcache),
    .aic_4_init_lt_Aw_Id(i_aic_4_init_lt_axi_s_awid),
    .aic_4_init_lt_Aw_Len(i_aic_4_init_lt_axi_s_awlen),
    .aic_4_init_lt_Aw_Lock(i_aic_4_init_lt_axi_s_awlock),
    .aic_4_init_lt_Aw_Prot(i_aic_4_init_lt_axi_s_awprot),
    .aic_4_init_lt_Aw_Qos(i_aic_4_init_lt_axi_s_awqos),
    .aic_4_init_lt_Aw_Ready(o_aic_4_init_lt_axi_s_awready),
    .aic_4_init_lt_Aw_Size(i_aic_4_init_lt_axi_s_awsize),
    .aic_4_init_lt_Aw_Valid(i_aic_4_init_lt_axi_s_awvalid),
    .aic_4_init_lt_B_Id(o_aic_4_init_lt_axi_s_bid),
    .aic_4_init_lt_B_Ready(i_aic_4_init_lt_axi_s_bready),
    .aic_4_init_lt_B_Resp(o_aic_4_init_lt_axi_s_bresp),
    .aic_4_init_lt_B_Valid(o_aic_4_init_lt_axi_s_bvalid),
    .aic_4_init_lt_R_Data(o_aic_4_init_lt_axi_s_rdata),
    .aic_4_init_lt_R_Id(o_aic_4_init_lt_axi_s_rid),
    .aic_4_init_lt_R_Last(o_aic_4_init_lt_axi_s_rlast),
    .aic_4_init_lt_R_Ready(i_aic_4_init_lt_axi_s_rready),
    .aic_4_init_lt_R_Resp(o_aic_4_init_lt_axi_s_rresp),
    .aic_4_init_lt_R_Valid(o_aic_4_init_lt_axi_s_rvalid),
    .aic_4_init_lt_W_Data(i_aic_4_init_lt_axi_s_wdata),
    .aic_4_init_lt_W_Last(i_aic_4_init_lt_axi_s_wlast),
    .aic_4_init_lt_W_Ready(o_aic_4_init_lt_axi_s_wready),
    .aic_4_init_lt_W_Strb(i_aic_4_init_lt_axi_s_wstrb),
    .aic_4_init_lt_W_Valid(i_aic_4_init_lt_axi_s_wvalid),
    .aic_4_pwr_Idle(o_aic_4_pwr_idle_val),
    .aic_4_pwr_IdleAck(o_aic_4_pwr_idle_ack),
    .aic_4_pwr_IdleReq(i_aic_4_pwr_idle_req),
    .aic_4_rst_n(i_aic_4_rst_n),
    .aic_4_targ_lt_Ar_Addr(aic_4_targ_lt_axi_m_araddr_msb_fixed),
    .aic_4_targ_lt_Ar_Burst(o_aic_4_targ_lt_axi_m_arburst),
    .aic_4_targ_lt_Ar_Cache(o_aic_4_targ_lt_axi_m_arcache),
    .aic_4_targ_lt_Ar_Id(o_aic_4_targ_lt_axi_m_arid),
    .aic_4_targ_lt_Ar_Len(o_aic_4_targ_lt_axi_m_arlen),
    .aic_4_targ_lt_Ar_Lock(o_aic_4_targ_lt_axi_m_arlock),
    .aic_4_targ_lt_Ar_Prot(o_aic_4_targ_lt_axi_m_arprot),
    .aic_4_targ_lt_Ar_Qos(o_aic_4_targ_lt_axi_m_arqos),
    .aic_4_targ_lt_Ar_Ready(i_aic_4_targ_lt_axi_m_arready),
    .aic_4_targ_lt_Ar_Size(o_aic_4_targ_lt_axi_m_arsize),
    .aic_4_targ_lt_Ar_Valid(o_aic_4_targ_lt_axi_m_arvalid),
    .aic_4_targ_lt_Aw_Addr(aic_4_targ_lt_axi_m_awaddr_msb_fixed),
    .aic_4_targ_lt_Aw_Burst(o_aic_4_targ_lt_axi_m_awburst),
    .aic_4_targ_lt_Aw_Cache(o_aic_4_targ_lt_axi_m_awcache),
    .aic_4_targ_lt_Aw_Id(o_aic_4_targ_lt_axi_m_awid),
    .aic_4_targ_lt_Aw_Len(o_aic_4_targ_lt_axi_m_awlen),
    .aic_4_targ_lt_Aw_Lock(o_aic_4_targ_lt_axi_m_awlock),
    .aic_4_targ_lt_Aw_Prot(o_aic_4_targ_lt_axi_m_awprot),
    .aic_4_targ_lt_Aw_Qos(o_aic_4_targ_lt_axi_m_awqos),
    .aic_4_targ_lt_Aw_Ready(i_aic_4_targ_lt_axi_m_awready),
    .aic_4_targ_lt_Aw_Size(o_aic_4_targ_lt_axi_m_awsize),
    .aic_4_targ_lt_Aw_Valid(o_aic_4_targ_lt_axi_m_awvalid),
    .aic_4_targ_lt_B_Id(i_aic_4_targ_lt_axi_m_bid),
    .aic_4_targ_lt_B_Ready(o_aic_4_targ_lt_axi_m_bready),
    .aic_4_targ_lt_B_Resp(i_aic_4_targ_lt_axi_m_bresp),
    .aic_4_targ_lt_B_Valid(i_aic_4_targ_lt_axi_m_bvalid),
    .aic_4_targ_lt_R_Data(i_aic_4_targ_lt_axi_m_rdata),
    .aic_4_targ_lt_R_Id(i_aic_4_targ_lt_axi_m_rid),
    .aic_4_targ_lt_R_Last(i_aic_4_targ_lt_axi_m_rlast),
    .aic_4_targ_lt_R_Ready(o_aic_4_targ_lt_axi_m_rready),
    .aic_4_targ_lt_R_Resp(i_aic_4_targ_lt_axi_m_rresp),
    .aic_4_targ_lt_R_Valid(i_aic_4_targ_lt_axi_m_rvalid),
    .aic_4_targ_lt_W_Data(o_aic_4_targ_lt_axi_m_wdata),
    .aic_4_targ_lt_W_Last(o_aic_4_targ_lt_axi_m_wlast),
    .aic_4_targ_lt_W_Ready(i_aic_4_targ_lt_axi_m_wready),
    .aic_4_targ_lt_W_Strb(o_aic_4_targ_lt_axi_m_wstrb),
    .aic_4_targ_lt_W_Valid(o_aic_4_targ_lt_axi_m_wvalid),
    .aic_4_targ_syscfg_PAddr(o_aic_4_targ_syscfg_apb_m_paddr),
    .aic_4_targ_syscfg_PEnable(o_aic_4_targ_syscfg_apb_m_penable),
    .aic_4_targ_syscfg_PProt(o_aic_4_targ_syscfg_apb_m_pprot),
    .aic_4_targ_syscfg_PRData(i_aic_4_targ_syscfg_apb_m_prdata),
    .aic_4_targ_syscfg_PReady(i_aic_4_targ_syscfg_apb_m_pready),
    .aic_4_targ_syscfg_PSel(o_aic_4_targ_syscfg_apb_m_psel),
    .aic_4_targ_syscfg_PSlvErr(i_aic_4_targ_syscfg_apb_m_pslverr),
    .aic_4_targ_syscfg_PStrb(o_aic_4_targ_syscfg_apb_m_pstrb),
    .aic_4_targ_syscfg_PWData(o_aic_4_targ_syscfg_apb_m_pwdata),
    .aic_4_targ_syscfg_PWrite(o_aic_4_targ_syscfg_apb_m_pwrite),
    .aic_5_aon_clk(i_aic_5_aon_clk),
    .aic_5_aon_rst_n(i_aic_5_aon_rst_n),
    .aic_5_clk(i_aic_5_clk),
    .aic_5_clken(i_aic_5_clken),
    .aic_5_init_ht_rd_Ar_Addr(aic_5_init_ht_axi_s_araddr_msb_fixed),
    .aic_5_init_ht_rd_Ar_Burst(i_aic_5_init_ht_axi_s_arburst),
    .aic_5_init_ht_rd_Ar_Cache(i_aic_5_init_ht_axi_s_arcache),
    .aic_5_init_ht_rd_Ar_Id(i_aic_5_init_ht_axi_s_arid),
    .aic_5_init_ht_rd_Ar_Len(i_aic_5_init_ht_axi_s_arlen),
    .aic_5_init_ht_rd_Ar_Lock(i_aic_5_init_ht_axi_s_arlock),
    .aic_5_init_ht_rd_Ar_Prot(i_aic_5_init_ht_axi_s_arprot),
    .aic_5_init_ht_rd_Ar_Ready(o_aic_5_init_ht_axi_s_arready),
    .aic_5_init_ht_rd_Ar_Size(i_aic_5_init_ht_axi_s_arsize),
    .aic_5_init_ht_rd_Ar_Valid(i_aic_5_init_ht_axi_s_arvalid),
    .aic_5_init_ht_rd_R_Data(o_aic_5_init_ht_axi_s_rdata),
    .aic_5_init_ht_rd_R_Id(o_aic_5_init_ht_axi_s_rid),
    .aic_5_init_ht_rd_R_Last(o_aic_5_init_ht_axi_s_rlast),
    .aic_5_init_ht_rd_R_Ready(i_aic_5_init_ht_axi_s_rready),
    .aic_5_init_ht_rd_R_Resp(o_aic_5_init_ht_axi_s_rresp),
    .aic_5_init_ht_rd_R_Valid(o_aic_5_init_ht_axi_s_rvalid),
    .aic_5_init_ht_wr_Aw_Addr(aic_5_init_ht_axi_s_awaddr_msb_fixed),
    .aic_5_init_ht_wr_Aw_Burst(i_aic_5_init_ht_axi_s_awburst),
    .aic_5_init_ht_wr_Aw_Cache(i_aic_5_init_ht_axi_s_awcache),
    .aic_5_init_ht_wr_Aw_Id(i_aic_5_init_ht_axi_s_awid),
    .aic_5_init_ht_wr_Aw_Len(i_aic_5_init_ht_axi_s_awlen),
    .aic_5_init_ht_wr_Aw_Lock(i_aic_5_init_ht_axi_s_awlock),
    .aic_5_init_ht_wr_Aw_Prot(i_aic_5_init_ht_axi_s_awprot),
    .aic_5_init_ht_wr_Aw_Ready(o_aic_5_init_ht_axi_s_awready),
    .aic_5_init_ht_wr_Aw_Size(i_aic_5_init_ht_axi_s_awsize),
    .aic_5_init_ht_wr_Aw_Valid(i_aic_5_init_ht_axi_s_awvalid),
    .aic_5_init_ht_wr_B_Id(o_aic_5_init_ht_axi_s_bid),
    .aic_5_init_ht_wr_B_Ready(i_aic_5_init_ht_axi_s_bready),
    .aic_5_init_ht_wr_B_Resp(o_aic_5_init_ht_axi_s_bresp),
    .aic_5_init_ht_wr_B_Valid(o_aic_5_init_ht_axi_s_bvalid),
    .aic_5_init_ht_wr_W_Data(i_aic_5_init_ht_axi_s_wdata),
    .aic_5_init_ht_wr_W_Last(i_aic_5_init_ht_axi_s_wlast),
    .aic_5_init_ht_wr_W_Ready(o_aic_5_init_ht_axi_s_wready),
    .aic_5_init_ht_wr_W_Strb(i_aic_5_init_ht_axi_s_wstrb),
    .aic_5_init_ht_wr_W_Valid(i_aic_5_init_ht_axi_s_wvalid),
    .aic_5_init_lt_Ar_Addr(aic_5_init_lt_axi_s_araddr_msb_fixed),
    .aic_5_init_lt_Ar_Burst(i_aic_5_init_lt_axi_s_arburst),
    .aic_5_init_lt_Ar_Cache(i_aic_5_init_lt_axi_s_arcache),
    .aic_5_init_lt_Ar_Id(i_aic_5_init_lt_axi_s_arid),
    .aic_5_init_lt_Ar_Len(i_aic_5_init_lt_axi_s_arlen),
    .aic_5_init_lt_Ar_Lock(i_aic_5_init_lt_axi_s_arlock),
    .aic_5_init_lt_Ar_Prot(i_aic_5_init_lt_axi_s_arprot),
    .aic_5_init_lt_Ar_Qos(i_aic_5_init_lt_axi_s_arqos),
    .aic_5_init_lt_Ar_Ready(o_aic_5_init_lt_axi_s_arready),
    .aic_5_init_lt_Ar_Size(i_aic_5_init_lt_axi_s_arsize),
    .aic_5_init_lt_Ar_Valid(i_aic_5_init_lt_axi_s_arvalid),
    .aic_5_init_lt_Aw_Addr(aic_5_init_lt_axi_s_awaddr_msb_fixed),
    .aic_5_init_lt_Aw_Burst(i_aic_5_init_lt_axi_s_awburst),
    .aic_5_init_lt_Aw_Cache(i_aic_5_init_lt_axi_s_awcache),
    .aic_5_init_lt_Aw_Id(i_aic_5_init_lt_axi_s_awid),
    .aic_5_init_lt_Aw_Len(i_aic_5_init_lt_axi_s_awlen),
    .aic_5_init_lt_Aw_Lock(i_aic_5_init_lt_axi_s_awlock),
    .aic_5_init_lt_Aw_Prot(i_aic_5_init_lt_axi_s_awprot),
    .aic_5_init_lt_Aw_Qos(i_aic_5_init_lt_axi_s_awqos),
    .aic_5_init_lt_Aw_Ready(o_aic_5_init_lt_axi_s_awready),
    .aic_5_init_lt_Aw_Size(i_aic_5_init_lt_axi_s_awsize),
    .aic_5_init_lt_Aw_Valid(i_aic_5_init_lt_axi_s_awvalid),
    .aic_5_init_lt_B_Id(o_aic_5_init_lt_axi_s_bid),
    .aic_5_init_lt_B_Ready(i_aic_5_init_lt_axi_s_bready),
    .aic_5_init_lt_B_Resp(o_aic_5_init_lt_axi_s_bresp),
    .aic_5_init_lt_B_Valid(o_aic_5_init_lt_axi_s_bvalid),
    .aic_5_init_lt_R_Data(o_aic_5_init_lt_axi_s_rdata),
    .aic_5_init_lt_R_Id(o_aic_5_init_lt_axi_s_rid),
    .aic_5_init_lt_R_Last(o_aic_5_init_lt_axi_s_rlast),
    .aic_5_init_lt_R_Ready(i_aic_5_init_lt_axi_s_rready),
    .aic_5_init_lt_R_Resp(o_aic_5_init_lt_axi_s_rresp),
    .aic_5_init_lt_R_Valid(o_aic_5_init_lt_axi_s_rvalid),
    .aic_5_init_lt_W_Data(i_aic_5_init_lt_axi_s_wdata),
    .aic_5_init_lt_W_Last(i_aic_5_init_lt_axi_s_wlast),
    .aic_5_init_lt_W_Ready(o_aic_5_init_lt_axi_s_wready),
    .aic_5_init_lt_W_Strb(i_aic_5_init_lt_axi_s_wstrb),
    .aic_5_init_lt_W_Valid(i_aic_5_init_lt_axi_s_wvalid),
    .aic_5_pwr_Idle(o_aic_5_pwr_idle_val),
    .aic_5_pwr_IdleAck(o_aic_5_pwr_idle_ack),
    .aic_5_pwr_IdleReq(i_aic_5_pwr_idle_req),
    .aic_5_rst_n(i_aic_5_rst_n),
    .aic_5_targ_lt_Ar_Addr(aic_5_targ_lt_axi_m_araddr_msb_fixed),
    .aic_5_targ_lt_Ar_Burst(o_aic_5_targ_lt_axi_m_arburst),
    .aic_5_targ_lt_Ar_Cache(o_aic_5_targ_lt_axi_m_arcache),
    .aic_5_targ_lt_Ar_Id(o_aic_5_targ_lt_axi_m_arid),
    .aic_5_targ_lt_Ar_Len(o_aic_5_targ_lt_axi_m_arlen),
    .aic_5_targ_lt_Ar_Lock(o_aic_5_targ_lt_axi_m_arlock),
    .aic_5_targ_lt_Ar_Prot(o_aic_5_targ_lt_axi_m_arprot),
    .aic_5_targ_lt_Ar_Qos(o_aic_5_targ_lt_axi_m_arqos),
    .aic_5_targ_lt_Ar_Ready(i_aic_5_targ_lt_axi_m_arready),
    .aic_5_targ_lt_Ar_Size(o_aic_5_targ_lt_axi_m_arsize),
    .aic_5_targ_lt_Ar_Valid(o_aic_5_targ_lt_axi_m_arvalid),
    .aic_5_targ_lt_Aw_Addr(aic_5_targ_lt_axi_m_awaddr_msb_fixed),
    .aic_5_targ_lt_Aw_Burst(o_aic_5_targ_lt_axi_m_awburst),
    .aic_5_targ_lt_Aw_Cache(o_aic_5_targ_lt_axi_m_awcache),
    .aic_5_targ_lt_Aw_Id(o_aic_5_targ_lt_axi_m_awid),
    .aic_5_targ_lt_Aw_Len(o_aic_5_targ_lt_axi_m_awlen),
    .aic_5_targ_lt_Aw_Lock(o_aic_5_targ_lt_axi_m_awlock),
    .aic_5_targ_lt_Aw_Prot(o_aic_5_targ_lt_axi_m_awprot),
    .aic_5_targ_lt_Aw_Qos(o_aic_5_targ_lt_axi_m_awqos),
    .aic_5_targ_lt_Aw_Ready(i_aic_5_targ_lt_axi_m_awready),
    .aic_5_targ_lt_Aw_Size(o_aic_5_targ_lt_axi_m_awsize),
    .aic_5_targ_lt_Aw_Valid(o_aic_5_targ_lt_axi_m_awvalid),
    .aic_5_targ_lt_B_Id(i_aic_5_targ_lt_axi_m_bid),
    .aic_5_targ_lt_B_Ready(o_aic_5_targ_lt_axi_m_bready),
    .aic_5_targ_lt_B_Resp(i_aic_5_targ_lt_axi_m_bresp),
    .aic_5_targ_lt_B_Valid(i_aic_5_targ_lt_axi_m_bvalid),
    .aic_5_targ_lt_R_Data(i_aic_5_targ_lt_axi_m_rdata),
    .aic_5_targ_lt_R_Id(i_aic_5_targ_lt_axi_m_rid),
    .aic_5_targ_lt_R_Last(i_aic_5_targ_lt_axi_m_rlast),
    .aic_5_targ_lt_R_Ready(o_aic_5_targ_lt_axi_m_rready),
    .aic_5_targ_lt_R_Resp(i_aic_5_targ_lt_axi_m_rresp),
    .aic_5_targ_lt_R_Valid(i_aic_5_targ_lt_axi_m_rvalid),
    .aic_5_targ_lt_W_Data(o_aic_5_targ_lt_axi_m_wdata),
    .aic_5_targ_lt_W_Last(o_aic_5_targ_lt_axi_m_wlast),
    .aic_5_targ_lt_W_Ready(i_aic_5_targ_lt_axi_m_wready),
    .aic_5_targ_lt_W_Strb(o_aic_5_targ_lt_axi_m_wstrb),
    .aic_5_targ_lt_W_Valid(o_aic_5_targ_lt_axi_m_wvalid),
    .aic_5_targ_syscfg_PAddr(o_aic_5_targ_syscfg_apb_m_paddr),
    .aic_5_targ_syscfg_PEnable(o_aic_5_targ_syscfg_apb_m_penable),
    .aic_5_targ_syscfg_PProt(o_aic_5_targ_syscfg_apb_m_pprot),
    .aic_5_targ_syscfg_PRData(i_aic_5_targ_syscfg_apb_m_prdata),
    .aic_5_targ_syscfg_PReady(i_aic_5_targ_syscfg_apb_m_pready),
    .aic_5_targ_syscfg_PSel(o_aic_5_targ_syscfg_apb_m_psel),
    .aic_5_targ_syscfg_PSlvErr(i_aic_5_targ_syscfg_apb_m_pslverr),
    .aic_5_targ_syscfg_PStrb(o_aic_5_targ_syscfg_apb_m_pstrb),
    .aic_5_targ_syscfg_PWData(o_aic_5_targ_syscfg_apb_m_pwdata),
    .aic_5_targ_syscfg_PWrite(o_aic_5_targ_syscfg_apb_m_pwrite),
    .aic_6_aon_clk(i_aic_6_aon_clk),
    .aic_6_aon_rst_n(i_aic_6_aon_rst_n),
    .aic_6_clk(i_aic_6_clk),
    .aic_6_clken(i_aic_6_clken),
    .aic_6_init_ht_rd_Ar_Addr(aic_6_init_ht_axi_s_araddr_msb_fixed),
    .aic_6_init_ht_rd_Ar_Burst(i_aic_6_init_ht_axi_s_arburst),
    .aic_6_init_ht_rd_Ar_Cache(i_aic_6_init_ht_axi_s_arcache),
    .aic_6_init_ht_rd_Ar_Id(i_aic_6_init_ht_axi_s_arid),
    .aic_6_init_ht_rd_Ar_Len(i_aic_6_init_ht_axi_s_arlen),
    .aic_6_init_ht_rd_Ar_Lock(i_aic_6_init_ht_axi_s_arlock),
    .aic_6_init_ht_rd_Ar_Prot(i_aic_6_init_ht_axi_s_arprot),
    .aic_6_init_ht_rd_Ar_Ready(o_aic_6_init_ht_axi_s_arready),
    .aic_6_init_ht_rd_Ar_Size(i_aic_6_init_ht_axi_s_arsize),
    .aic_6_init_ht_rd_Ar_Valid(i_aic_6_init_ht_axi_s_arvalid),
    .aic_6_init_ht_rd_R_Data(o_aic_6_init_ht_axi_s_rdata),
    .aic_6_init_ht_rd_R_Id(o_aic_6_init_ht_axi_s_rid),
    .aic_6_init_ht_rd_R_Last(o_aic_6_init_ht_axi_s_rlast),
    .aic_6_init_ht_rd_R_Ready(i_aic_6_init_ht_axi_s_rready),
    .aic_6_init_ht_rd_R_Resp(o_aic_6_init_ht_axi_s_rresp),
    .aic_6_init_ht_rd_R_Valid(o_aic_6_init_ht_axi_s_rvalid),
    .aic_6_init_ht_wr_Aw_Addr(aic_6_init_ht_axi_s_awaddr_msb_fixed),
    .aic_6_init_ht_wr_Aw_Burst(i_aic_6_init_ht_axi_s_awburst),
    .aic_6_init_ht_wr_Aw_Cache(i_aic_6_init_ht_axi_s_awcache),
    .aic_6_init_ht_wr_Aw_Id(i_aic_6_init_ht_axi_s_awid),
    .aic_6_init_ht_wr_Aw_Len(i_aic_6_init_ht_axi_s_awlen),
    .aic_6_init_ht_wr_Aw_Lock(i_aic_6_init_ht_axi_s_awlock),
    .aic_6_init_ht_wr_Aw_Prot(i_aic_6_init_ht_axi_s_awprot),
    .aic_6_init_ht_wr_Aw_Ready(o_aic_6_init_ht_axi_s_awready),
    .aic_6_init_ht_wr_Aw_Size(i_aic_6_init_ht_axi_s_awsize),
    .aic_6_init_ht_wr_Aw_Valid(i_aic_6_init_ht_axi_s_awvalid),
    .aic_6_init_ht_wr_B_Id(o_aic_6_init_ht_axi_s_bid),
    .aic_6_init_ht_wr_B_Ready(i_aic_6_init_ht_axi_s_bready),
    .aic_6_init_ht_wr_B_Resp(o_aic_6_init_ht_axi_s_bresp),
    .aic_6_init_ht_wr_B_Valid(o_aic_6_init_ht_axi_s_bvalid),
    .aic_6_init_ht_wr_W_Data(i_aic_6_init_ht_axi_s_wdata),
    .aic_6_init_ht_wr_W_Last(i_aic_6_init_ht_axi_s_wlast),
    .aic_6_init_ht_wr_W_Ready(o_aic_6_init_ht_axi_s_wready),
    .aic_6_init_ht_wr_W_Strb(i_aic_6_init_ht_axi_s_wstrb),
    .aic_6_init_ht_wr_W_Valid(i_aic_6_init_ht_axi_s_wvalid),
    .aic_6_init_lt_Ar_Addr(aic_6_init_lt_axi_s_araddr_msb_fixed),
    .aic_6_init_lt_Ar_Burst(i_aic_6_init_lt_axi_s_arburst),
    .aic_6_init_lt_Ar_Cache(i_aic_6_init_lt_axi_s_arcache),
    .aic_6_init_lt_Ar_Id(i_aic_6_init_lt_axi_s_arid),
    .aic_6_init_lt_Ar_Len(i_aic_6_init_lt_axi_s_arlen),
    .aic_6_init_lt_Ar_Lock(i_aic_6_init_lt_axi_s_arlock),
    .aic_6_init_lt_Ar_Prot(i_aic_6_init_lt_axi_s_arprot),
    .aic_6_init_lt_Ar_Qos(i_aic_6_init_lt_axi_s_arqos),
    .aic_6_init_lt_Ar_Ready(o_aic_6_init_lt_axi_s_arready),
    .aic_6_init_lt_Ar_Size(i_aic_6_init_lt_axi_s_arsize),
    .aic_6_init_lt_Ar_Valid(i_aic_6_init_lt_axi_s_arvalid),
    .aic_6_init_lt_Aw_Addr(aic_6_init_lt_axi_s_awaddr_msb_fixed),
    .aic_6_init_lt_Aw_Burst(i_aic_6_init_lt_axi_s_awburst),
    .aic_6_init_lt_Aw_Cache(i_aic_6_init_lt_axi_s_awcache),
    .aic_6_init_lt_Aw_Id(i_aic_6_init_lt_axi_s_awid),
    .aic_6_init_lt_Aw_Len(i_aic_6_init_lt_axi_s_awlen),
    .aic_6_init_lt_Aw_Lock(i_aic_6_init_lt_axi_s_awlock),
    .aic_6_init_lt_Aw_Prot(i_aic_6_init_lt_axi_s_awprot),
    .aic_6_init_lt_Aw_Qos(i_aic_6_init_lt_axi_s_awqos),
    .aic_6_init_lt_Aw_Ready(o_aic_6_init_lt_axi_s_awready),
    .aic_6_init_lt_Aw_Size(i_aic_6_init_lt_axi_s_awsize),
    .aic_6_init_lt_Aw_Valid(i_aic_6_init_lt_axi_s_awvalid),
    .aic_6_init_lt_B_Id(o_aic_6_init_lt_axi_s_bid),
    .aic_6_init_lt_B_Ready(i_aic_6_init_lt_axi_s_bready),
    .aic_6_init_lt_B_Resp(o_aic_6_init_lt_axi_s_bresp),
    .aic_6_init_lt_B_Valid(o_aic_6_init_lt_axi_s_bvalid),
    .aic_6_init_lt_R_Data(o_aic_6_init_lt_axi_s_rdata),
    .aic_6_init_lt_R_Id(o_aic_6_init_lt_axi_s_rid),
    .aic_6_init_lt_R_Last(o_aic_6_init_lt_axi_s_rlast),
    .aic_6_init_lt_R_Ready(i_aic_6_init_lt_axi_s_rready),
    .aic_6_init_lt_R_Resp(o_aic_6_init_lt_axi_s_rresp),
    .aic_6_init_lt_R_Valid(o_aic_6_init_lt_axi_s_rvalid),
    .aic_6_init_lt_W_Data(i_aic_6_init_lt_axi_s_wdata),
    .aic_6_init_lt_W_Last(i_aic_6_init_lt_axi_s_wlast),
    .aic_6_init_lt_W_Ready(o_aic_6_init_lt_axi_s_wready),
    .aic_6_init_lt_W_Strb(i_aic_6_init_lt_axi_s_wstrb),
    .aic_6_init_lt_W_Valid(i_aic_6_init_lt_axi_s_wvalid),
    .aic_6_pwr_Idle(o_aic_6_pwr_idle_val),
    .aic_6_pwr_IdleAck(o_aic_6_pwr_idle_ack),
    .aic_6_pwr_IdleReq(i_aic_6_pwr_idle_req),
    .aic_6_rst_n(i_aic_6_rst_n),
    .aic_6_targ_lt_Ar_Addr(aic_6_targ_lt_axi_m_araddr_msb_fixed),
    .aic_6_targ_lt_Ar_Burst(o_aic_6_targ_lt_axi_m_arburst),
    .aic_6_targ_lt_Ar_Cache(o_aic_6_targ_lt_axi_m_arcache),
    .aic_6_targ_lt_Ar_Id(o_aic_6_targ_lt_axi_m_arid),
    .aic_6_targ_lt_Ar_Len(o_aic_6_targ_lt_axi_m_arlen),
    .aic_6_targ_lt_Ar_Lock(o_aic_6_targ_lt_axi_m_arlock),
    .aic_6_targ_lt_Ar_Prot(o_aic_6_targ_lt_axi_m_arprot),
    .aic_6_targ_lt_Ar_Qos(o_aic_6_targ_lt_axi_m_arqos),
    .aic_6_targ_lt_Ar_Ready(i_aic_6_targ_lt_axi_m_arready),
    .aic_6_targ_lt_Ar_Size(o_aic_6_targ_lt_axi_m_arsize),
    .aic_6_targ_lt_Ar_Valid(o_aic_6_targ_lt_axi_m_arvalid),
    .aic_6_targ_lt_Aw_Addr(aic_6_targ_lt_axi_m_awaddr_msb_fixed),
    .aic_6_targ_lt_Aw_Burst(o_aic_6_targ_lt_axi_m_awburst),
    .aic_6_targ_lt_Aw_Cache(o_aic_6_targ_lt_axi_m_awcache),
    .aic_6_targ_lt_Aw_Id(o_aic_6_targ_lt_axi_m_awid),
    .aic_6_targ_lt_Aw_Len(o_aic_6_targ_lt_axi_m_awlen),
    .aic_6_targ_lt_Aw_Lock(o_aic_6_targ_lt_axi_m_awlock),
    .aic_6_targ_lt_Aw_Prot(o_aic_6_targ_lt_axi_m_awprot),
    .aic_6_targ_lt_Aw_Qos(o_aic_6_targ_lt_axi_m_awqos),
    .aic_6_targ_lt_Aw_Ready(i_aic_6_targ_lt_axi_m_awready),
    .aic_6_targ_lt_Aw_Size(o_aic_6_targ_lt_axi_m_awsize),
    .aic_6_targ_lt_Aw_Valid(o_aic_6_targ_lt_axi_m_awvalid),
    .aic_6_targ_lt_B_Id(i_aic_6_targ_lt_axi_m_bid),
    .aic_6_targ_lt_B_Ready(o_aic_6_targ_lt_axi_m_bready),
    .aic_6_targ_lt_B_Resp(i_aic_6_targ_lt_axi_m_bresp),
    .aic_6_targ_lt_B_Valid(i_aic_6_targ_lt_axi_m_bvalid),
    .aic_6_targ_lt_R_Data(i_aic_6_targ_lt_axi_m_rdata),
    .aic_6_targ_lt_R_Id(i_aic_6_targ_lt_axi_m_rid),
    .aic_6_targ_lt_R_Last(i_aic_6_targ_lt_axi_m_rlast),
    .aic_6_targ_lt_R_Ready(o_aic_6_targ_lt_axi_m_rready),
    .aic_6_targ_lt_R_Resp(i_aic_6_targ_lt_axi_m_rresp),
    .aic_6_targ_lt_R_Valid(i_aic_6_targ_lt_axi_m_rvalid),
    .aic_6_targ_lt_W_Data(o_aic_6_targ_lt_axi_m_wdata),
    .aic_6_targ_lt_W_Last(o_aic_6_targ_lt_axi_m_wlast),
    .aic_6_targ_lt_W_Ready(i_aic_6_targ_lt_axi_m_wready),
    .aic_6_targ_lt_W_Strb(o_aic_6_targ_lt_axi_m_wstrb),
    .aic_6_targ_lt_W_Valid(o_aic_6_targ_lt_axi_m_wvalid),
    .aic_6_targ_syscfg_PAddr(o_aic_6_targ_syscfg_apb_m_paddr),
    .aic_6_targ_syscfg_PEnable(o_aic_6_targ_syscfg_apb_m_penable),
    .aic_6_targ_syscfg_PProt(o_aic_6_targ_syscfg_apb_m_pprot),
    .aic_6_targ_syscfg_PRData(i_aic_6_targ_syscfg_apb_m_prdata),
    .aic_6_targ_syscfg_PReady(i_aic_6_targ_syscfg_apb_m_pready),
    .aic_6_targ_syscfg_PSel(o_aic_6_targ_syscfg_apb_m_psel),
    .aic_6_targ_syscfg_PSlvErr(i_aic_6_targ_syscfg_apb_m_pslverr),
    .aic_6_targ_syscfg_PStrb(o_aic_6_targ_syscfg_apb_m_pstrb),
    .aic_6_targ_syscfg_PWData(o_aic_6_targ_syscfg_apb_m_pwdata),
    .aic_6_targ_syscfg_PWrite(o_aic_6_targ_syscfg_apb_m_pwrite),
    .aic_7_aon_clk(i_aic_7_aon_clk),
    .aic_7_aon_rst_n(i_aic_7_aon_rst_n),
    .aic_7_clk(i_aic_7_clk),
    .aic_7_clken(i_aic_7_clken),
    .aic_7_init_ht_rd_Ar_Addr(aic_7_init_ht_axi_s_araddr_msb_fixed),
    .aic_7_init_ht_rd_Ar_Burst(i_aic_7_init_ht_axi_s_arburst),
    .aic_7_init_ht_rd_Ar_Cache(i_aic_7_init_ht_axi_s_arcache),
    .aic_7_init_ht_rd_Ar_Id(i_aic_7_init_ht_axi_s_arid),
    .aic_7_init_ht_rd_Ar_Len(i_aic_7_init_ht_axi_s_arlen),
    .aic_7_init_ht_rd_Ar_Lock(i_aic_7_init_ht_axi_s_arlock),
    .aic_7_init_ht_rd_Ar_Prot(i_aic_7_init_ht_axi_s_arprot),
    .aic_7_init_ht_rd_Ar_Ready(o_aic_7_init_ht_axi_s_arready),
    .aic_7_init_ht_rd_Ar_Size(i_aic_7_init_ht_axi_s_arsize),
    .aic_7_init_ht_rd_Ar_Valid(i_aic_7_init_ht_axi_s_arvalid),
    .aic_7_init_ht_rd_R_Data(o_aic_7_init_ht_axi_s_rdata),
    .aic_7_init_ht_rd_R_Id(o_aic_7_init_ht_axi_s_rid),
    .aic_7_init_ht_rd_R_Last(o_aic_7_init_ht_axi_s_rlast),
    .aic_7_init_ht_rd_R_Ready(i_aic_7_init_ht_axi_s_rready),
    .aic_7_init_ht_rd_R_Resp(o_aic_7_init_ht_axi_s_rresp),
    .aic_7_init_ht_rd_R_Valid(o_aic_7_init_ht_axi_s_rvalid),
    .aic_7_init_ht_wr_Aw_Addr(aic_7_init_ht_axi_s_awaddr_msb_fixed),
    .aic_7_init_ht_wr_Aw_Burst(i_aic_7_init_ht_axi_s_awburst),
    .aic_7_init_ht_wr_Aw_Cache(i_aic_7_init_ht_axi_s_awcache),
    .aic_7_init_ht_wr_Aw_Id(i_aic_7_init_ht_axi_s_awid),
    .aic_7_init_ht_wr_Aw_Len(i_aic_7_init_ht_axi_s_awlen),
    .aic_7_init_ht_wr_Aw_Lock(i_aic_7_init_ht_axi_s_awlock),
    .aic_7_init_ht_wr_Aw_Prot(i_aic_7_init_ht_axi_s_awprot),
    .aic_7_init_ht_wr_Aw_Ready(o_aic_7_init_ht_axi_s_awready),
    .aic_7_init_ht_wr_Aw_Size(i_aic_7_init_ht_axi_s_awsize),
    .aic_7_init_ht_wr_Aw_Valid(i_aic_7_init_ht_axi_s_awvalid),
    .aic_7_init_ht_wr_B_Id(o_aic_7_init_ht_axi_s_bid),
    .aic_7_init_ht_wr_B_Ready(i_aic_7_init_ht_axi_s_bready),
    .aic_7_init_ht_wr_B_Resp(o_aic_7_init_ht_axi_s_bresp),
    .aic_7_init_ht_wr_B_Valid(o_aic_7_init_ht_axi_s_bvalid),
    .aic_7_init_ht_wr_W_Data(i_aic_7_init_ht_axi_s_wdata),
    .aic_7_init_ht_wr_W_Last(i_aic_7_init_ht_axi_s_wlast),
    .aic_7_init_ht_wr_W_Ready(o_aic_7_init_ht_axi_s_wready),
    .aic_7_init_ht_wr_W_Strb(i_aic_7_init_ht_axi_s_wstrb),
    .aic_7_init_ht_wr_W_Valid(i_aic_7_init_ht_axi_s_wvalid),
    .aic_7_init_lt_Ar_Addr(aic_7_init_lt_axi_s_araddr_msb_fixed),
    .aic_7_init_lt_Ar_Burst(i_aic_7_init_lt_axi_s_arburst),
    .aic_7_init_lt_Ar_Cache(i_aic_7_init_lt_axi_s_arcache),
    .aic_7_init_lt_Ar_Id(i_aic_7_init_lt_axi_s_arid),
    .aic_7_init_lt_Ar_Len(i_aic_7_init_lt_axi_s_arlen),
    .aic_7_init_lt_Ar_Lock(i_aic_7_init_lt_axi_s_arlock),
    .aic_7_init_lt_Ar_Prot(i_aic_7_init_lt_axi_s_arprot),
    .aic_7_init_lt_Ar_Qos(i_aic_7_init_lt_axi_s_arqos),
    .aic_7_init_lt_Ar_Ready(o_aic_7_init_lt_axi_s_arready),
    .aic_7_init_lt_Ar_Size(i_aic_7_init_lt_axi_s_arsize),
    .aic_7_init_lt_Ar_Valid(i_aic_7_init_lt_axi_s_arvalid),
    .aic_7_init_lt_Aw_Addr(aic_7_init_lt_axi_s_awaddr_msb_fixed),
    .aic_7_init_lt_Aw_Burst(i_aic_7_init_lt_axi_s_awburst),
    .aic_7_init_lt_Aw_Cache(i_aic_7_init_lt_axi_s_awcache),
    .aic_7_init_lt_Aw_Id(i_aic_7_init_lt_axi_s_awid),
    .aic_7_init_lt_Aw_Len(i_aic_7_init_lt_axi_s_awlen),
    .aic_7_init_lt_Aw_Lock(i_aic_7_init_lt_axi_s_awlock),
    .aic_7_init_lt_Aw_Prot(i_aic_7_init_lt_axi_s_awprot),
    .aic_7_init_lt_Aw_Qos(i_aic_7_init_lt_axi_s_awqos),
    .aic_7_init_lt_Aw_Ready(o_aic_7_init_lt_axi_s_awready),
    .aic_7_init_lt_Aw_Size(i_aic_7_init_lt_axi_s_awsize),
    .aic_7_init_lt_Aw_Valid(i_aic_7_init_lt_axi_s_awvalid),
    .aic_7_init_lt_B_Id(o_aic_7_init_lt_axi_s_bid),
    .aic_7_init_lt_B_Ready(i_aic_7_init_lt_axi_s_bready),
    .aic_7_init_lt_B_Resp(o_aic_7_init_lt_axi_s_bresp),
    .aic_7_init_lt_B_Valid(o_aic_7_init_lt_axi_s_bvalid),
    .aic_7_init_lt_R_Data(o_aic_7_init_lt_axi_s_rdata),
    .aic_7_init_lt_R_Id(o_aic_7_init_lt_axi_s_rid),
    .aic_7_init_lt_R_Last(o_aic_7_init_lt_axi_s_rlast),
    .aic_7_init_lt_R_Ready(i_aic_7_init_lt_axi_s_rready),
    .aic_7_init_lt_R_Resp(o_aic_7_init_lt_axi_s_rresp),
    .aic_7_init_lt_R_Valid(o_aic_7_init_lt_axi_s_rvalid),
    .aic_7_init_lt_W_Data(i_aic_7_init_lt_axi_s_wdata),
    .aic_7_init_lt_W_Last(i_aic_7_init_lt_axi_s_wlast),
    .aic_7_init_lt_W_Ready(o_aic_7_init_lt_axi_s_wready),
    .aic_7_init_lt_W_Strb(i_aic_7_init_lt_axi_s_wstrb),
    .aic_7_init_lt_W_Valid(i_aic_7_init_lt_axi_s_wvalid),
    .aic_7_pwr_Idle(o_aic_7_pwr_idle_val),
    .aic_7_pwr_IdleAck(o_aic_7_pwr_idle_ack),
    .aic_7_pwr_IdleReq(i_aic_7_pwr_idle_req),
    .aic_7_rst_n(i_aic_7_rst_n),
    .aic_7_targ_lt_Ar_Addr(aic_7_targ_lt_axi_m_araddr_msb_fixed),
    .aic_7_targ_lt_Ar_Burst(o_aic_7_targ_lt_axi_m_arburst),
    .aic_7_targ_lt_Ar_Cache(o_aic_7_targ_lt_axi_m_arcache),
    .aic_7_targ_lt_Ar_Id(o_aic_7_targ_lt_axi_m_arid),
    .aic_7_targ_lt_Ar_Len(o_aic_7_targ_lt_axi_m_arlen),
    .aic_7_targ_lt_Ar_Lock(o_aic_7_targ_lt_axi_m_arlock),
    .aic_7_targ_lt_Ar_Prot(o_aic_7_targ_lt_axi_m_arprot),
    .aic_7_targ_lt_Ar_Qos(o_aic_7_targ_lt_axi_m_arqos),
    .aic_7_targ_lt_Ar_Ready(i_aic_7_targ_lt_axi_m_arready),
    .aic_7_targ_lt_Ar_Size(o_aic_7_targ_lt_axi_m_arsize),
    .aic_7_targ_lt_Ar_Valid(o_aic_7_targ_lt_axi_m_arvalid),
    .aic_7_targ_lt_Aw_Addr(aic_7_targ_lt_axi_m_awaddr_msb_fixed),
    .aic_7_targ_lt_Aw_Burst(o_aic_7_targ_lt_axi_m_awburst),
    .aic_7_targ_lt_Aw_Cache(o_aic_7_targ_lt_axi_m_awcache),
    .aic_7_targ_lt_Aw_Id(o_aic_7_targ_lt_axi_m_awid),
    .aic_7_targ_lt_Aw_Len(o_aic_7_targ_lt_axi_m_awlen),
    .aic_7_targ_lt_Aw_Lock(o_aic_7_targ_lt_axi_m_awlock),
    .aic_7_targ_lt_Aw_Prot(o_aic_7_targ_lt_axi_m_awprot),
    .aic_7_targ_lt_Aw_Qos(o_aic_7_targ_lt_axi_m_awqos),
    .aic_7_targ_lt_Aw_Ready(i_aic_7_targ_lt_axi_m_awready),
    .aic_7_targ_lt_Aw_Size(o_aic_7_targ_lt_axi_m_awsize),
    .aic_7_targ_lt_Aw_Valid(o_aic_7_targ_lt_axi_m_awvalid),
    .aic_7_targ_lt_B_Id(i_aic_7_targ_lt_axi_m_bid),
    .aic_7_targ_lt_B_Ready(o_aic_7_targ_lt_axi_m_bready),
    .aic_7_targ_lt_B_Resp(i_aic_7_targ_lt_axi_m_bresp),
    .aic_7_targ_lt_B_Valid(i_aic_7_targ_lt_axi_m_bvalid),
    .aic_7_targ_lt_R_Data(i_aic_7_targ_lt_axi_m_rdata),
    .aic_7_targ_lt_R_Id(i_aic_7_targ_lt_axi_m_rid),
    .aic_7_targ_lt_R_Last(i_aic_7_targ_lt_axi_m_rlast),
    .aic_7_targ_lt_R_Ready(o_aic_7_targ_lt_axi_m_rready),
    .aic_7_targ_lt_R_Resp(i_aic_7_targ_lt_axi_m_rresp),
    .aic_7_targ_lt_R_Valid(i_aic_7_targ_lt_axi_m_rvalid),
    .aic_7_targ_lt_W_Data(o_aic_7_targ_lt_axi_m_wdata),
    .aic_7_targ_lt_W_Last(o_aic_7_targ_lt_axi_m_wlast),
    .aic_7_targ_lt_W_Ready(i_aic_7_targ_lt_axi_m_wready),
    .aic_7_targ_lt_W_Strb(o_aic_7_targ_lt_axi_m_wstrb),
    .aic_7_targ_lt_W_Valid(o_aic_7_targ_lt_axi_m_wvalid),
    .aic_7_targ_syscfg_PAddr(o_aic_7_targ_syscfg_apb_m_paddr),
    .aic_7_targ_syscfg_PEnable(o_aic_7_targ_syscfg_apb_m_penable),
    .aic_7_targ_syscfg_PProt(o_aic_7_targ_syscfg_apb_m_pprot),
    .aic_7_targ_syscfg_PRData(i_aic_7_targ_syscfg_apb_m_prdata),
    .aic_7_targ_syscfg_PReady(i_aic_7_targ_syscfg_apb_m_pready),
    .aic_7_targ_syscfg_PSel(o_aic_7_targ_syscfg_apb_m_psel),
    .aic_7_targ_syscfg_PSlvErr(i_aic_7_targ_syscfg_apb_m_pslverr),
    .aic_7_targ_syscfg_PStrb(o_aic_7_targ_syscfg_apb_m_pstrb),
    .aic_7_targ_syscfg_PWData(o_aic_7_targ_syscfg_apb_m_pwdata),
    .aic_7_targ_syscfg_PWrite(o_aic_7_targ_syscfg_apb_m_pwrite),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Data(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Head(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Data(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Head(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Data(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Head(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Data(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Head(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Data(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Head(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Data(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Head(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Data(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Head(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Data(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Head(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Data(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Head(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Data(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Head(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Data(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Head(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Rdy(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Tail(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail),
    .dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_Vld(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Data(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Head(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Data(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Head(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Rdy(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Tail(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail),
    .dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_Vld(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Data(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Head(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Rdy(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Tail(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail),
    .dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_Vld(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Data(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Head(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Rdy(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Tail(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail),
    .dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_Vld(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Data(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Head(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Rdy(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Tail(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail),
    .dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_Vld(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Data(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Head(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Rdy(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Tail(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_Vld(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Data(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Head(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Data(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Head(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Rdy(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Tail(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_Vld(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Data(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Head(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Data(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Head(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Rdy(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Tail(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_Vld(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Data(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Head(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Data(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Head(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Rdy(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Tail(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_Vld(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Data(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Head(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Data(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Head(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Rdy(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Tail(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_Vld(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Data(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Head(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Data(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Head(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Rdy(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Tail(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_Vld(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Data(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Head(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Data(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Head(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Rdy(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Tail(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_Vld(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Data(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Head(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Data(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Head(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Rdy(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Tail(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_Vld(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Data(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Head(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Data(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Head(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Rdy(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Tail(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_Vld(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Data(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Head(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Data(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Head(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Rdy(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Tail(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_Vld(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Data(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Head(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Data(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Head(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Rdy(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Tail(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail),
    .dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_Vld(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Data(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Head(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Data(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Head(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Rdy(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Tail(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail),
    .dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_Vld(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Data(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Head(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Rdy(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Tail(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail),
    .dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_Vld(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Data(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Head(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Rdy(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Tail(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail),
    .dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_Vld(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Data(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Head(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Rdy(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Tail(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail),
    .dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_Vld(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld),
    .l2_4_aon_clk(i_l2_4_aon_clk),
    .l2_4_aon_rst_n(i_l2_4_aon_rst_n),
    .l2_4_clk(i_l2_4_clk),
    .l2_4_clken(i_l2_4_clken),
    .l2_4_pwr_Idle(o_l2_4_pwr_idle_val),
    .l2_4_pwr_IdleAck(o_l2_4_pwr_idle_ack),
    .l2_4_pwr_IdleReq(i_l2_4_pwr_idle_req),
    .l2_4_rst_n(i_l2_4_rst_n),
    .l2_4_targ_ht_rd_Ar_Addr(l2_4_targ_ht_axi_m_araddr_msb_fixed),
    .l2_4_targ_ht_rd_Ar_Burst(o_l2_4_targ_ht_axi_m_arburst),
    .l2_4_targ_ht_rd_Ar_Cache(o_l2_4_targ_ht_axi_m_arcache),
    .l2_4_targ_ht_rd_Ar_Id(o_l2_4_targ_ht_axi_m_arid),
    .l2_4_targ_ht_rd_Ar_Len(o_l2_4_targ_ht_axi_m_arlen),
    .l2_4_targ_ht_rd_Ar_Lock(o_l2_4_targ_ht_axi_m_arlock),
    .l2_4_targ_ht_rd_Ar_Prot(o_l2_4_targ_ht_axi_m_arprot),
    .l2_4_targ_ht_rd_Ar_Ready(i_l2_4_targ_ht_axi_m_arready),
    .l2_4_targ_ht_rd_Ar_Size(o_l2_4_targ_ht_axi_m_arsize),
    .l2_4_targ_ht_rd_Ar_Valid(o_l2_4_targ_ht_axi_m_arvalid),
    .l2_4_targ_ht_rd_R_Data(i_l2_4_targ_ht_axi_m_rdata),
    .l2_4_targ_ht_rd_R_Id(i_l2_4_targ_ht_axi_m_rid),
    .l2_4_targ_ht_rd_R_Last(i_l2_4_targ_ht_axi_m_rlast),
    .l2_4_targ_ht_rd_R_Ready(o_l2_4_targ_ht_axi_m_rready),
    .l2_4_targ_ht_rd_R_Resp(i_l2_4_targ_ht_axi_m_rresp),
    .l2_4_targ_ht_rd_R_Valid(i_l2_4_targ_ht_axi_m_rvalid),
    .l2_4_targ_ht_wr_Aw_Addr(l2_4_targ_ht_axi_m_awaddr_msb_fixed),
    .l2_4_targ_ht_wr_Aw_Burst(o_l2_4_targ_ht_axi_m_awburst),
    .l2_4_targ_ht_wr_Aw_Cache(o_l2_4_targ_ht_axi_m_awcache),
    .l2_4_targ_ht_wr_Aw_Id(o_l2_4_targ_ht_axi_m_awid),
    .l2_4_targ_ht_wr_Aw_Len(o_l2_4_targ_ht_axi_m_awlen),
    .l2_4_targ_ht_wr_Aw_Lock(o_l2_4_targ_ht_axi_m_awlock),
    .l2_4_targ_ht_wr_Aw_Prot(o_l2_4_targ_ht_axi_m_awprot),
    .l2_4_targ_ht_wr_Aw_Ready(i_l2_4_targ_ht_axi_m_awready),
    .l2_4_targ_ht_wr_Aw_Size(o_l2_4_targ_ht_axi_m_awsize),
    .l2_4_targ_ht_wr_Aw_Valid(o_l2_4_targ_ht_axi_m_awvalid),
    .l2_4_targ_ht_wr_B_Id(i_l2_4_targ_ht_axi_m_bid),
    .l2_4_targ_ht_wr_B_Ready(o_l2_4_targ_ht_axi_m_bready),
    .l2_4_targ_ht_wr_B_Resp(i_l2_4_targ_ht_axi_m_bresp),
    .l2_4_targ_ht_wr_B_Valid(i_l2_4_targ_ht_axi_m_bvalid),
    .l2_4_targ_ht_wr_W_Data(o_l2_4_targ_ht_axi_m_wdata),
    .l2_4_targ_ht_wr_W_Last(o_l2_4_targ_ht_axi_m_wlast),
    .l2_4_targ_ht_wr_W_Ready(i_l2_4_targ_ht_axi_m_wready),
    .l2_4_targ_ht_wr_W_Strb(o_l2_4_targ_ht_axi_m_wstrb),
    .l2_4_targ_ht_wr_W_Valid(o_l2_4_targ_ht_axi_m_wvalid),
    .l2_4_targ_syscfg_PAddr(o_l2_4_targ_syscfg_apb_m_paddr),
    .l2_4_targ_syscfg_PEnable(o_l2_4_targ_syscfg_apb_m_penable),
    .l2_4_targ_syscfg_PProt(o_l2_4_targ_syscfg_apb_m_pprot),
    .l2_4_targ_syscfg_PRData(i_l2_4_targ_syscfg_apb_m_prdata),
    .l2_4_targ_syscfg_PReady(i_l2_4_targ_syscfg_apb_m_pready),
    .l2_4_targ_syscfg_PSel(o_l2_4_targ_syscfg_apb_m_psel),
    .l2_4_targ_syscfg_PSlvErr(i_l2_4_targ_syscfg_apb_m_pslverr),
    .l2_4_targ_syscfg_PStrb(o_l2_4_targ_syscfg_apb_m_pstrb),
    .l2_4_targ_syscfg_PWData(o_l2_4_targ_syscfg_apb_m_pwdata),
    .l2_4_targ_syscfg_PWrite(o_l2_4_targ_syscfg_apb_m_pwrite),
    .l2_5_aon_clk(i_l2_5_aon_clk),
    .l2_5_aon_rst_n(i_l2_5_aon_rst_n),
    .l2_5_clk(i_l2_5_clk),
    .l2_5_clken(i_l2_5_clken),
    .l2_5_pwr_Idle(o_l2_5_pwr_idle_val),
    .l2_5_pwr_IdleAck(o_l2_5_pwr_idle_ack),
    .l2_5_pwr_IdleReq(i_l2_5_pwr_idle_req),
    .l2_5_rst_n(i_l2_5_rst_n),
    .l2_5_targ_ht_rd_Ar_Addr(l2_5_targ_ht_axi_m_araddr_msb_fixed),
    .l2_5_targ_ht_rd_Ar_Burst(o_l2_5_targ_ht_axi_m_arburst),
    .l2_5_targ_ht_rd_Ar_Cache(o_l2_5_targ_ht_axi_m_arcache),
    .l2_5_targ_ht_rd_Ar_Id(o_l2_5_targ_ht_axi_m_arid),
    .l2_5_targ_ht_rd_Ar_Len(o_l2_5_targ_ht_axi_m_arlen),
    .l2_5_targ_ht_rd_Ar_Lock(o_l2_5_targ_ht_axi_m_arlock),
    .l2_5_targ_ht_rd_Ar_Prot(o_l2_5_targ_ht_axi_m_arprot),
    .l2_5_targ_ht_rd_Ar_Ready(i_l2_5_targ_ht_axi_m_arready),
    .l2_5_targ_ht_rd_Ar_Size(o_l2_5_targ_ht_axi_m_arsize),
    .l2_5_targ_ht_rd_Ar_Valid(o_l2_5_targ_ht_axi_m_arvalid),
    .l2_5_targ_ht_rd_R_Data(i_l2_5_targ_ht_axi_m_rdata),
    .l2_5_targ_ht_rd_R_Id(i_l2_5_targ_ht_axi_m_rid),
    .l2_5_targ_ht_rd_R_Last(i_l2_5_targ_ht_axi_m_rlast),
    .l2_5_targ_ht_rd_R_Ready(o_l2_5_targ_ht_axi_m_rready),
    .l2_5_targ_ht_rd_R_Resp(i_l2_5_targ_ht_axi_m_rresp),
    .l2_5_targ_ht_rd_R_Valid(i_l2_5_targ_ht_axi_m_rvalid),
    .l2_5_targ_ht_wr_Aw_Addr(l2_5_targ_ht_axi_m_awaddr_msb_fixed),
    .l2_5_targ_ht_wr_Aw_Burst(o_l2_5_targ_ht_axi_m_awburst),
    .l2_5_targ_ht_wr_Aw_Cache(o_l2_5_targ_ht_axi_m_awcache),
    .l2_5_targ_ht_wr_Aw_Id(o_l2_5_targ_ht_axi_m_awid),
    .l2_5_targ_ht_wr_Aw_Len(o_l2_5_targ_ht_axi_m_awlen),
    .l2_5_targ_ht_wr_Aw_Lock(o_l2_5_targ_ht_axi_m_awlock),
    .l2_5_targ_ht_wr_Aw_Prot(o_l2_5_targ_ht_axi_m_awprot),
    .l2_5_targ_ht_wr_Aw_Ready(i_l2_5_targ_ht_axi_m_awready),
    .l2_5_targ_ht_wr_Aw_Size(o_l2_5_targ_ht_axi_m_awsize),
    .l2_5_targ_ht_wr_Aw_Valid(o_l2_5_targ_ht_axi_m_awvalid),
    .l2_5_targ_ht_wr_B_Id(i_l2_5_targ_ht_axi_m_bid),
    .l2_5_targ_ht_wr_B_Ready(o_l2_5_targ_ht_axi_m_bready),
    .l2_5_targ_ht_wr_B_Resp(i_l2_5_targ_ht_axi_m_bresp),
    .l2_5_targ_ht_wr_B_Valid(i_l2_5_targ_ht_axi_m_bvalid),
    .l2_5_targ_ht_wr_W_Data(o_l2_5_targ_ht_axi_m_wdata),
    .l2_5_targ_ht_wr_W_Last(o_l2_5_targ_ht_axi_m_wlast),
    .l2_5_targ_ht_wr_W_Ready(i_l2_5_targ_ht_axi_m_wready),
    .l2_5_targ_ht_wr_W_Strb(o_l2_5_targ_ht_axi_m_wstrb),
    .l2_5_targ_ht_wr_W_Valid(o_l2_5_targ_ht_axi_m_wvalid),
    .l2_5_targ_syscfg_PAddr(o_l2_5_targ_syscfg_apb_m_paddr),
    .l2_5_targ_syscfg_PEnable(o_l2_5_targ_syscfg_apb_m_penable),
    .l2_5_targ_syscfg_PProt(o_l2_5_targ_syscfg_apb_m_pprot),
    .l2_5_targ_syscfg_PRData(i_l2_5_targ_syscfg_apb_m_prdata),
    .l2_5_targ_syscfg_PReady(i_l2_5_targ_syscfg_apb_m_pready),
    .l2_5_targ_syscfg_PSel(o_l2_5_targ_syscfg_apb_m_psel),
    .l2_5_targ_syscfg_PSlvErr(i_l2_5_targ_syscfg_apb_m_pslverr),
    .l2_5_targ_syscfg_PStrb(o_l2_5_targ_syscfg_apb_m_pstrb),
    .l2_5_targ_syscfg_PWData(o_l2_5_targ_syscfg_apb_m_pwdata),
    .l2_5_targ_syscfg_PWrite(o_l2_5_targ_syscfg_apb_m_pwrite),
    .l2_6_aon_clk(i_l2_6_aon_clk),
    .l2_6_aon_rst_n(i_l2_6_aon_rst_n),
    .l2_6_clk(i_l2_6_clk),
    .l2_6_clken(i_l2_6_clken),
    .l2_6_pwr_Idle(o_l2_6_pwr_idle_val),
    .l2_6_pwr_IdleAck(o_l2_6_pwr_idle_ack),
    .l2_6_pwr_IdleReq(i_l2_6_pwr_idle_req),
    .l2_6_rst_n(i_l2_6_rst_n),
    .l2_6_targ_ht_rd_Ar_Addr(l2_6_targ_ht_axi_m_araddr_msb_fixed),
    .l2_6_targ_ht_rd_Ar_Burst(o_l2_6_targ_ht_axi_m_arburst),
    .l2_6_targ_ht_rd_Ar_Cache(o_l2_6_targ_ht_axi_m_arcache),
    .l2_6_targ_ht_rd_Ar_Id(o_l2_6_targ_ht_axi_m_arid),
    .l2_6_targ_ht_rd_Ar_Len(o_l2_6_targ_ht_axi_m_arlen),
    .l2_6_targ_ht_rd_Ar_Lock(o_l2_6_targ_ht_axi_m_arlock),
    .l2_6_targ_ht_rd_Ar_Prot(o_l2_6_targ_ht_axi_m_arprot),
    .l2_6_targ_ht_rd_Ar_Ready(i_l2_6_targ_ht_axi_m_arready),
    .l2_6_targ_ht_rd_Ar_Size(o_l2_6_targ_ht_axi_m_arsize),
    .l2_6_targ_ht_rd_Ar_Valid(o_l2_6_targ_ht_axi_m_arvalid),
    .l2_6_targ_ht_rd_R_Data(i_l2_6_targ_ht_axi_m_rdata),
    .l2_6_targ_ht_rd_R_Id(i_l2_6_targ_ht_axi_m_rid),
    .l2_6_targ_ht_rd_R_Last(i_l2_6_targ_ht_axi_m_rlast),
    .l2_6_targ_ht_rd_R_Ready(o_l2_6_targ_ht_axi_m_rready),
    .l2_6_targ_ht_rd_R_Resp(i_l2_6_targ_ht_axi_m_rresp),
    .l2_6_targ_ht_rd_R_Valid(i_l2_6_targ_ht_axi_m_rvalid),
    .l2_6_targ_ht_wr_Aw_Addr(l2_6_targ_ht_axi_m_awaddr_msb_fixed),
    .l2_6_targ_ht_wr_Aw_Burst(o_l2_6_targ_ht_axi_m_awburst),
    .l2_6_targ_ht_wr_Aw_Cache(o_l2_6_targ_ht_axi_m_awcache),
    .l2_6_targ_ht_wr_Aw_Id(o_l2_6_targ_ht_axi_m_awid),
    .l2_6_targ_ht_wr_Aw_Len(o_l2_6_targ_ht_axi_m_awlen),
    .l2_6_targ_ht_wr_Aw_Lock(o_l2_6_targ_ht_axi_m_awlock),
    .l2_6_targ_ht_wr_Aw_Prot(o_l2_6_targ_ht_axi_m_awprot),
    .l2_6_targ_ht_wr_Aw_Ready(i_l2_6_targ_ht_axi_m_awready),
    .l2_6_targ_ht_wr_Aw_Size(o_l2_6_targ_ht_axi_m_awsize),
    .l2_6_targ_ht_wr_Aw_Valid(o_l2_6_targ_ht_axi_m_awvalid),
    .l2_6_targ_ht_wr_B_Id(i_l2_6_targ_ht_axi_m_bid),
    .l2_6_targ_ht_wr_B_Ready(o_l2_6_targ_ht_axi_m_bready),
    .l2_6_targ_ht_wr_B_Resp(i_l2_6_targ_ht_axi_m_bresp),
    .l2_6_targ_ht_wr_B_Valid(i_l2_6_targ_ht_axi_m_bvalid),
    .l2_6_targ_ht_wr_W_Data(o_l2_6_targ_ht_axi_m_wdata),
    .l2_6_targ_ht_wr_W_Last(o_l2_6_targ_ht_axi_m_wlast),
    .l2_6_targ_ht_wr_W_Ready(i_l2_6_targ_ht_axi_m_wready),
    .l2_6_targ_ht_wr_W_Strb(o_l2_6_targ_ht_axi_m_wstrb),
    .l2_6_targ_ht_wr_W_Valid(o_l2_6_targ_ht_axi_m_wvalid),
    .l2_6_targ_syscfg_PAddr(o_l2_6_targ_syscfg_apb_m_paddr),
    .l2_6_targ_syscfg_PEnable(o_l2_6_targ_syscfg_apb_m_penable),
    .l2_6_targ_syscfg_PProt(o_l2_6_targ_syscfg_apb_m_pprot),
    .l2_6_targ_syscfg_PRData(i_l2_6_targ_syscfg_apb_m_prdata),
    .l2_6_targ_syscfg_PReady(i_l2_6_targ_syscfg_apb_m_pready),
    .l2_6_targ_syscfg_PSel(o_l2_6_targ_syscfg_apb_m_psel),
    .l2_6_targ_syscfg_PSlvErr(i_l2_6_targ_syscfg_apb_m_pslverr),
    .l2_6_targ_syscfg_PStrb(o_l2_6_targ_syscfg_apb_m_pstrb),
    .l2_6_targ_syscfg_PWData(o_l2_6_targ_syscfg_apb_m_pwdata),
    .l2_6_targ_syscfg_PWrite(o_l2_6_targ_syscfg_apb_m_pwrite),
    .l2_7_aon_clk(i_l2_7_aon_clk),
    .l2_7_aon_rst_n(i_l2_7_aon_rst_n),
    .l2_7_clk(i_l2_7_clk),
    .l2_7_clken(i_l2_7_clken),
    .l2_7_pwr_Idle(o_l2_7_pwr_idle_val),
    .l2_7_pwr_IdleAck(o_l2_7_pwr_idle_ack),
    .l2_7_pwr_IdleReq(i_l2_7_pwr_idle_req),
    .l2_7_rst_n(i_l2_7_rst_n),
    .l2_7_targ_ht_rd_Ar_Addr(l2_7_targ_ht_axi_m_araddr_msb_fixed),
    .l2_7_targ_ht_rd_Ar_Burst(o_l2_7_targ_ht_axi_m_arburst),
    .l2_7_targ_ht_rd_Ar_Cache(o_l2_7_targ_ht_axi_m_arcache),
    .l2_7_targ_ht_rd_Ar_Id(o_l2_7_targ_ht_axi_m_arid),
    .l2_7_targ_ht_rd_Ar_Len(o_l2_7_targ_ht_axi_m_arlen),
    .l2_7_targ_ht_rd_Ar_Lock(o_l2_7_targ_ht_axi_m_arlock),
    .l2_7_targ_ht_rd_Ar_Prot(o_l2_7_targ_ht_axi_m_arprot),
    .l2_7_targ_ht_rd_Ar_Ready(i_l2_7_targ_ht_axi_m_arready),
    .l2_7_targ_ht_rd_Ar_Size(o_l2_7_targ_ht_axi_m_arsize),
    .l2_7_targ_ht_rd_Ar_Valid(o_l2_7_targ_ht_axi_m_arvalid),
    .l2_7_targ_ht_rd_R_Data(i_l2_7_targ_ht_axi_m_rdata),
    .l2_7_targ_ht_rd_R_Id(i_l2_7_targ_ht_axi_m_rid),
    .l2_7_targ_ht_rd_R_Last(i_l2_7_targ_ht_axi_m_rlast),
    .l2_7_targ_ht_rd_R_Ready(o_l2_7_targ_ht_axi_m_rready),
    .l2_7_targ_ht_rd_R_Resp(i_l2_7_targ_ht_axi_m_rresp),
    .l2_7_targ_ht_rd_R_Valid(i_l2_7_targ_ht_axi_m_rvalid),
    .l2_7_targ_ht_wr_Aw_Addr(l2_7_targ_ht_axi_m_awaddr_msb_fixed),
    .l2_7_targ_ht_wr_Aw_Burst(o_l2_7_targ_ht_axi_m_awburst),
    .l2_7_targ_ht_wr_Aw_Cache(o_l2_7_targ_ht_axi_m_awcache),
    .l2_7_targ_ht_wr_Aw_Id(o_l2_7_targ_ht_axi_m_awid),
    .l2_7_targ_ht_wr_Aw_Len(o_l2_7_targ_ht_axi_m_awlen),
    .l2_7_targ_ht_wr_Aw_Lock(o_l2_7_targ_ht_axi_m_awlock),
    .l2_7_targ_ht_wr_Aw_Prot(o_l2_7_targ_ht_axi_m_awprot),
    .l2_7_targ_ht_wr_Aw_Ready(i_l2_7_targ_ht_axi_m_awready),
    .l2_7_targ_ht_wr_Aw_Size(o_l2_7_targ_ht_axi_m_awsize),
    .l2_7_targ_ht_wr_Aw_Valid(o_l2_7_targ_ht_axi_m_awvalid),
    .l2_7_targ_ht_wr_B_Id(i_l2_7_targ_ht_axi_m_bid),
    .l2_7_targ_ht_wr_B_Ready(o_l2_7_targ_ht_axi_m_bready),
    .l2_7_targ_ht_wr_B_Resp(i_l2_7_targ_ht_axi_m_bresp),
    .l2_7_targ_ht_wr_B_Valid(i_l2_7_targ_ht_axi_m_bvalid),
    .l2_7_targ_ht_wr_W_Data(o_l2_7_targ_ht_axi_m_wdata),
    .l2_7_targ_ht_wr_W_Last(o_l2_7_targ_ht_axi_m_wlast),
    .l2_7_targ_ht_wr_W_Ready(i_l2_7_targ_ht_axi_m_wready),
    .l2_7_targ_ht_wr_W_Strb(o_l2_7_targ_ht_axi_m_wstrb),
    .l2_7_targ_ht_wr_W_Valid(o_l2_7_targ_ht_axi_m_wvalid),
    .l2_7_targ_syscfg_PAddr(o_l2_7_targ_syscfg_apb_m_paddr),
    .l2_7_targ_syscfg_PEnable(o_l2_7_targ_syscfg_apb_m_penable),
    .l2_7_targ_syscfg_PProt(o_l2_7_targ_syscfg_apb_m_pprot),
    .l2_7_targ_syscfg_PRData(i_l2_7_targ_syscfg_apb_m_prdata),
    .l2_7_targ_syscfg_PReady(i_l2_7_targ_syscfg_apb_m_pready),
    .l2_7_targ_syscfg_PSel(o_l2_7_targ_syscfg_apb_m_psel),
    .l2_7_targ_syscfg_PSlvErr(i_l2_7_targ_syscfg_apb_m_pslverr),
    .l2_7_targ_syscfg_PStrb(o_l2_7_targ_syscfg_apb_m_pstrb),
    .l2_7_targ_syscfg_PWData(o_l2_7_targ_syscfg_apb_m_pwdata),
    .l2_7_targ_syscfg_PWrite(o_l2_7_targ_syscfg_apb_m_pwrite),
    .l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .noc_clk(i_noc_clk),
    .noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
);

endmodule
