const phy_init_data_t ddrctl_init_details[string][] = '{
"A" : '{
'{step_type:POLL,reg_addr : 32'h10ff8,value : 32'd0},
'{step_type:POLL,reg_addr : 32'h10ffc,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h10b84,value : 32'd1},
'{step_type:REG_WRITE,reg_addr : 32'h10000,value : 32'd50855944},
'{step_type:REG_WRITE,reg_addr : 32'h10010,value : 32'd273},
'{step_type:REG_WRITE,reg_addr : 32'h10100,value : 32'd1},
'{step_type:REG_WRITE,reg_addr : 32'h10104,value : 32'd15},
'{step_type:REG_WRITE,reg_addr : 32'h10108,value : 32'd15},
'{step_type:REG_WRITE,reg_addr : 32'h10118,value : 32'd1},
'{step_type:REG_WRITE,reg_addr : 32'h10180,value : 32'd1},
'{step_type:REG_WRITE,reg_addr : 32'h10184,value : 32'd2},
'{step_type:REG_WRITE,reg_addr : 32'h1018c,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h10200,value : 32'd4},
'{step_type:REG_WRITE,reg_addr : 32'h10220,value : 32'd520093953},
'{step_type:REG_WRITE,reg_addr : 32'h10224,value : 32'd14},
'{step_type:REG_WRITE,reg_addr : 32'h10300,value : 32'd6160478},
'{step_type:REG_WRITE,reg_addr : 32'h10308,value : 32'd1},
'{step_type:REG_WRITE,reg_addr : 32'h10380,value : 32'd671202832},
'{step_type:REG_WRITE,reg_addr : 32'h10390,value : 32'd138151952},
'{step_type:REG_WRITE,reg_addr : 32'h10394,value : 32'd7453},
'{step_type:REG_WRITE,reg_addr : 32'h10400,value : 32'd2147483728},
'{step_type:REG_WRITE,reg_addr : 32'h10500,value : 32'd1048849},
'{step_type:REG_WRITE,reg_addr : 32'h10508,value : 32'd1610645504},
'{step_type:REG_WRITE,reg_addr : 32'h10510,value : 32'd65541},
'{step_type:REG_WRITE,reg_addr : 32'h10518,value : 32'd2097152001},
'{step_type:REG_WRITE,reg_addr : 32'h10600,value : 32'd3829349504},
'{step_type:REG_WRITE,reg_addr : 32'h10604,value : 32'd8114},
'{step_type:REG_WRITE,reg_addr : 32'h10648,value : 32'd16778112},
'{step_type:REG_WRITE,reg_addr : 32'h1064c,value : 32'd146926},
'{step_type:REG_WRITE,reg_addr : 32'h10658,value : 32'd4078640039},
'{step_type:REG_WRITE,reg_addr : 32'h10660,value : 32'd254},
'{step_type:REG_WRITE,reg_addr : 32'h10c90,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h10cb0,value : 32'd17},
'{step_type:REG_WRITE,reg_addr : 32'h10d00,value : 32'd1073938436},
'{step_type:REG_WRITE,reg_addr : 32'h10f00,value : 32'd2149081472},
'{step_type:REG_WRITE,reg_addr : 32'h20000,value : 32'd16},
'{step_type:REG_WRITE,reg_addr : 32'h20004,value : 32'd6316032},
'{step_type:REG_WRITE,reg_addr : 32'h20008,value : 32'd16384},
'{step_type:REG_WRITE,reg_addr : 32'h20094,value : 32'd16780812},
'{step_type:REG_WRITE,reg_addr : 32'h20098,value : 32'd97124609},
'{step_type:REG_WRITE,reg_addr : 32'h2009c,value : 32'd16779779},
'{step_type:REG_WRITE,reg_addr : 32'h200a0,value : 32'd44631896},
'{step_type:REG_WRITE,reg_addr : 32'h200e0,value : 32'd268458000},
'{step_type:REG_WRITE,reg_addr : 32'h200f0,value : 32'd1303953134},
'{step_type:REG_WRITE,reg_addr : 32'h200f8,value : 32'd1352986425},
'{step_type:REG_WRITE,reg_addr : 32'h0     ,value : 32'd688928290},
'{step_type:REG_WRITE,reg_addr : 32'h4     ,value : 32'd84281392},
'{step_type:REG_WRITE,reg_addr : 32'h8     ,value : 32'd152179225},
'{step_type:REG_WRITE,reg_addr : 32'hc     ,value : 32'd795184},
'{step_type:REG_WRITE,reg_addr : 32'h10    ,value : 32'd251921423},
'{step_type:REG_WRITE,reg_addr : 32'h14    ,value : 32'd33819657},
'{step_type:REG_WRITE,reg_addr : 32'h18    ,value : 32'd8},
'{step_type:REG_WRITE,reg_addr : 32'h1c    ,value : 32'd3},
'{step_type:REG_WRITE,reg_addr : 32'h24    ,value : 32'd132114},
'{step_type:REG_WRITE,reg_addr : 32'h30    ,value : 32'd196608},
'{step_type:REG_WRITE,reg_addr : 32'h34    ,value : 32'd202375170},
'{step_type:REG_WRITE,reg_addr : 32'h38    ,value : 32'd3735862},
'{step_type:REG_WRITE,reg_addr : 32'h44    ,value : 32'd7864400},
'{step_type:REG_WRITE,reg_addr : 32'h5c    ,value : 32'd10289161},
'{step_type:REG_WRITE,reg_addr : 32'h60    ,value : 32'd1054478},
'{step_type:REG_WRITE,reg_addr : 32'h64    ,value : 32'd10502},
'{step_type:REG_WRITE,reg_addr : 32'h78    ,value : 32'd1709081},
'{step_type:REG_WRITE,reg_addr : 32'h500   ,value : 32'd1296},
'{step_type:REG_WRITE,reg_addr : 32'h504   ,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h508   ,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h50c   ,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h580   ,value : 32'd54198815},
'{step_type:REG_WRITE,reg_addr : 32'h584   ,value : 32'd525059},
'{step_type:REG_WRITE,reg_addr : 32'h588   ,value : 32'd1587999},
'{step_type:REG_WRITE,reg_addr : 32'h590   ,value : 32'd470549521},
'{step_type:REG_WRITE,reg_addr : 32'h594   ,value : 32'd68157455},
'{step_type:REG_WRITE,reg_addr : 32'h598   ,value : 32'd279},
'{step_type:REG_WRITE,reg_addr : 32'h5a0   ,value : 32'd197379},
'{step_type:REG_WRITE,reg_addr : 32'h5a4   ,value : 32'd770},
'{step_type:REG_WRITE,reg_addr : 32'h5a8   ,value : 32'd26214415},
'{step_type:REG_WRITE,reg_addr : 32'h5ac   ,value : 32'd851983},
'{step_type:REG_WRITE,reg_addr : 32'h5b4   ,value : 32'd1073741838},
'{step_type:REG_WRITE,reg_addr : 32'h5b8   ,value : 32'd327},
'{step_type:REG_WRITE,reg_addr : 32'h600   ,value : 32'd3224833076},
'{step_type:REG_WRITE,reg_addr : 32'h604   ,value : 32'd19923248},
'{step_type:REG_WRITE,reg_addr : 32'h608   ,value : 32'd105381888},
'{step_type:REG_WRITE,reg_addr : 32'h60c   ,value : 32'd16777216},
'{step_type:REG_WRITE,reg_addr : 32'h650   ,value : 32'd208},
'{step_type:REG_WRITE,reg_addr : 32'h800   ,value : 32'd1574103},
'{step_type:REG_WRITE,reg_addr : 32'h804   ,value : 32'd41943138},
'{step_type:REG_WRITE,reg_addr : 32'ha80   ,value : 32'd10468},
'{step_type:REG_WRITE,reg_addr : 32'hb00   ,value : 32'd2383496020},
'{step_type:REG_WRITE,reg_addr : 32'hb04   ,value : 32'd270798858},
'{step_type:REG_WRITE,reg_addr : 32'hb08   ,value : 32'd1331},
'{step_type:REG_WRITE,reg_addr : 32'hb80   ,value : 32'd64356352},
'{step_type:REG_WRITE,reg_addr : 32'hc88   ,value : 32'd251658283},
'{step_type:REG_WRITE,reg_addr : 32'hd00   ,value : 32'd1},
'{step_type:REG_WRITE,reg_addr : 32'hd04   ,value : 32'd2823},
'{step_type:REG_WRITE,reg_addr : 32'hd08   ,value : 32'd4610},
'{step_type:REG_WRITE,reg_addr : 32'hd0c   ,value : 32'd52691067},
'{step_type:REG_WRITE,reg_addr : 32'hd30   ,value : 32'd2151451263},
'{step_type:REG_WRITE,reg_addr : 32'hd34   ,value : 32'd536892214},
'{step_type:REG_WRITE,reg_addr : 32'h100500,value : 32'd1296},
'{step_type:REG_WRITE,reg_addr : 32'h100504,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h100508,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h10050c,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h200500,value : 32'd1296},
'{step_type:REG_WRITE,reg_addr : 32'h200504,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h200508,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h20050c,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h300500,value : 32'd1296},
'{step_type:REG_WRITE,reg_addr : 32'h300504,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h300508,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h30050c,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h30004 ,value : 32'd26},
'{step_type:REG_WRITE,reg_addr : 32'h3000c ,value : 32'd4131075},
'{step_type:REG_WRITE,reg_addr : 32'h30010 ,value : 32'd257},
'{step_type:REG_WRITE,reg_addr : 32'h30014 ,value : 32'd520291075},
'{step_type:REG_WRITE,reg_addr : 32'h30018 ,value : 32'd50529024},
'{step_type:REG_WRITE,reg_addr : 32'h3001c ,value : 32'd134744072},
'{step_type:REG_WRITE,reg_addr : 32'h30020 ,value : 32'd134744072},
'{step_type:REG_WRITE,reg_addr : 32'h30024 ,value : 32'd134744072},
'{step_type:REG_WRITE,reg_addr : 32'h30028 ,value : 32'd134744072},
'{step_type:REG_WRITE,reg_addr : 32'h3002c ,value : 32'd2056},
'{step_type:REG_WRITE,reg_addr : 32'h30030 ,value : 32'd16},
'{step_type:REG_WRITE,reg_addr : 32'h10b84 ,value : 32'd0},
'{step_type:REG_WRITE,reg_addr : 32'h20090 ,value : 32'd1},
'{step_type:REG_WRITE,reg_addr : 32'h10208 ,value : 32'd1},
'{step_type:REG_WRITE,reg_addr : 32'h10208 ,value : 32'd1}
}};
