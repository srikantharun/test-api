// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: {{ cookiecutter.author_full_name }} <{{ cookiecutter.author_email }}>

/// TODO:__one_line_summary_of_{{ cookiecutter.ip_name }}__
///
module {{ cookiecutter.ip_name }} #(
  /// TODO:description_of_parameter
  parameter int unsigned __parameter
)(
  /// Clock, positive edge triggered
  input  wire i_clk,
  /// Asynchronous reset, active low
  input  wire i_rst_n,


);


endmodule
