// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: Manuel Oliveira <manuel.oliveira@axelera.ai>

/// SVA of ai_core
///

`ifndef AI_CORE_SVA_SV
`define AI_CORE_SVA_SV

module ai_core_sva #(
  /// TODO:description_of_parameter
  parameter int unsigned __parameter
)(
  /// Clock, positive edge triggered
  input  wire i_clk,
  /// Asynchronous reset, active low
  input  wire i_rst_n,


);
  // =====================================================
  // Local parameters
  // =====================================================

  // =====================================================
  // Type definition
  // =====================================================

  // =====================================================
  // Signal declarations
  // =====================================================

  // =====================================================
  // Bind signals
  // =====================================================

  // =====================================================
  // Properties
  // =====================================================

  // =====================================================
  // Assumes
  // =====================================================

  // =====================================================
  // Assertions
  // =====================================================

  // =====================================================
  // Covers
  // =====================================================

endmodule

`endif // AI_CORE_SVA_SV
