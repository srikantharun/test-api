// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_h_west
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_h_west_p (
    output logic [182:0]  o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data,
    output logic          o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head,
    input  logic          i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail,
    output logic          o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld,
    input  logic [182:0]  i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data,
    input  logic          i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head,
    output logic          o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy,
    input  logic          i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail,
    input  logic          i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld,
    output logic [398:0]  o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld,
    input  logic [398:0]  i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld,
    output logic [398:0]  o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld,
    input  logic [398:0]  i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld,
    output logic [398:0]  o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld,
    input  logic [398:0]  i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld,
    output logic [398:0]  o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld,
    input  logic [398:0]  i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld,
    output logic [146:0]  o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data,
    output logic          o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head,
    input  logic          i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy,
    output logic          o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail,
    output logic          o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld,
    input  logic [146:0]  i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data,
    input  logic          i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head,
    output logic          o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy,
    input  logic          i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail,
    input  logic          i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld,
    input  wire           i_noc_clk,
    input  wire           i_noc_rst_n,
    // DFT Interface
    input  wire           tck,
    input  wire           trst,
    input  logic          tms,
    input  logic          tdi,
    output logic          tdo_en,
    output logic          tdo,
    input  wire           test_clk,
    input  logic          test_mode,
    input  logic          edt_update,
    input  logic          scan_en,
    input  logic [12-1:0] scan_in,
    output logic [12-1:0] scan_out,
    input  wire            bisr_clk,
    input  wire            bisr_reset,
    input  logic           bisr_shift_en,
    input  logic           bisr_si,
    output logic           bisr_so
);
    // -- Automatically-generated Memory Interface -- //
    localparam int unsigned MEM_INTERFACES = 8;

    axe_tcl_sram_pkg::impl_inp_t mem_impl_in;
    axe_tcl_sram_pkg::impl_oup_t mem_impl_out;
    axe_tcl_sram_pkg::impl_inp_t[MEM_INTERFACES-1:0] impl_to_mem;
    axe_tcl_sram_pkg::impl_oup_t[MEM_INTERFACES-1:0] impl_from_mem;

    logic mem_pde;
    logic mem_prn;
    logic mem_ret;

    // TODO(psarras; bronze; drive mem_pde by CSRs)
    assign mem_pde = '0;
    // TODO(psarras; bronze; connect mem_prn to CSRs)
    // assign CSR = mem_prn;
    // Wiring: 1st interface in the chain
    assign mem_impl_in = axe_tcl_sram_pkg::impl_inp_t'{
        ret: mem_ret,
        pde: mem_pde,
        se: scan_en,
        default: '0
    };
    // Wiring: Last interface in the chain
    assign mem_prn = mem_impl_out.prn;
    // Wiring: Intermediate interfaces
    axe_tcl_sram_cfg #(
        .NUM_SRAMS(MEM_INTERFACES)
    ) u_sram_cfg_impl (
        .i_s(mem_impl_in),
        .o_s(mem_impl_out),
        .o_m(impl_to_mem),
        .i_m(impl_from_mem)
    );

    noc_h_west u_noc_h_west (
    .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data),
    .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head),
    .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy(i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy),
    .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail),
    .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld(o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld),
    .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data),
    .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head),
    .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy(o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy),
    .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail),
    .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld(i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld),
    .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data),
    .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head),
    .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy(i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy),
    .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail),
    .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld(o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld),
    .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data),
    .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head),
    .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy(o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy),
    .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail),
    .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld(i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld),
    .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data),
    .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head),
    .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy(i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy),
    .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail),
    .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld(o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld),
    .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data),
    .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head),
    .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy(o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy),
    .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail),
    .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld(i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld),
    .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data),
    .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head),
    .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy(i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy),
    .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail),
    .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld(o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld),
    .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data),
    .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head),
    .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy(o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy),
    .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail),
    .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld(i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld),
    .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data),
    .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head),
    .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy(i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy),
    .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail),
    .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld(o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld),
    .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data),
    .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head),
    .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy(o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy),
    .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail),
    .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld(i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld),
    .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data),
    .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head),
    .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy),
    .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail),
    .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld),
    .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data),
    .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head),
    .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy),
    .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail),
    .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld),
    .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data),
    .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head),
    .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy),
    .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail),
    .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld),
    .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data),
    .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head),
    .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy),
    .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail),
    .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld),
    .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data),
    .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head),
    .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy),
    .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail),
    .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld),
    .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data),
    .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head),
    .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy),
    .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail),
    .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld),
    .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data),
    .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head),
    .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy),
    .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail),
    .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld),
    .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data),
    .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head),
    .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy),
    .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail),
    .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld),
    .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data),
    .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head),
    .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy),
    .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail),
    .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld),
    .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data),
    .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head),
    .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy),
    .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail),
    .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_mainpde(impl_to_mem[0].pde),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_mainprn(impl_from_mem[0].prn),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_mainret(impl_to_mem[0].ret),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_mainse(impl_to_mem[0].se),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainpde(impl_to_mem[1].pde),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainprn(impl_from_mem[1].prn),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainret(impl_to_mem[1].ret),
    .lnk_buff_512_to_256_west_to_ddr_w0_req_resp_mainse(impl_to_mem[1].se),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_mainpde(impl_to_mem[2].pde),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_mainprn(impl_from_mem[2].prn),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_mainret(impl_to_mem[2].ret),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_mainse(impl_to_mem[2].se),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainpde(impl_to_mem[3].pde),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainprn(impl_from_mem[3].prn),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainret(impl_to_mem[3].ret),
    .lnk_buff_512_to_256_west_to_ddr_w1_req_resp_mainse(impl_to_mem[3].se),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_mainpde(impl_to_mem[4].pde),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_mainprn(impl_from_mem[4].prn),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_mainret(impl_to_mem[4].ret),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_mainse(impl_to_mem[4].se),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainpde(impl_to_mem[5].pde),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainprn(impl_from_mem[5].prn),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainret(impl_to_mem[5].ret),
    .lnk_buff_512_to_256_west_to_ddr_w2_req_resp_mainse(impl_to_mem[5].se),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_mainpde(impl_to_mem[6].pde),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_mainprn(impl_from_mem[6].prn),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_mainret(impl_to_mem[6].ret),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_mainse(impl_to_mem[6].se),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainpde(impl_to_mem[7].pde),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainprn(impl_from_mem[7].prn),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainret(impl_to_mem[7].ret),
    .lnk_buff_512_to_256_west_to_ddr_w3_req_resp_mainse(impl_to_mem[7].se),
    .i_noc_clk(i_noc_clk),
    .i_noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
);

endmodule
