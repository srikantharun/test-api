`ifndef RAL_DWC_DDRCTL_MAP_REGB_ARB_PORT0_PKG
`define RAL_DWC_DDRCTL_MAP_REGB_ARB_PORT0_PKG

package ral_DWC_ddrctl_map_REGB_ARB_PORT0_pkg;
import uvm_pkg::*;

class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCCFG extends uvm_reg;
	rand uvm_reg_field go2critical_en;
	rand uvm_reg_field pagematch_limit;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   go2critical_en: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   pagematch_limit: coverpoint {m_data[4:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PCCFG");
		super.new(name, 8,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.go2critical_en = uvm_reg_field::type_id::create("go2critical_en",,get_full_name());
      this.go2critical_en.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.pagematch_limit = uvm_reg_field::type_id::create("pagematch_limit",,get_full_name());
      this.pagematch_limit.configure(this, 1, 4, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCCFG)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCCFG


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGR extends uvm_reg;
	rand uvm_reg_field rd_port_priority;
	rand uvm_reg_field rd_port_aging_en;
	rand uvm_reg_field rd_port_urgent_en;
	rand uvm_reg_field rd_port_pagematch_en;
	rand uvm_reg_field rrb_lock_threshold;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   rd_port_priority: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	   rd_port_aging_en: coverpoint {m_data[12:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   rd_port_urgent_en: coverpoint {m_data[13:13], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   rd_port_pagematch_en: coverpoint {m_data[14:14], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   rrb_lock_threshold: coverpoint {m_data[23:20], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PCFGR");
		super.new(name, 24,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.rd_port_priority = uvm_reg_field::type_id::create("rd_port_priority",,get_full_name());
      this.rd_port_priority.configure(this, 10, 0, "RW", 0, 10'h1f, 1, 0, 0);
      this.rd_port_aging_en = uvm_reg_field::type_id::create("rd_port_aging_en",,get_full_name());
      this.rd_port_aging_en.configure(this, 1, 12, "RW", 0, 1'h1, 1, 0, 0);
      this.rd_port_urgent_en = uvm_reg_field::type_id::create("rd_port_urgent_en",,get_full_name());
      this.rd_port_urgent_en.configure(this, 1, 13, "RW", 0, 1'h0, 1, 0, 0);
      this.rd_port_pagematch_en = uvm_reg_field::type_id::create("rd_port_pagematch_en",,get_full_name());
      this.rd_port_pagematch_en.configure(this, 1, 14, "RW", 0, 1'h1, 1, 0, 0);
      this.rrb_lock_threshold = uvm_reg_field::type_id::create("rrb_lock_threshold",,get_full_name());
      this.rrb_lock_threshold.configure(this, 4, 20, "RW", 0, 4'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGR)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGR


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGW extends uvm_reg;
	rand uvm_reg_field wr_port_priority;
	rand uvm_reg_field wr_port_aging_en;
	rand uvm_reg_field wr_port_urgent_en;
	rand uvm_reg_field wr_port_pagematch_en;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   wr_port_priority: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	   wr_port_aging_en: coverpoint {m_data[12:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   wr_port_urgent_en: coverpoint {m_data[13:13], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   wr_port_pagematch_en: coverpoint {m_data[14:14], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PCFGW");
		super.new(name, 16,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.wr_port_priority = uvm_reg_field::type_id::create("wr_port_priority",,get_full_name());
      this.wr_port_priority.configure(this, 10, 0, "RW", 0, 10'h1f, 1, 0, 0);
      this.wr_port_aging_en = uvm_reg_field::type_id::create("wr_port_aging_en",,get_full_name());
      this.wr_port_aging_en.configure(this, 1, 12, "RW", 0, 1'h1, 1, 0, 0);
      this.wr_port_urgent_en = uvm_reg_field::type_id::create("wr_port_urgent_en",,get_full_name());
      this.wr_port_urgent_en.configure(this, 1, 13, "RW", 0, 1'h0, 1, 0, 0);
      this.wr_port_pagematch_en = uvm_reg_field::type_id::create("wr_port_pagematch_en",,get_full_name());
      this.wr_port_pagematch_en.configure(this, 1, 14, "RW", 0, 1'h1, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGW)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGW


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCTRL extends uvm_reg;
	rand uvm_reg_field port_en;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   port_en: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PCTRL");
		super.new(name, 8,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.port_en = uvm_reg_field::type_id::create("port_en",,get_full_name());
      this.port_en.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCTRL)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCTRL


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS0 extends uvm_reg;
	rand uvm_reg_field rqos_map_level1;
	rand uvm_reg_field rqos_map_level2;
	rand uvm_reg_field rqos_map_region0;
	rand uvm_reg_field rqos_map_region1;
	rand uvm_reg_field rqos_map_region2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   rqos_map_level1: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   rqos_map_level2: coverpoint {m_data[11:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   rqos_map_region0: coverpoint {m_data[17:16], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	   rqos_map_region1: coverpoint {m_data[21:20], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	   rqos_map_region2: coverpoint {m_data[25:24], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS0");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.rqos_map_level1 = uvm_reg_field::type_id::create("rqos_map_level1",,get_full_name());
      this.rqos_map_level1.configure(this, 4, 0, "RW", 1, 4'h0, 1, 0, 1);
      this.rqos_map_level2 = uvm_reg_field::type_id::create("rqos_map_level2",,get_full_name());
      this.rqos_map_level2.configure(this, 4, 8, "RW", 1, 4'he, 1, 0, 1);
      this.rqos_map_region0 = uvm_reg_field::type_id::create("rqos_map_region0",,get_full_name());
      this.rqos_map_region0.configure(this, 2, 16, "RW", 1, 2'h0, 1, 0, 0);
      this.rqos_map_region1 = uvm_reg_field::type_id::create("rqos_map_region1",,get_full_name());
      this.rqos_map_region1.configure(this, 2, 20, "RW", 1, 2'h0, 1, 0, 0);
      this.rqos_map_region2 = uvm_reg_field::type_id::create("rqos_map_region2",,get_full_name());
      this.rqos_map_region2.configure(this, 2, 24, "RW", 1, 2'h2, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS0


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS1 extends uvm_reg;
	rand uvm_reg_field rqos_map_timeoutb;
	rand uvm_reg_field rqos_map_timeoutr;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   rqos_map_timeoutb: coverpoint {m_data[10:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {12'b??????????00};
	      wildcard bins bit_0_wr_as_1 = {12'b??????????10};
	      wildcard bins bit_0_rd_as_0 = {12'b??????????01};
	      wildcard bins bit_0_rd_as_1 = {12'b??????????11};
	      wildcard bins bit_1_wr_as_0 = {12'b?????????0?0};
	      wildcard bins bit_1_wr_as_1 = {12'b?????????1?0};
	      wildcard bins bit_1_rd_as_0 = {12'b?????????0?1};
	      wildcard bins bit_1_rd_as_1 = {12'b?????????1?1};
	      wildcard bins bit_2_wr_as_0 = {12'b????????0??0};
	      wildcard bins bit_2_wr_as_1 = {12'b????????1??0};
	      wildcard bins bit_2_rd_as_0 = {12'b????????0??1};
	      wildcard bins bit_2_rd_as_1 = {12'b????????1??1};
	      wildcard bins bit_3_wr_as_0 = {12'b???????0???0};
	      wildcard bins bit_3_wr_as_1 = {12'b???????1???0};
	      wildcard bins bit_3_rd_as_0 = {12'b???????0???1};
	      wildcard bins bit_3_rd_as_1 = {12'b???????1???1};
	      wildcard bins bit_4_wr_as_0 = {12'b??????0????0};
	      wildcard bins bit_4_wr_as_1 = {12'b??????1????0};
	      wildcard bins bit_4_rd_as_0 = {12'b??????0????1};
	      wildcard bins bit_4_rd_as_1 = {12'b??????1????1};
	      wildcard bins bit_5_wr_as_0 = {12'b?????0?????0};
	      wildcard bins bit_5_wr_as_1 = {12'b?????1?????0};
	      wildcard bins bit_5_rd_as_0 = {12'b?????0?????1};
	      wildcard bins bit_5_rd_as_1 = {12'b?????1?????1};
	      wildcard bins bit_6_wr_as_0 = {12'b????0??????0};
	      wildcard bins bit_6_wr_as_1 = {12'b????1??????0};
	      wildcard bins bit_6_rd_as_0 = {12'b????0??????1};
	      wildcard bins bit_6_rd_as_1 = {12'b????1??????1};
	      wildcard bins bit_7_wr_as_0 = {12'b???0???????0};
	      wildcard bins bit_7_wr_as_1 = {12'b???1???????0};
	      wildcard bins bit_7_rd_as_0 = {12'b???0???????1};
	      wildcard bins bit_7_rd_as_1 = {12'b???1???????1};
	      wildcard bins bit_8_wr_as_0 = {12'b??0????????0};
	      wildcard bins bit_8_wr_as_1 = {12'b??1????????0};
	      wildcard bins bit_8_rd_as_0 = {12'b??0????????1};
	      wildcard bins bit_8_rd_as_1 = {12'b??1????????1};
	      wildcard bins bit_9_wr_as_0 = {12'b?0?????????0};
	      wildcard bins bit_9_wr_as_1 = {12'b?1?????????0};
	      wildcard bins bit_9_rd_as_0 = {12'b?0?????????1};
	      wildcard bins bit_9_rd_as_1 = {12'b?1?????????1};
	      wildcard bins bit_10_wr_as_0 = {12'b0??????????0};
	      wildcard bins bit_10_wr_as_1 = {12'b1??????????0};
	      wildcard bins bit_10_rd_as_0 = {12'b0??????????1};
	      wildcard bins bit_10_rd_as_1 = {12'b1??????????1};
	      option.weight = 44;
	   }
	   rqos_map_timeoutr: coverpoint {m_data[26:16], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {12'b??????????00};
	      wildcard bins bit_0_wr_as_1 = {12'b??????????10};
	      wildcard bins bit_0_rd_as_0 = {12'b??????????01};
	      wildcard bins bit_0_rd_as_1 = {12'b??????????11};
	      wildcard bins bit_1_wr_as_0 = {12'b?????????0?0};
	      wildcard bins bit_1_wr_as_1 = {12'b?????????1?0};
	      wildcard bins bit_1_rd_as_0 = {12'b?????????0?1};
	      wildcard bins bit_1_rd_as_1 = {12'b?????????1?1};
	      wildcard bins bit_2_wr_as_0 = {12'b????????0??0};
	      wildcard bins bit_2_wr_as_1 = {12'b????????1??0};
	      wildcard bins bit_2_rd_as_0 = {12'b????????0??1};
	      wildcard bins bit_2_rd_as_1 = {12'b????????1??1};
	      wildcard bins bit_3_wr_as_0 = {12'b???????0???0};
	      wildcard bins bit_3_wr_as_1 = {12'b???????1???0};
	      wildcard bins bit_3_rd_as_0 = {12'b???????0???1};
	      wildcard bins bit_3_rd_as_1 = {12'b???????1???1};
	      wildcard bins bit_4_wr_as_0 = {12'b??????0????0};
	      wildcard bins bit_4_wr_as_1 = {12'b??????1????0};
	      wildcard bins bit_4_rd_as_0 = {12'b??????0????1};
	      wildcard bins bit_4_rd_as_1 = {12'b??????1????1};
	      wildcard bins bit_5_wr_as_0 = {12'b?????0?????0};
	      wildcard bins bit_5_wr_as_1 = {12'b?????1?????0};
	      wildcard bins bit_5_rd_as_0 = {12'b?????0?????1};
	      wildcard bins bit_5_rd_as_1 = {12'b?????1?????1};
	      wildcard bins bit_6_wr_as_0 = {12'b????0??????0};
	      wildcard bins bit_6_wr_as_1 = {12'b????1??????0};
	      wildcard bins bit_6_rd_as_0 = {12'b????0??????1};
	      wildcard bins bit_6_rd_as_1 = {12'b????1??????1};
	      wildcard bins bit_7_wr_as_0 = {12'b???0???????0};
	      wildcard bins bit_7_wr_as_1 = {12'b???1???????0};
	      wildcard bins bit_7_rd_as_0 = {12'b???0???????1};
	      wildcard bins bit_7_rd_as_1 = {12'b???1???????1};
	      wildcard bins bit_8_wr_as_0 = {12'b??0????????0};
	      wildcard bins bit_8_wr_as_1 = {12'b??1????????0};
	      wildcard bins bit_8_rd_as_0 = {12'b??0????????1};
	      wildcard bins bit_8_rd_as_1 = {12'b??1????????1};
	      wildcard bins bit_9_wr_as_0 = {12'b?0?????????0};
	      wildcard bins bit_9_wr_as_1 = {12'b?1?????????0};
	      wildcard bins bit_9_rd_as_0 = {12'b?0?????????1};
	      wildcard bins bit_9_rd_as_1 = {12'b?1?????????1};
	      wildcard bins bit_10_wr_as_0 = {12'b0??????????0};
	      wildcard bins bit_10_wr_as_1 = {12'b1??????????0};
	      wildcard bins bit_10_rd_as_0 = {12'b0??????????1};
	      wildcard bins bit_10_rd_as_1 = {12'b1??????????1};
	      option.weight = 44;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS1");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.rqos_map_timeoutb = uvm_reg_field::type_id::create("rqos_map_timeoutb",,get_full_name());
      this.rqos_map_timeoutb.configure(this, 11, 0, "RW", 1, 11'h0, 1, 0, 1);
      this.rqos_map_timeoutr = uvm_reg_field::type_id::create("rqos_map_timeoutr",,get_full_name());
      this.rqos_map_timeoutr.configure(this, 11, 16, "RW", 1, 11'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS1


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS0 extends uvm_reg;
	rand uvm_reg_field wqos_map_level1;
	rand uvm_reg_field wqos_map_level2;
	rand uvm_reg_field wqos_map_region0;
	rand uvm_reg_field wqos_map_region1;
	rand uvm_reg_field wqos_map_region2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   wqos_map_level1: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   wqos_map_level2: coverpoint {m_data[11:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   wqos_map_region0: coverpoint {m_data[17:16], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	   wqos_map_region1: coverpoint {m_data[21:20], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	   wqos_map_region2: coverpoint {m_data[25:24], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	constraint wqos_map_level1_valid {
		wqos_map_level1.value < 14; 			
	}
	constraint wqos_map_level2_valid {
		wqos_map_level2.value < 15; 			
	}
	constraint wqos_map_region0_valid {
		wqos_map_region0.value < 2; 			
	}
	constraint wqos_map_region1_valid {
		wqos_map_region1.value < 2; 			
	}
	constraint wqos_map_region2_valid {
		wqos_map_region2.value < 2; 			
	}

	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS0");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.wqos_map_level1 = uvm_reg_field::type_id::create("wqos_map_level1",,get_full_name());
      this.wqos_map_level1.configure(this, 4, 0, "RW", 1, 4'h0, 1, 1, 1);
      this.wqos_map_level2 = uvm_reg_field::type_id::create("wqos_map_level2",,get_full_name());
      this.wqos_map_level2.configure(this, 4, 8, "RW", 1, 4'he, 1, 1, 1);
      this.wqos_map_region0 = uvm_reg_field::type_id::create("wqos_map_region0",,get_full_name());
      this.wqos_map_region0.configure(this, 2, 16, "RW", 1, 2'h0, 1, 1, 0);
      this.wqos_map_region1 = uvm_reg_field::type_id::create("wqos_map_region1",,get_full_name());
      this.wqos_map_region1.configure(this, 2, 20, "RW", 1, 2'h0, 1, 1, 0);
      this.wqos_map_region2 = uvm_reg_field::type_id::create("wqos_map_region2",,get_full_name());
      this.wqos_map_region2.configure(this, 2, 24, "RW", 1, 2'h0, 1, 1, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS0


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS1 extends uvm_reg;
	rand uvm_reg_field wqos_map_timeout1;
	rand uvm_reg_field wqos_map_timeout2;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   wqos_map_timeout1: coverpoint {m_data[10:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {12'b??????????00};
	      wildcard bins bit_0_wr_as_1 = {12'b??????????10};
	      wildcard bins bit_0_rd_as_0 = {12'b??????????01};
	      wildcard bins bit_0_rd_as_1 = {12'b??????????11};
	      wildcard bins bit_1_wr_as_0 = {12'b?????????0?0};
	      wildcard bins bit_1_wr_as_1 = {12'b?????????1?0};
	      wildcard bins bit_1_rd_as_0 = {12'b?????????0?1};
	      wildcard bins bit_1_rd_as_1 = {12'b?????????1?1};
	      wildcard bins bit_2_wr_as_0 = {12'b????????0??0};
	      wildcard bins bit_2_wr_as_1 = {12'b????????1??0};
	      wildcard bins bit_2_rd_as_0 = {12'b????????0??1};
	      wildcard bins bit_2_rd_as_1 = {12'b????????1??1};
	      wildcard bins bit_3_wr_as_0 = {12'b???????0???0};
	      wildcard bins bit_3_wr_as_1 = {12'b???????1???0};
	      wildcard bins bit_3_rd_as_0 = {12'b???????0???1};
	      wildcard bins bit_3_rd_as_1 = {12'b???????1???1};
	      wildcard bins bit_4_wr_as_0 = {12'b??????0????0};
	      wildcard bins bit_4_wr_as_1 = {12'b??????1????0};
	      wildcard bins bit_4_rd_as_0 = {12'b??????0????1};
	      wildcard bins bit_4_rd_as_1 = {12'b??????1????1};
	      wildcard bins bit_5_wr_as_0 = {12'b?????0?????0};
	      wildcard bins bit_5_wr_as_1 = {12'b?????1?????0};
	      wildcard bins bit_5_rd_as_0 = {12'b?????0?????1};
	      wildcard bins bit_5_rd_as_1 = {12'b?????1?????1};
	      wildcard bins bit_6_wr_as_0 = {12'b????0??????0};
	      wildcard bins bit_6_wr_as_1 = {12'b????1??????0};
	      wildcard bins bit_6_rd_as_0 = {12'b????0??????1};
	      wildcard bins bit_6_rd_as_1 = {12'b????1??????1};
	      wildcard bins bit_7_wr_as_0 = {12'b???0???????0};
	      wildcard bins bit_7_wr_as_1 = {12'b???1???????0};
	      wildcard bins bit_7_rd_as_0 = {12'b???0???????1};
	      wildcard bins bit_7_rd_as_1 = {12'b???1???????1};
	      wildcard bins bit_8_wr_as_0 = {12'b??0????????0};
	      wildcard bins bit_8_wr_as_1 = {12'b??1????????0};
	      wildcard bins bit_8_rd_as_0 = {12'b??0????????1};
	      wildcard bins bit_8_rd_as_1 = {12'b??1????????1};
	      wildcard bins bit_9_wr_as_0 = {12'b?0?????????0};
	      wildcard bins bit_9_wr_as_1 = {12'b?1?????????0};
	      wildcard bins bit_9_rd_as_0 = {12'b?0?????????1};
	      wildcard bins bit_9_rd_as_1 = {12'b?1?????????1};
	      wildcard bins bit_10_wr_as_0 = {12'b0??????????0};
	      wildcard bins bit_10_wr_as_1 = {12'b1??????????0};
	      wildcard bins bit_10_rd_as_0 = {12'b0??????????1};
	      wildcard bins bit_10_rd_as_1 = {12'b1??????????1};
	      option.weight = 44;
	   }
	   wqos_map_timeout2: coverpoint {m_data[26:16], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {12'b??????????00};
	      wildcard bins bit_0_wr_as_1 = {12'b??????????10};
	      wildcard bins bit_0_rd_as_0 = {12'b??????????01};
	      wildcard bins bit_0_rd_as_1 = {12'b??????????11};
	      wildcard bins bit_1_wr_as_0 = {12'b?????????0?0};
	      wildcard bins bit_1_wr_as_1 = {12'b?????????1?0};
	      wildcard bins bit_1_rd_as_0 = {12'b?????????0?1};
	      wildcard bins bit_1_rd_as_1 = {12'b?????????1?1};
	      wildcard bins bit_2_wr_as_0 = {12'b????????0??0};
	      wildcard bins bit_2_wr_as_1 = {12'b????????1??0};
	      wildcard bins bit_2_rd_as_0 = {12'b????????0??1};
	      wildcard bins bit_2_rd_as_1 = {12'b????????1??1};
	      wildcard bins bit_3_wr_as_0 = {12'b???????0???0};
	      wildcard bins bit_3_wr_as_1 = {12'b???????1???0};
	      wildcard bins bit_3_rd_as_0 = {12'b???????0???1};
	      wildcard bins bit_3_rd_as_1 = {12'b???????1???1};
	      wildcard bins bit_4_wr_as_0 = {12'b??????0????0};
	      wildcard bins bit_4_wr_as_1 = {12'b??????1????0};
	      wildcard bins bit_4_rd_as_0 = {12'b??????0????1};
	      wildcard bins bit_4_rd_as_1 = {12'b??????1????1};
	      wildcard bins bit_5_wr_as_0 = {12'b?????0?????0};
	      wildcard bins bit_5_wr_as_1 = {12'b?????1?????0};
	      wildcard bins bit_5_rd_as_0 = {12'b?????0?????1};
	      wildcard bins bit_5_rd_as_1 = {12'b?????1?????1};
	      wildcard bins bit_6_wr_as_0 = {12'b????0??????0};
	      wildcard bins bit_6_wr_as_1 = {12'b????1??????0};
	      wildcard bins bit_6_rd_as_0 = {12'b????0??????1};
	      wildcard bins bit_6_rd_as_1 = {12'b????1??????1};
	      wildcard bins bit_7_wr_as_0 = {12'b???0???????0};
	      wildcard bins bit_7_wr_as_1 = {12'b???1???????0};
	      wildcard bins bit_7_rd_as_0 = {12'b???0???????1};
	      wildcard bins bit_7_rd_as_1 = {12'b???1???????1};
	      wildcard bins bit_8_wr_as_0 = {12'b??0????????0};
	      wildcard bins bit_8_wr_as_1 = {12'b??1????????0};
	      wildcard bins bit_8_rd_as_0 = {12'b??0????????1};
	      wildcard bins bit_8_rd_as_1 = {12'b??1????????1};
	      wildcard bins bit_9_wr_as_0 = {12'b?0?????????0};
	      wildcard bins bit_9_wr_as_1 = {12'b?1?????????0};
	      wildcard bins bit_9_rd_as_0 = {12'b?0?????????1};
	      wildcard bins bit_9_rd_as_1 = {12'b?1?????????1};
	      wildcard bins bit_10_wr_as_0 = {12'b0??????????0};
	      wildcard bins bit_10_wr_as_1 = {12'b1??????????0};
	      wildcard bins bit_10_rd_as_0 = {12'b0??????????1};
	      wildcard bins bit_10_rd_as_1 = {12'b1??????????1};
	      option.weight = 44;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS1");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.wqos_map_timeout1 = uvm_reg_field::type_id::create("wqos_map_timeout1",,get_full_name());
      this.wqos_map_timeout1.configure(this, 11, 0, "RW", 1, 11'h0, 1, 0, 1);
      this.wqos_map_timeout2 = uvm_reg_field::type_id::create("wqos_map_timeout2",,get_full_name());
      this.wqos_map_timeout2.configure(this, 11, 16, "RW", 1, 11'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS1


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRCTL extends uvm_reg;
	rand uvm_reg_field scrub_en;
	rand uvm_reg_field scrub_during_lowpower;
	rand uvm_reg_field scrub_burst_length_nm;
	rand uvm_reg_field scrub_interval;
	rand uvm_reg_field scrub_cmd_type;
	rand uvm_reg_field scrub_burst_length_lp;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   scrub_en: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   scrub_during_lowpower: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   scrub_burst_length_nm: coverpoint {m_data[6:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	   scrub_interval: coverpoint {m_data[20:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {14'b????????????00};
	      wildcard bins bit_0_wr_as_1 = {14'b????????????10};
	      wildcard bins bit_0_rd_as_0 = {14'b????????????01};
	      wildcard bins bit_0_rd_as_1 = {14'b????????????11};
	      wildcard bins bit_1_wr_as_0 = {14'b???????????0?0};
	      wildcard bins bit_1_wr_as_1 = {14'b???????????1?0};
	      wildcard bins bit_1_rd_as_0 = {14'b???????????0?1};
	      wildcard bins bit_1_rd_as_1 = {14'b???????????1?1};
	      wildcard bins bit_2_wr_as_0 = {14'b??????????0??0};
	      wildcard bins bit_2_wr_as_1 = {14'b??????????1??0};
	      wildcard bins bit_2_rd_as_0 = {14'b??????????0??1};
	      wildcard bins bit_2_rd_as_1 = {14'b??????????1??1};
	      wildcard bins bit_3_wr_as_0 = {14'b?????????0???0};
	      wildcard bins bit_3_wr_as_1 = {14'b?????????1???0};
	      wildcard bins bit_3_rd_as_0 = {14'b?????????0???1};
	      wildcard bins bit_3_rd_as_1 = {14'b?????????1???1};
	      wildcard bins bit_4_wr_as_0 = {14'b????????0????0};
	      wildcard bins bit_4_wr_as_1 = {14'b????????1????0};
	      wildcard bins bit_4_rd_as_0 = {14'b????????0????1};
	      wildcard bins bit_4_rd_as_1 = {14'b????????1????1};
	      wildcard bins bit_5_wr_as_0 = {14'b???????0?????0};
	      wildcard bins bit_5_wr_as_1 = {14'b???????1?????0};
	      wildcard bins bit_5_rd_as_0 = {14'b???????0?????1};
	      wildcard bins bit_5_rd_as_1 = {14'b???????1?????1};
	      wildcard bins bit_6_wr_as_0 = {14'b??????0??????0};
	      wildcard bins bit_6_wr_as_1 = {14'b??????1??????0};
	      wildcard bins bit_6_rd_as_0 = {14'b??????0??????1};
	      wildcard bins bit_6_rd_as_1 = {14'b??????1??????1};
	      wildcard bins bit_7_wr_as_0 = {14'b?????0???????0};
	      wildcard bins bit_7_wr_as_1 = {14'b?????1???????0};
	      wildcard bins bit_7_rd_as_0 = {14'b?????0???????1};
	      wildcard bins bit_7_rd_as_1 = {14'b?????1???????1};
	      wildcard bins bit_8_wr_as_0 = {14'b????0????????0};
	      wildcard bins bit_8_wr_as_1 = {14'b????1????????0};
	      wildcard bins bit_8_rd_as_0 = {14'b????0????????1};
	      wildcard bins bit_8_rd_as_1 = {14'b????1????????1};
	      wildcard bins bit_9_wr_as_0 = {14'b???0?????????0};
	      wildcard bins bit_9_wr_as_1 = {14'b???1?????????0};
	      wildcard bins bit_9_rd_as_0 = {14'b???0?????????1};
	      wildcard bins bit_9_rd_as_1 = {14'b???1?????????1};
	      wildcard bins bit_10_wr_as_0 = {14'b??0??????????0};
	      wildcard bins bit_10_wr_as_1 = {14'b??1??????????0};
	      wildcard bins bit_10_rd_as_0 = {14'b??0??????????1};
	      wildcard bins bit_10_rd_as_1 = {14'b??1??????????1};
	      wildcard bins bit_11_wr_as_0 = {14'b?0???????????0};
	      wildcard bins bit_11_wr_as_1 = {14'b?1???????????0};
	      wildcard bins bit_11_rd_as_0 = {14'b?0???????????1};
	      wildcard bins bit_11_rd_as_1 = {14'b?1???????????1};
	      wildcard bins bit_12_wr_as_0 = {14'b0????????????0};
	      wildcard bins bit_12_wr_as_1 = {14'b1????????????0};
	      wildcard bins bit_12_rd_as_0 = {14'b0????????????1};
	      wildcard bins bit_12_rd_as_1 = {14'b1????????????1};
	      option.weight = 52;
	   }
	   scrub_cmd_type: coverpoint {m_data[25:24], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	   scrub_burst_length_lp: coverpoint {m_data[30:28], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_SBRCTL");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.scrub_en = uvm_reg_field::type_id::create("scrub_en",,get_full_name());
      this.scrub_en.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.scrub_during_lowpower = uvm_reg_field::type_id::create("scrub_during_lowpower",,get_full_name());
      this.scrub_during_lowpower.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.scrub_burst_length_nm = uvm_reg_field::type_id::create("scrub_burst_length_nm",,get_full_name());
      this.scrub_burst_length_nm.configure(this, 3, 4, "RW", 0, 3'h1, 1, 0, 0);
      this.scrub_interval = uvm_reg_field::type_id::create("scrub_interval",,get_full_name());
      this.scrub_interval.configure(this, 13, 8, "RW", 0, 13'hff, 1, 0, 1);
      this.scrub_cmd_type = uvm_reg_field::type_id::create("scrub_cmd_type",,get_full_name());
      this.scrub_cmd_type.configure(this, 2, 24, "RW", 0, 2'h0, 1, 0, 0);
      this.scrub_burst_length_lp = uvm_reg_field::type_id::create("scrub_burst_length_lp",,get_full_name());
      this.scrub_burst_length_lp.configure(this, 3, 28, "RW", 0, 3'h1, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRCTL)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRCTL


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTAT extends uvm_reg;
	uvm_reg_field scrub_busy;
	uvm_reg_field scrub_done;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   scrub_busy: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   scrub_done: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTAT");
		super.new(name, 8,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.scrub_busy = uvm_reg_field::type_id::create("scrub_busy",,get_full_name());
      this.scrub_busy.configure(this, 1, 0, "RO", 0, 1'h0, 1, 0, 0);
      this.scrub_done = uvm_reg_field::type_id::create("scrub_done",,get_full_name());
      this.scrub_done.configure(this, 1, 1, "RO", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTAT)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTAT


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRWDATA0 extends uvm_reg;
	rand uvm_reg_field scrub_pattern0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   scrub_pattern0: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_SBRWDATA0");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.scrub_pattern0 = uvm_reg_field::type_id::create("scrub_pattern0",,get_full_name());
      this.scrub_pattern0.configure(this, 32, 0, "RW", 0, 32'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRWDATA0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRWDATA0


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART0 extends uvm_reg;
	rand uvm_reg_field sbr_address_start_mask_0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   sbr_address_start_mask_0: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART0");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.sbr_address_start_mask_0 = uvm_reg_field::type_id::create("sbr_address_start_mask_0",,get_full_name());
      this.sbr_address_start_mask_0.configure(this, 32, 0, "RW", 0, 32'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART0


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART1 extends uvm_reg;
	rand uvm_reg_field sbr_address_start_mask_1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   sbr_address_start_mask_1: coverpoint {m_data[7:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd_as_0 = {9'b???????01};
	      wildcard bins bit_0_rd_as_1 = {9'b???????11};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd_as_0 = {9'b??????0?1};
	      wildcard bins bit_1_rd_as_1 = {9'b??????1?1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd_as_0 = {9'b?????0??1};
	      wildcard bins bit_2_rd_as_1 = {9'b?????1??1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd_as_0 = {9'b????0???1};
	      wildcard bins bit_3_rd_as_1 = {9'b????1???1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd_as_0 = {9'b???0????1};
	      wildcard bins bit_4_rd_as_1 = {9'b???1????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd_as_0 = {9'b??0?????1};
	      wildcard bins bit_5_rd_as_1 = {9'b??1?????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd_as_0 = {9'b?0??????1};
	      wildcard bins bit_6_rd_as_1 = {9'b?1??????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd_as_0 = {9'b0???????1};
	      wildcard bins bit_7_rd_as_1 = {9'b1???????1};
	      option.weight = 32;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART1");
		super.new(name, 8,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.sbr_address_start_mask_1 = uvm_reg_field::type_id::create("sbr_address_start_mask_1",,get_full_name());
      this.sbr_address_start_mask_1.configure(this, 8, 0, "RW", 0, 8'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART1


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE0 extends uvm_reg;
	rand uvm_reg_field sbr_address_range_mask_0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   sbr_address_range_mask_0: coverpoint {m_data[31:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {33'b???????????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {33'b???????????????????????????????10};
	      wildcard bins bit_0_rd_as_0 = {33'b???????????????????????????????01};
	      wildcard bins bit_0_rd_as_1 = {33'b???????????????????????????????11};
	      wildcard bins bit_1_wr_as_0 = {33'b??????????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {33'b??????????????????????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {33'b??????????????????????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {33'b??????????????????????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {33'b?????????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {33'b?????????????????????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {33'b?????????????????????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {33'b?????????????????????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {33'b????????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {33'b????????????????????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {33'b????????????????????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {33'b????????????????????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {33'b???????????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {33'b???????????????????????????1????0};
	      wildcard bins bit_4_rd_as_0 = {33'b???????????????????????????0????1};
	      wildcard bins bit_4_rd_as_1 = {33'b???????????????????????????1????1};
	      wildcard bins bit_5_wr_as_0 = {33'b??????????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {33'b??????????????????????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {33'b??????????????????????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {33'b??????????????????????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {33'b?????????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {33'b?????????????????????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {33'b?????????????????????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {33'b?????????????????????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {33'b????????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {33'b????????????????????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {33'b????????????????????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {33'b????????????????????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {33'b???????????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {33'b???????????????????????1????????0};
	      wildcard bins bit_8_rd_as_0 = {33'b???????????????????????0????????1};
	      wildcard bins bit_8_rd_as_1 = {33'b???????????????????????1????????1};
	      wildcard bins bit_9_wr_as_0 = {33'b??????????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {33'b??????????????????????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {33'b??????????????????????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {33'b??????????????????????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {33'b?????????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {33'b?????????????????????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {33'b?????????????????????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {33'b?????????????????????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {33'b????????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {33'b????????????????????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {33'b????????????????????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {33'b????????????????????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {33'b???????????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {33'b???????????????????1????????????0};
	      wildcard bins bit_12_rd_as_0 = {33'b???????????????????0????????????1};
	      wildcard bins bit_12_rd_as_1 = {33'b???????????????????1????????????1};
	      wildcard bins bit_13_wr_as_0 = {33'b??????????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {33'b??????????????????1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {33'b??????????????????0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {33'b??????????????????1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {33'b?????????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {33'b?????????????????1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {33'b?????????????????0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {33'b?????????????????1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {33'b????????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {33'b????????????????1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {33'b????????????????0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {33'b????????????????1???????????????1};
	      wildcard bins bit_16_wr_as_0 = {33'b???????????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {33'b???????????????1????????????????0};
	      wildcard bins bit_16_rd_as_0 = {33'b???????????????0????????????????1};
	      wildcard bins bit_16_rd_as_1 = {33'b???????????????1????????????????1};
	      wildcard bins bit_17_wr_as_0 = {33'b??????????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {33'b??????????????1?????????????????0};
	      wildcard bins bit_17_rd_as_0 = {33'b??????????????0?????????????????1};
	      wildcard bins bit_17_rd_as_1 = {33'b??????????????1?????????????????1};
	      wildcard bins bit_18_wr_as_0 = {33'b?????????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {33'b?????????????1??????????????????0};
	      wildcard bins bit_18_rd_as_0 = {33'b?????????????0??????????????????1};
	      wildcard bins bit_18_rd_as_1 = {33'b?????????????1??????????????????1};
	      wildcard bins bit_19_wr_as_0 = {33'b????????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {33'b????????????1???????????????????0};
	      wildcard bins bit_19_rd_as_0 = {33'b????????????0???????????????????1};
	      wildcard bins bit_19_rd_as_1 = {33'b????????????1???????????????????1};
	      wildcard bins bit_20_wr_as_0 = {33'b???????????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {33'b???????????1????????????????????0};
	      wildcard bins bit_20_rd_as_0 = {33'b???????????0????????????????????1};
	      wildcard bins bit_20_rd_as_1 = {33'b???????????1????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {33'b??????????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {33'b??????????1?????????????????????0};
	      wildcard bins bit_21_rd_as_0 = {33'b??????????0?????????????????????1};
	      wildcard bins bit_21_rd_as_1 = {33'b??????????1?????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {33'b?????????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {33'b?????????1??????????????????????0};
	      wildcard bins bit_22_rd_as_0 = {33'b?????????0??????????????????????1};
	      wildcard bins bit_22_rd_as_1 = {33'b?????????1??????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {33'b????????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {33'b????????1???????????????????????0};
	      wildcard bins bit_23_rd_as_0 = {33'b????????0???????????????????????1};
	      wildcard bins bit_23_rd_as_1 = {33'b????????1???????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {33'b???????0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {33'b???????1????????????????????????0};
	      wildcard bins bit_24_rd_as_0 = {33'b???????0????????????????????????1};
	      wildcard bins bit_24_rd_as_1 = {33'b???????1????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {33'b??????0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {33'b??????1?????????????????????????0};
	      wildcard bins bit_25_rd_as_0 = {33'b??????0?????????????????????????1};
	      wildcard bins bit_25_rd_as_1 = {33'b??????1?????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {33'b?????0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {33'b?????1??????????????????????????0};
	      wildcard bins bit_26_rd_as_0 = {33'b?????0??????????????????????????1};
	      wildcard bins bit_26_rd_as_1 = {33'b?????1??????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {33'b????0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {33'b????1???????????????????????????0};
	      wildcard bins bit_27_rd_as_0 = {33'b????0???????????????????????????1};
	      wildcard bins bit_27_rd_as_1 = {33'b????1???????????????????????????1};
	      wildcard bins bit_28_wr_as_0 = {33'b???0????????????????????????????0};
	      wildcard bins bit_28_wr_as_1 = {33'b???1????????????????????????????0};
	      wildcard bins bit_28_rd_as_0 = {33'b???0????????????????????????????1};
	      wildcard bins bit_28_rd_as_1 = {33'b???1????????????????????????????1};
	      wildcard bins bit_29_wr_as_0 = {33'b??0?????????????????????????????0};
	      wildcard bins bit_29_wr_as_1 = {33'b??1?????????????????????????????0};
	      wildcard bins bit_29_rd_as_0 = {33'b??0?????????????????????????????1};
	      wildcard bins bit_29_rd_as_1 = {33'b??1?????????????????????????????1};
	      wildcard bins bit_30_wr_as_0 = {33'b?0??????????????????????????????0};
	      wildcard bins bit_30_wr_as_1 = {33'b?1??????????????????????????????0};
	      wildcard bins bit_30_rd_as_0 = {33'b?0??????????????????????????????1};
	      wildcard bins bit_30_rd_as_1 = {33'b?1??????????????????????????????1};
	      wildcard bins bit_31_wr_as_0 = {33'b0???????????????????????????????0};
	      wildcard bins bit_31_wr_as_1 = {33'b1???????????????????????????????0};
	      wildcard bins bit_31_rd_as_0 = {33'b0???????????????????????????????1};
	      wildcard bins bit_31_rd_as_1 = {33'b1???????????????????????????????1};
	      option.weight = 128;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE0");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.sbr_address_range_mask_0 = uvm_reg_field::type_id::create("sbr_address_range_mask_0",,get_full_name());
      this.sbr_address_range_mask_0.configure(this, 32, 0, "RW", 0, 32'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE0)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE0


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE1 extends uvm_reg;
	rand uvm_reg_field sbr_address_range_mask_1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   sbr_address_range_mask_1: coverpoint {m_data[7:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd_as_0 = {9'b???????01};
	      wildcard bins bit_0_rd_as_1 = {9'b???????11};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd_as_0 = {9'b??????0?1};
	      wildcard bins bit_1_rd_as_1 = {9'b??????1?1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd_as_0 = {9'b?????0??1};
	      wildcard bins bit_2_rd_as_1 = {9'b?????1??1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd_as_0 = {9'b????0???1};
	      wildcard bins bit_3_rd_as_1 = {9'b????1???1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd_as_0 = {9'b???0????1};
	      wildcard bins bit_4_rd_as_1 = {9'b???1????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd_as_0 = {9'b??0?????1};
	      wildcard bins bit_5_rd_as_1 = {9'b??1?????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd_as_0 = {9'b?0??????1};
	      wildcard bins bit_6_rd_as_1 = {9'b?1??????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd_as_0 = {9'b0???????1};
	      wildcard bins bit_7_rd_as_1 = {9'b1???????1};
	      option.weight = 32;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE1");
		super.new(name, 8,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.sbr_address_range_mask_1 = uvm_reg_field::type_id::create("sbr_address_range_mask_1",,get_full_name());
      this.sbr_address_range_mask_1.configure(this, 8, 0, "RW", 0, 8'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE1


class ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PSTAT extends uvm_reg;
	uvm_reg_field rd_port_busy_0;
	uvm_reg_field wr_port_busy_0;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   rd_port_busy_0: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   wr_port_busy_0: coverpoint {m_data[16:16], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0_PSTAT");
		super.new(name, 24,build_coverage(UVM_CVR_REG_BITS));
		add_coverage(build_coverage(UVM_CVR_REG_BITS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.rd_port_busy_0 = uvm_reg_field::type_id::create("rd_port_busy_0",,get_full_name());
      this.rd_port_busy_0.configure(this, 1, 0, "RO", 0, 1'h0, 1, 0, 1);
      this.wr_port_busy_0 = uvm_reg_field::type_id::create("wr_port_busy_0",,get_full_name());
      this.wr_port_busy_0.configure(this, 1, 16, "RO", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PSTAT)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PSTAT


class ral_block_DWC_ddrctl_map_REGB_ARB_PORT0 extends uvm_reg_block;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCCFG PCCFG;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGR PCFGR;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGW PCFGW;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCTRL PCTRL;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS0 PCFGQOS0;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS1 PCFGQOS1;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS0 PCFGWQOS0;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS1 PCFGWQOS1;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRCTL SBRCTL;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTAT SBRSTAT;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRWDATA0 SBRWDATA0;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART0 SBRSTART0;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART1 SBRSTART1;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE0 SBRRANGE0;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE1 SBRRANGE1;
	rand ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PSTAT PSTAT;
   local uvm_reg_data_t m_offset;
	rand uvm_reg_field PCCFG_go2critical_en;
	rand uvm_reg_field go2critical_en;
	rand uvm_reg_field PCCFG_pagematch_limit;
	rand uvm_reg_field pagematch_limit;
	rand uvm_reg_field PCFGR_rd_port_priority;
	rand uvm_reg_field rd_port_priority;
	rand uvm_reg_field PCFGR_rd_port_aging_en;
	rand uvm_reg_field rd_port_aging_en;
	rand uvm_reg_field PCFGR_rd_port_urgent_en;
	rand uvm_reg_field rd_port_urgent_en;
	rand uvm_reg_field PCFGR_rd_port_pagematch_en;
	rand uvm_reg_field rd_port_pagematch_en;
	rand uvm_reg_field PCFGR_rrb_lock_threshold;
	rand uvm_reg_field rrb_lock_threshold;
	rand uvm_reg_field PCFGW_wr_port_priority;
	rand uvm_reg_field wr_port_priority;
	rand uvm_reg_field PCFGW_wr_port_aging_en;
	rand uvm_reg_field wr_port_aging_en;
	rand uvm_reg_field PCFGW_wr_port_urgent_en;
	rand uvm_reg_field wr_port_urgent_en;
	rand uvm_reg_field PCFGW_wr_port_pagematch_en;
	rand uvm_reg_field wr_port_pagematch_en;
	rand uvm_reg_field PCTRL_port_en;
	rand uvm_reg_field port_en;
	rand uvm_reg_field PCFGQOS0_rqos_map_level1;
	rand uvm_reg_field rqos_map_level1;
	rand uvm_reg_field PCFGQOS0_rqos_map_level2;
	rand uvm_reg_field rqos_map_level2;
	rand uvm_reg_field PCFGQOS0_rqos_map_region0;
	rand uvm_reg_field rqos_map_region0;
	rand uvm_reg_field PCFGQOS0_rqos_map_region1;
	rand uvm_reg_field rqos_map_region1;
	rand uvm_reg_field PCFGQOS0_rqos_map_region2;
	rand uvm_reg_field rqos_map_region2;
	rand uvm_reg_field PCFGQOS1_rqos_map_timeoutb;
	rand uvm_reg_field rqos_map_timeoutb;
	rand uvm_reg_field PCFGQOS1_rqos_map_timeoutr;
	rand uvm_reg_field rqos_map_timeoutr;
	rand uvm_reg_field PCFGWQOS0_wqos_map_level1;
	rand uvm_reg_field wqos_map_level1;
	rand uvm_reg_field PCFGWQOS0_wqos_map_level2;
	rand uvm_reg_field wqos_map_level2;
	rand uvm_reg_field PCFGWQOS0_wqos_map_region0;
	rand uvm_reg_field wqos_map_region0;
	rand uvm_reg_field PCFGWQOS0_wqos_map_region1;
	rand uvm_reg_field wqos_map_region1;
	rand uvm_reg_field PCFGWQOS0_wqos_map_region2;
	rand uvm_reg_field wqos_map_region2;
	rand uvm_reg_field PCFGWQOS1_wqos_map_timeout1;
	rand uvm_reg_field wqos_map_timeout1;
	rand uvm_reg_field PCFGWQOS1_wqos_map_timeout2;
	rand uvm_reg_field wqos_map_timeout2;
	rand uvm_reg_field SBRCTL_scrub_en;
	rand uvm_reg_field scrub_en;
	rand uvm_reg_field SBRCTL_scrub_during_lowpower;
	rand uvm_reg_field scrub_during_lowpower;
	rand uvm_reg_field SBRCTL_scrub_burst_length_nm;
	rand uvm_reg_field scrub_burst_length_nm;
	rand uvm_reg_field SBRCTL_scrub_interval;
	rand uvm_reg_field scrub_interval;
	rand uvm_reg_field SBRCTL_scrub_cmd_type;
	rand uvm_reg_field scrub_cmd_type;
	rand uvm_reg_field SBRCTL_scrub_burst_length_lp;
	rand uvm_reg_field scrub_burst_length_lp;
	uvm_reg_field SBRSTAT_scrub_busy;
	uvm_reg_field scrub_busy;
	uvm_reg_field SBRSTAT_scrub_done;
	uvm_reg_field scrub_done;
	rand uvm_reg_field SBRWDATA0_scrub_pattern0;
	rand uvm_reg_field scrub_pattern0;
	rand uvm_reg_field SBRSTART0_sbr_address_start_mask_0;
	rand uvm_reg_field sbr_address_start_mask_0;
	rand uvm_reg_field SBRSTART1_sbr_address_start_mask_1;
	rand uvm_reg_field sbr_address_start_mask_1;
	rand uvm_reg_field SBRRANGE0_sbr_address_range_mask_0;
	rand uvm_reg_field sbr_address_range_mask_0;
	rand uvm_reg_field SBRRANGE1_sbr_address_range_mask_1;
	rand uvm_reg_field sbr_address_range_mask_1;
	uvm_reg_field PSTAT_rd_port_busy_0;
	uvm_reg_field rd_port_busy_0;
	uvm_reg_field PSTAT_wr_port_busy_0;
	uvm_reg_field wr_port_busy_0;


	covergroup cg_addr (input string name);
	option.per_instance = 1;
option.name = get_name();

	PCCFG : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h0 };
		option.weight = 1;
	}

	PCFGR : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h4 };
		option.weight = 1;
	}

	PCFGW : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h8 };
		option.weight = 1;
	}

	PCTRL : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h90 };
		option.weight = 1;
	}

	PCFGQOS0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h94 };
		option.weight = 1;
	}

	PCFGQOS1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h98 };
		option.weight = 1;
	}

	PCFGWQOS0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h9C };
		option.weight = 1;
	}

	PCFGWQOS1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hA0 };
		option.weight = 1;
	}

	SBRCTL : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE0 };
		option.weight = 1;
	}

	SBRSTAT : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE4 };
		option.weight = 1;
	}

	SBRWDATA0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE8 };
		option.weight = 1;
	}

	SBRSTART0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hF0 };
		option.weight = 1;
	}

	SBRSTART1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hF4 };
		option.weight = 1;
	}

	SBRRANGE0 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hF8 };
		option.weight = 1;
	}

	SBRRANGE1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hFC };
		option.weight = 1;
	}

	PSTAT : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h114 };
		option.weight = 1;
	}
endgroup
	function new(string name = "DWC_ddrctl_map_REGB_ARB_PORT0");
		super.new(name, build_coverage(UVM_CVR_ADDR_MAP));
		add_coverage(build_coverage(UVM_CVR_ADDR_MAP));
		if (has_coverage(UVM_CVR_ADDR_MAP))
			cg_addr = new("cg_addr");
	endfunction: new

   virtual function void build();
      this.default_map = create_map("", 0, 4, UVM_LITTLE_ENDIAN, 0);
      this.PCCFG = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCCFG::type_id::create("PCCFG",,get_full_name());
      if(this.PCCFG.has_coverage(UVM_CVR_REG_BITS))
      	this.PCCFG.cg_bits.option.name = {get_name(), ".", "PCCFG_bits"};
      this.PCCFG.configure(this, null, "");
      this.PCCFG.build();
	  uvm_resource_db#(string)::set({"REG::", PCCFG.get_full_name()}, "accessType", "NONSECURE", this);
         this.PCCFG.add_hdl_path('{
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_go2critical_en", 0, 1},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_pagematch_limit", 4, 1}
         });
      this.default_map.add_reg(this.PCCFG, `UVM_REG_ADDR_WIDTH'h0, "RW", 0);
		this.PCCFG_go2critical_en = this.PCCFG.go2critical_en;
		this.go2critical_en = this.PCCFG.go2critical_en;
		this.PCCFG_pagematch_limit = this.PCCFG.pagematch_limit;
		this.pagematch_limit = this.PCCFG.pagematch_limit;
      this.PCFGR = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGR::type_id::create("PCFGR",,get_full_name());
      if(this.PCFGR.has_coverage(UVM_CVR_REG_BITS))
      	this.PCFGR.cg_bits.option.name = {get_name(), ".", "PCFGR_bits"};
      this.PCFGR.configure(this, null, "");
      this.PCFGR.build();
	  uvm_resource_db#(string)::set({"REG::", PCFGR.get_full_name()}, "accessType", "NONSECURE", this);
         this.PCFGR.add_hdl_path('{
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rd_port_priority", 0, 10},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rd_port_aging_en", 12, 1},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rd_port_urgent_en", 13, 1},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rd_port_pagematch_en", 14, 1},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rrb_lock_threshold", 20, 4}
         });
      this.default_map.add_reg(this.PCFGR, `UVM_REG_ADDR_WIDTH'h4, "RW", 0);
		this.PCFGR_rd_port_priority = this.PCFGR.rd_port_priority;
		this.rd_port_priority = this.PCFGR.rd_port_priority;
		this.PCFGR_rd_port_aging_en = this.PCFGR.rd_port_aging_en;
		this.rd_port_aging_en = this.PCFGR.rd_port_aging_en;
		this.PCFGR_rd_port_urgent_en = this.PCFGR.rd_port_urgent_en;
		this.rd_port_urgent_en = this.PCFGR.rd_port_urgent_en;
		this.PCFGR_rd_port_pagematch_en = this.PCFGR.rd_port_pagematch_en;
		this.rd_port_pagematch_en = this.PCFGR.rd_port_pagematch_en;
		this.PCFGR_rrb_lock_threshold = this.PCFGR.rrb_lock_threshold;
		this.rrb_lock_threshold = this.PCFGR.rrb_lock_threshold;
      this.PCFGW = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGW::type_id::create("PCFGW",,get_full_name());
      if(this.PCFGW.has_coverage(UVM_CVR_REG_BITS))
      	this.PCFGW.cg_bits.option.name = {get_name(), ".", "PCFGW_bits"};
      this.PCFGW.configure(this, null, "");
      this.PCFGW.build();
	  uvm_resource_db#(string)::set({"REG::", PCFGW.get_full_name()}, "accessType", "NONSECURE", this);
         this.PCFGW.add_hdl_path('{
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wr_port_priority", 0, 10},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wr_port_aging_en", 12, 1},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wr_port_urgent_en", 13, 1},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wr_port_pagematch_en", 14, 1}
         });
      this.default_map.add_reg(this.PCFGW, `UVM_REG_ADDR_WIDTH'h8, "RW", 0);
		this.PCFGW_wr_port_priority = this.PCFGW.wr_port_priority;
		this.wr_port_priority = this.PCFGW.wr_port_priority;
		this.PCFGW_wr_port_aging_en = this.PCFGW.wr_port_aging_en;
		this.wr_port_aging_en = this.PCFGW.wr_port_aging_en;
		this.PCFGW_wr_port_urgent_en = this.PCFGW.wr_port_urgent_en;
		this.wr_port_urgent_en = this.PCFGW.wr_port_urgent_en;
		this.PCFGW_wr_port_pagematch_en = this.PCFGW.wr_port_pagematch_en;
		this.wr_port_pagematch_en = this.PCFGW.wr_port_pagematch_en;
      this.PCTRL = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCTRL::type_id::create("PCTRL",,get_full_name());
      if(this.PCTRL.has_coverage(UVM_CVR_REG_BITS))
      	this.PCTRL.cg_bits.option.name = {get_name(), ".", "PCTRL_bits"};
      this.PCTRL.configure(this, null, "");
      this.PCTRL.build();
	  uvm_resource_db#(string)::set({"REG::", PCTRL.get_full_name()}, "accessType", "NONSECURE", this);
         this.PCTRL.add_hdl_path('{
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_port_en", 0, 1}
         });
      this.default_map.add_reg(this.PCTRL, `UVM_REG_ADDR_WIDTH'h90, "RW", 0);
		this.PCTRL_port_en = this.PCTRL.port_en;
		this.port_en = this.PCTRL.port_en;
      this.PCFGQOS0 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS0::type_id::create("PCFGQOS0",,get_full_name());
      if(this.PCFGQOS0.has_coverage(UVM_CVR_REG_BITS))
      	this.PCFGQOS0.cg_bits.option.name = {get_name(), ".", "PCFGQOS0_bits"};
      this.PCFGQOS0.configure(this, null, "");
      this.PCFGQOS0.build();
	  uvm_resource_db#(string)::set({"REG::", PCFGQOS0.get_full_name()}, "accessType", "NONSECURE", this);
         this.PCFGQOS0.add_hdl_path('{
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rqos_map_level1", 0, 4},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rqos_map_level2", 8, 4},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rqos_map_region0", 16, 2},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rqos_map_region1", 20, 2},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rqos_map_region2", 24, 2}
         });
      this.default_map.add_reg(this.PCFGQOS0, `UVM_REG_ADDR_WIDTH'h94, "RW", 0);
		this.PCFGQOS0_rqos_map_level1 = this.PCFGQOS0.rqos_map_level1;
		this.rqos_map_level1 = this.PCFGQOS0.rqos_map_level1;
		this.PCFGQOS0_rqos_map_level2 = this.PCFGQOS0.rqos_map_level2;
		this.rqos_map_level2 = this.PCFGQOS0.rqos_map_level2;
		this.PCFGQOS0_rqos_map_region0 = this.PCFGQOS0.rqos_map_region0;
		this.rqos_map_region0 = this.PCFGQOS0.rqos_map_region0;
		this.PCFGQOS0_rqos_map_region1 = this.PCFGQOS0.rqos_map_region1;
		this.rqos_map_region1 = this.PCFGQOS0.rqos_map_region1;
		this.PCFGQOS0_rqos_map_region2 = this.PCFGQOS0.rqos_map_region2;
		this.rqos_map_region2 = this.PCFGQOS0.rqos_map_region2;
      this.PCFGQOS1 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGQOS1::type_id::create("PCFGQOS1",,get_full_name());
      if(this.PCFGQOS1.has_coverage(UVM_CVR_REG_BITS))
      	this.PCFGQOS1.cg_bits.option.name = {get_name(), ".", "PCFGQOS1_bits"};
      this.PCFGQOS1.configure(this, null, "");
      this.PCFGQOS1.build();
	  uvm_resource_db#(string)::set({"REG::", PCFGQOS1.get_full_name()}, "accessType", "NONSECURE", this);
         this.PCFGQOS1.add_hdl_path('{
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rqos_map_timeoutb", 0, 11},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_rqos_map_timeoutr", 16, 11}
         });
      this.default_map.add_reg(this.PCFGQOS1, `UVM_REG_ADDR_WIDTH'h98, "RW", 0);
		this.PCFGQOS1_rqos_map_timeoutb = this.PCFGQOS1.rqos_map_timeoutb;
		this.rqos_map_timeoutb = this.PCFGQOS1.rqos_map_timeoutb;
		this.PCFGQOS1_rqos_map_timeoutr = this.PCFGQOS1.rqos_map_timeoutr;
		this.rqos_map_timeoutr = this.PCFGQOS1.rqos_map_timeoutr;
      this.PCFGWQOS0 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS0::type_id::create("PCFGWQOS0",,get_full_name());
      if(this.PCFGWQOS0.has_coverage(UVM_CVR_REG_BITS))
      	this.PCFGWQOS0.cg_bits.option.name = {get_name(), ".", "PCFGWQOS0_bits"};
      this.PCFGWQOS0.configure(this, null, "");
      this.PCFGWQOS0.build();
	  uvm_resource_db#(string)::set({"REG::", PCFGWQOS0.get_full_name()}, "accessType", "NONSECURE", this);
         this.PCFGWQOS0.add_hdl_path('{
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wqos_map_level1", 0, 4},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wqos_map_level2", 8, 4},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wqos_map_region0", 16, 2},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wqos_map_region1", 20, 2},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wqos_map_region2", 24, 2}
         });
      this.default_map.add_reg(this.PCFGWQOS0, `UVM_REG_ADDR_WIDTH'h9C, "RW", 0);
		this.PCFGWQOS0_wqos_map_level1 = this.PCFGWQOS0.wqos_map_level1;
		this.wqos_map_level1 = this.PCFGWQOS0.wqos_map_level1;
		this.PCFGWQOS0_wqos_map_level2 = this.PCFGWQOS0.wqos_map_level2;
		this.wqos_map_level2 = this.PCFGWQOS0.wqos_map_level2;
		this.PCFGWQOS0_wqos_map_region0 = this.PCFGWQOS0.wqos_map_region0;
		this.wqos_map_region0 = this.PCFGWQOS0.wqos_map_region0;
		this.PCFGWQOS0_wqos_map_region1 = this.PCFGWQOS0.wqos_map_region1;
		this.wqos_map_region1 = this.PCFGWQOS0.wqos_map_region1;
		this.PCFGWQOS0_wqos_map_region2 = this.PCFGWQOS0.wqos_map_region2;
		this.wqos_map_region2 = this.PCFGWQOS0.wqos_map_region2;
      this.PCFGWQOS1 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PCFGWQOS1::type_id::create("PCFGWQOS1",,get_full_name());
      if(this.PCFGWQOS1.has_coverage(UVM_CVR_REG_BITS))
      	this.PCFGWQOS1.cg_bits.option.name = {get_name(), ".", "PCFGWQOS1_bits"};
      this.PCFGWQOS1.configure(this, null, "");
      this.PCFGWQOS1.build();
	  uvm_resource_db#(string)::set({"REG::", PCFGWQOS1.get_full_name()}, "accessType", "NONSECURE", this);
         this.PCFGWQOS1.add_hdl_path('{
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wqos_map_timeout1", 0, 11},
            '{"U_apb_slvtop.slvif.cfgs_ff_regb_arb_port0_wqos_map_timeout2", 16, 11}
         });
      this.default_map.add_reg(this.PCFGWQOS1, `UVM_REG_ADDR_WIDTH'hA0, "RW", 0);
		this.PCFGWQOS1_wqos_map_timeout1 = this.PCFGWQOS1.wqos_map_timeout1;
		this.wqos_map_timeout1 = this.PCFGWQOS1.wqos_map_timeout1;
		this.PCFGWQOS1_wqos_map_timeout2 = this.PCFGWQOS1.wqos_map_timeout2;
		this.wqos_map_timeout2 = this.PCFGWQOS1.wqos_map_timeout2;
      this.SBRCTL = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRCTL::type_id::create("SBRCTL",,get_full_name());
      if(this.SBRCTL.has_coverage(UVM_CVR_REG_BITS))
      	this.SBRCTL.cg_bits.option.name = {get_name(), ".", "SBRCTL_bits"};
      this.SBRCTL.configure(this, null, "");
      this.SBRCTL.build();
	  uvm_resource_db#(string)::set({"REG::", SBRCTL.get_full_name()}, "accessType", "NONSECURE", this);
         this.SBRCTL.add_hdl_path('{
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_scrub_en", 0, 1},
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_scrub_during_lowpower", 1, 1},
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_scrub_burst_length_nm", 4, 3},
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_scrub_interval", 8, 13},
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_scrub_cmd_type", 24, 2},
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_scrub_burst_length_lp", 28, 3}
         });
      this.default_map.add_reg(this.SBRCTL, `UVM_REG_ADDR_WIDTH'hE0, "RW", 0);
		this.SBRCTL_scrub_en = this.SBRCTL.scrub_en;
		this.scrub_en = this.SBRCTL.scrub_en;
		this.SBRCTL_scrub_during_lowpower = this.SBRCTL.scrub_during_lowpower;
		this.scrub_during_lowpower = this.SBRCTL.scrub_during_lowpower;
		this.SBRCTL_scrub_burst_length_nm = this.SBRCTL.scrub_burst_length_nm;
		this.scrub_burst_length_nm = this.SBRCTL.scrub_burst_length_nm;
		this.SBRCTL_scrub_interval = this.SBRCTL.scrub_interval;
		this.scrub_interval = this.SBRCTL.scrub_interval;
		this.SBRCTL_scrub_cmd_type = this.SBRCTL.scrub_cmd_type;
		this.scrub_cmd_type = this.SBRCTL.scrub_cmd_type;
		this.SBRCTL_scrub_burst_length_lp = this.SBRCTL.scrub_burst_length_lp;
		this.scrub_burst_length_lp = this.SBRCTL.scrub_burst_length_lp;
      this.SBRSTAT = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTAT::type_id::create("SBRSTAT",,get_full_name());
      if(this.SBRSTAT.has_coverage(UVM_CVR_REG_BITS))
      	this.SBRSTAT.cg_bits.option.name = {get_name(), ".", "SBRSTAT_bits"};
      this.SBRSTAT.configure(this, null, "");
      this.SBRSTAT.build();
	  uvm_resource_db#(string)::set({"REG::", SBRSTAT.get_full_name()}, "accessType", "NONSECURE", this);
         this.SBRSTAT.add_hdl_path('{
            '{"arb_reg_scrub_busy", 0, 1},
            '{"arb_reg_scrub_done", 1, 1}
         });
      this.default_map.add_reg(this.SBRSTAT, `UVM_REG_ADDR_WIDTH'hE4, "RO", 0);
		this.SBRSTAT_scrub_busy = this.SBRSTAT.scrub_busy;
		this.scrub_busy = this.SBRSTAT.scrub_busy;
		this.SBRSTAT_scrub_done = this.SBRSTAT.scrub_done;
		this.scrub_done = this.SBRSTAT.scrub_done;
      this.SBRWDATA0 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRWDATA0::type_id::create("SBRWDATA0",,get_full_name());
      if(this.SBRWDATA0.has_coverage(UVM_CVR_REG_BITS))
      	this.SBRWDATA0.cg_bits.option.name = {get_name(), ".", "SBRWDATA0_bits"};
      this.SBRWDATA0.configure(this, null, "");
      this.SBRWDATA0.build();
	  uvm_resource_db#(string)::set({"REG::", SBRWDATA0.get_full_name()}, "accessType", "NONSECURE", this);
         this.SBRWDATA0.add_hdl_path('{
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_scrub_pattern0", 0, 32}
         });
      this.default_map.add_reg(this.SBRWDATA0, `UVM_REG_ADDR_WIDTH'hE8, "RW", 0);
		this.SBRWDATA0_scrub_pattern0 = this.SBRWDATA0.scrub_pattern0;
		this.scrub_pattern0 = this.SBRWDATA0.scrub_pattern0;
      this.SBRSTART0 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART0::type_id::create("SBRSTART0",,get_full_name());
      if(this.SBRSTART0.has_coverage(UVM_CVR_REG_BITS))
      	this.SBRSTART0.cg_bits.option.name = {get_name(), ".", "SBRSTART0_bits"};
      this.SBRSTART0.configure(this, null, "");
      this.SBRSTART0.build();
	  uvm_resource_db#(string)::set({"REG::", SBRSTART0.get_full_name()}, "accessType", "NONSECURE", this);
         this.SBRSTART0.add_hdl_path('{
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_sbr_address_start_mask_0", 0, 32}
         });
      this.default_map.add_reg(this.SBRSTART0, `UVM_REG_ADDR_WIDTH'hF0, "RW", 0);
		this.SBRSTART0_sbr_address_start_mask_0 = this.SBRSTART0.sbr_address_start_mask_0;
		this.sbr_address_start_mask_0 = this.SBRSTART0.sbr_address_start_mask_0;
      this.SBRSTART1 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRSTART1::type_id::create("SBRSTART1",,get_full_name());
      if(this.SBRSTART1.has_coverage(UVM_CVR_REG_BITS))
      	this.SBRSTART1.cg_bits.option.name = {get_name(), ".", "SBRSTART1_bits"};
      this.SBRSTART1.configure(this, null, "");
      this.SBRSTART1.build();
	  uvm_resource_db#(string)::set({"REG::", SBRSTART1.get_full_name()}, "accessType", "NONSECURE", this);
         this.SBRSTART1.add_hdl_path('{
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_sbr_address_start_mask_1", 0, 8}
         });
      this.default_map.add_reg(this.SBRSTART1, `UVM_REG_ADDR_WIDTH'hF4, "RW", 0);
		this.SBRSTART1_sbr_address_start_mask_1 = this.SBRSTART1.sbr_address_start_mask_1;
		this.sbr_address_start_mask_1 = this.SBRSTART1.sbr_address_start_mask_1;
      this.SBRRANGE0 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE0::type_id::create("SBRRANGE0",,get_full_name());
      if(this.SBRRANGE0.has_coverage(UVM_CVR_REG_BITS))
      	this.SBRRANGE0.cg_bits.option.name = {get_name(), ".", "SBRRANGE0_bits"};
      this.SBRRANGE0.configure(this, null, "");
      this.SBRRANGE0.build();
	  uvm_resource_db#(string)::set({"REG::", SBRRANGE0.get_full_name()}, "accessType", "NONSECURE", this);
         this.SBRRANGE0.add_hdl_path('{
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_sbr_address_range_mask_0", 0, 32}
         });
      this.default_map.add_reg(this.SBRRANGE0, `UVM_REG_ADDR_WIDTH'hF8, "RW", 0);
		this.SBRRANGE0_sbr_address_range_mask_0 = this.SBRRANGE0.sbr_address_range_mask_0;
		this.sbr_address_range_mask_0 = this.SBRRANGE0.sbr_address_range_mask_0;
      this.SBRRANGE1 = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_SBRRANGE1::type_id::create("SBRRANGE1",,get_full_name());
      if(this.SBRRANGE1.has_coverage(UVM_CVR_REG_BITS))
      	this.SBRRANGE1.cg_bits.option.name = {get_name(), ".", "SBRRANGE1_bits"};
      this.SBRRANGE1.configure(this, null, "");
      this.SBRRANGE1.build();
	  uvm_resource_db#(string)::set({"REG::", SBRRANGE1.get_full_name()}, "accessType", "NONSECURE", this);
         this.SBRRANGE1.add_hdl_path('{
            '{"U_apb_slvtop.slvif.ff_regb_arb_port0_sbr_address_range_mask_1", 0, 8}
         });
      this.default_map.add_reg(this.SBRRANGE1, `UVM_REG_ADDR_WIDTH'hFC, "RW", 0);
		this.SBRRANGE1_sbr_address_range_mask_1 = this.SBRRANGE1.sbr_address_range_mask_1;
		this.sbr_address_range_mask_1 = this.SBRRANGE1.sbr_address_range_mask_1;
      this.PSTAT = ral_reg_DWC_ddrctl_map_REGB_ARB_PORT0_PSTAT::type_id::create("PSTAT",,get_full_name());
      if(this.PSTAT.has_coverage(UVM_CVR_REG_BITS))
      	this.PSTAT.cg_bits.option.name = {get_name(), ".", "PSTAT_bits"};
      this.PSTAT.configure(this, null, "");
      this.PSTAT.build();
	  uvm_resource_db#(string)::set({"REG::", PSTAT.get_full_name()}, "accessType", "NONSECURE", this);
         this.PSTAT.add_hdl_path('{
            '{"arb_reg_rd_port_busy_0", 0, 1},
            '{"arb_reg_wr_port_busy_0", 16, 1}
         });
      this.default_map.add_reg(this.PSTAT, `UVM_REG_ADDR_WIDTH'h114, "RO", 0);
		this.PSTAT_rd_port_busy_0 = this.PSTAT.rd_port_busy_0;
		this.rd_port_busy_0 = this.PSTAT.rd_port_busy_0;
		this.PSTAT_wr_port_busy_0 = this.PSTAT.wr_port_busy_0;
		this.wr_port_busy_0 = this.PSTAT.wr_port_busy_0;
   endfunction : build

	`uvm_object_utils(ral_block_DWC_ddrctl_map_REGB_ARB_PORT0)


function void sample(uvm_reg_addr_t offset,
                     bit            is_read,
                     uvm_reg_map    map);
  if (get_coverage(UVM_CVR_ADDR_MAP)) begin
    m_offset = offset;
    cg_addr.sample();
  end
endfunction
endclass : ral_block_DWC_ddrctl_map_REGB_ARB_PORT0


endpackage
`endif
