// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_h_north
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_h_north_p (
  input logic [7:0] i_aic_4_init_tok_ocpl_s_maddr,
  input logic i_aic_4_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_4_init_tok_ocpl_s_mdata,
  output logic  o_aic_4_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_4_pwr_tok_idle_val,
  output logic  o_aic_4_pwr_tok_idle_ack,
  input logic  i_aic_4_pwr_tok_idle_req,
  output logic [7:0] o_aic_4_targ_tok_ocpl_m_maddr,
  output logic o_aic_4_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_4_targ_tok_ocpl_m_mdata,
  input logic  i_aic_4_targ_tok_ocpl_m_scmdaccept,
  input logic [7:0] i_aic_5_init_tok_ocpl_s_maddr,
  input logic i_aic_5_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_5_init_tok_ocpl_s_mdata,
  output logic  o_aic_5_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_5_pwr_tok_idle_val,
  output logic  o_aic_5_pwr_tok_idle_ack,
  input logic  i_aic_5_pwr_tok_idle_req,
  output logic [7:0] o_aic_5_targ_tok_ocpl_m_maddr,
  output logic o_aic_5_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_5_targ_tok_ocpl_m_mdata,
  input logic  i_aic_5_targ_tok_ocpl_m_scmdaccept,
  input logic [7:0] i_aic_6_init_tok_ocpl_s_maddr,
  input logic i_aic_6_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_6_init_tok_ocpl_s_mdata,
  output logic  o_aic_6_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_6_pwr_tok_idle_val,
  output logic  o_aic_6_pwr_tok_idle_ack,
  input logic  i_aic_6_pwr_tok_idle_req,
  output logic [7:0] o_aic_6_targ_tok_ocpl_m_maddr,
  output logic o_aic_6_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_6_targ_tok_ocpl_m_mdata,
  input logic  i_aic_6_targ_tok_ocpl_m_scmdaccept,
  input logic [7:0] i_aic_7_init_tok_ocpl_s_maddr,
  input logic i_aic_7_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_7_init_tok_ocpl_s_mdata,
  output logic  o_aic_7_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_7_pwr_tok_idle_val,
  output logic  o_aic_7_pwr_tok_idle_ack,
  input logic  i_aic_7_pwr_tok_idle_req,
  output logic [7:0] o_aic_7_targ_tok_ocpl_m_maddr,
  output logic o_aic_7_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_7_targ_tok_ocpl_m_mdata,
  input logic  i_aic_7_targ_tok_ocpl_m_scmdaccept,
  input logic [41:0] i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld,

    input  wire                                    i_aic_4_aon_clk,
    input  wire                                    i_aic_4_aon_rst_n,
    input  wire                                    i_aic_4_clk,
    input  wire                                    i_aic_4_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_4_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_4_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_4_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_4_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_4_init_ht_axi_s_arlen,
    input  logic                                   i_aic_4_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_4_init_ht_axi_s_arprot,
    output logic                                   o_aic_4_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_4_init_ht_axi_s_arsize,
    input  logic                                   i_aic_4_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_4_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_4_init_ht_axi_s_rid,
    output logic                                   o_aic_4_init_ht_axi_s_rlast,
    input  logic                                   i_aic_4_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_4_init_ht_axi_s_rresp,
    output logic                                   o_aic_4_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_4_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_4_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_4_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_4_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_4_init_ht_axi_s_awlen,
    input  logic                                   i_aic_4_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_4_init_ht_axi_s_awprot,
    output logic                                   o_aic_4_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_4_init_ht_axi_s_awsize,
    input  logic                                   i_aic_4_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_4_init_ht_axi_s_bid,
    input  logic                                   i_aic_4_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_4_init_ht_axi_s_bresp,
    output logic                                   o_aic_4_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_4_init_ht_axi_s_wdata,
    input  logic                                   i_aic_4_init_ht_axi_s_wlast,
    output logic                                   o_aic_4_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_4_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_4_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_4_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_4_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_4_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_4_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_4_init_lt_axi_s_arlen,
    input  logic                                   i_aic_4_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_4_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_4_init_lt_axi_s_arqos,
    output logic                                   o_aic_4_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_4_init_lt_axi_s_arsize,
    input  logic                                   i_aic_4_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_4_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_4_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_4_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_4_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_4_init_lt_axi_s_awlen,
    input  logic                                   i_aic_4_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_4_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_4_init_lt_axi_s_awqos,
    output logic                                   o_aic_4_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_4_init_lt_axi_s_awsize,
    input  logic                                   i_aic_4_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_4_init_lt_axi_s_bid,
    input  logic                                   i_aic_4_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_4_init_lt_axi_s_bresp,
    output logic                                   o_aic_4_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_4_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_4_init_lt_axi_s_rid,
    output logic                                   o_aic_4_init_lt_axi_s_rlast,
    input  logic                                   i_aic_4_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_4_init_lt_axi_s_rresp,
    output logic                                   o_aic_4_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_4_init_lt_axi_s_wdata,
    input  logic                                   i_aic_4_init_lt_axi_s_wlast,
    output logic                                   o_aic_4_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_4_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_4_init_lt_axi_s_wvalid,
    output logic                                   o_aic_4_pwr_idle_val,
    output logic                                   o_aic_4_pwr_idle_ack,
    input  logic                                   i_aic_4_pwr_idle_req,
    input  wire                                    i_aic_4_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_4_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_4_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_4_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_4_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_4_targ_lt_axi_m_arlen,
    output logic                                   o_aic_4_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_4_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_4_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_4_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_4_targ_lt_axi_m_arsize,
    output logic                                   o_aic_4_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_4_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_4_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_4_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_4_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_4_targ_lt_axi_m_awlen,
    output logic                                   o_aic_4_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_4_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_4_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_4_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_4_targ_lt_axi_m_awsize,
    output logic                                   o_aic_4_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_4_targ_lt_axi_m_bid,
    output logic                                   o_aic_4_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_4_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_4_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_4_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_4_targ_lt_axi_m_rid,
    input  logic                                   i_aic_4_targ_lt_axi_m_rlast,
    output logic                                   o_aic_4_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_4_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_4_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_4_targ_lt_axi_m_wdata,
    output logic                                   o_aic_4_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_4_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_4_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_4_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_4_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_4_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_4_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_4_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_4_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_4_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_4_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_4_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_4_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_4_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_5_aon_clk,
    input  wire                                    i_aic_5_aon_rst_n,
    input  wire                                    i_aic_5_clk,
    input  wire                                    i_aic_5_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_5_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_5_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_5_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_5_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_5_init_ht_axi_s_arlen,
    input  logic                                   i_aic_5_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_5_init_ht_axi_s_arprot,
    output logic                                   o_aic_5_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_5_init_ht_axi_s_arsize,
    input  logic                                   i_aic_5_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_5_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_5_init_ht_axi_s_rid,
    output logic                                   o_aic_5_init_ht_axi_s_rlast,
    input  logic                                   i_aic_5_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_5_init_ht_axi_s_rresp,
    output logic                                   o_aic_5_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_5_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_5_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_5_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_5_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_5_init_ht_axi_s_awlen,
    input  logic                                   i_aic_5_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_5_init_ht_axi_s_awprot,
    output logic                                   o_aic_5_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_5_init_ht_axi_s_awsize,
    input  logic                                   i_aic_5_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_5_init_ht_axi_s_bid,
    input  logic                                   i_aic_5_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_5_init_ht_axi_s_bresp,
    output logic                                   o_aic_5_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_5_init_ht_axi_s_wdata,
    input  logic                                   i_aic_5_init_ht_axi_s_wlast,
    output logic                                   o_aic_5_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_5_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_5_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_5_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_5_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_5_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_5_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_5_init_lt_axi_s_arlen,
    input  logic                                   i_aic_5_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_5_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_5_init_lt_axi_s_arqos,
    output logic                                   o_aic_5_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_5_init_lt_axi_s_arsize,
    input  logic                                   i_aic_5_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_5_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_5_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_5_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_5_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_5_init_lt_axi_s_awlen,
    input  logic                                   i_aic_5_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_5_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_5_init_lt_axi_s_awqos,
    output logic                                   o_aic_5_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_5_init_lt_axi_s_awsize,
    input  logic                                   i_aic_5_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_5_init_lt_axi_s_bid,
    input  logic                                   i_aic_5_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_5_init_lt_axi_s_bresp,
    output logic                                   o_aic_5_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_5_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_5_init_lt_axi_s_rid,
    output logic                                   o_aic_5_init_lt_axi_s_rlast,
    input  logic                                   i_aic_5_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_5_init_lt_axi_s_rresp,
    output logic                                   o_aic_5_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_5_init_lt_axi_s_wdata,
    input  logic                                   i_aic_5_init_lt_axi_s_wlast,
    output logic                                   o_aic_5_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_5_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_5_init_lt_axi_s_wvalid,
    output logic                                   o_aic_5_pwr_idle_val,
    output logic                                   o_aic_5_pwr_idle_ack,
    input  logic                                   i_aic_5_pwr_idle_req,
    input  wire                                    i_aic_5_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_5_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_5_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_5_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_5_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_5_targ_lt_axi_m_arlen,
    output logic                                   o_aic_5_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_5_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_5_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_5_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_5_targ_lt_axi_m_arsize,
    output logic                                   o_aic_5_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_5_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_5_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_5_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_5_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_5_targ_lt_axi_m_awlen,
    output logic                                   o_aic_5_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_5_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_5_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_5_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_5_targ_lt_axi_m_awsize,
    output logic                                   o_aic_5_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_5_targ_lt_axi_m_bid,
    output logic                                   o_aic_5_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_5_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_5_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_5_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_5_targ_lt_axi_m_rid,
    input  logic                                   i_aic_5_targ_lt_axi_m_rlast,
    output logic                                   o_aic_5_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_5_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_5_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_5_targ_lt_axi_m_wdata,
    output logic                                   o_aic_5_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_5_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_5_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_5_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_5_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_5_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_5_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_5_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_5_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_5_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_5_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_5_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_5_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_5_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_6_aon_clk,
    input  wire                                    i_aic_6_aon_rst_n,
    input  wire                                    i_aic_6_clk,
    input  wire                                    i_aic_6_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_6_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_6_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_6_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_6_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_6_init_ht_axi_s_arlen,
    input  logic                                   i_aic_6_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_6_init_ht_axi_s_arprot,
    output logic                                   o_aic_6_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_6_init_ht_axi_s_arsize,
    input  logic                                   i_aic_6_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_6_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_6_init_ht_axi_s_rid,
    output logic                                   o_aic_6_init_ht_axi_s_rlast,
    input  logic                                   i_aic_6_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_6_init_ht_axi_s_rresp,
    output logic                                   o_aic_6_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_6_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_6_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_6_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_6_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_6_init_ht_axi_s_awlen,
    input  logic                                   i_aic_6_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_6_init_ht_axi_s_awprot,
    output logic                                   o_aic_6_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_6_init_ht_axi_s_awsize,
    input  logic                                   i_aic_6_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_6_init_ht_axi_s_bid,
    input  logic                                   i_aic_6_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_6_init_ht_axi_s_bresp,
    output logic                                   o_aic_6_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_6_init_ht_axi_s_wdata,
    input  logic                                   i_aic_6_init_ht_axi_s_wlast,
    output logic                                   o_aic_6_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_6_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_6_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_6_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_6_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_6_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_6_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_6_init_lt_axi_s_arlen,
    input  logic                                   i_aic_6_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_6_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_6_init_lt_axi_s_arqos,
    output logic                                   o_aic_6_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_6_init_lt_axi_s_arsize,
    input  logic                                   i_aic_6_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_6_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_6_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_6_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_6_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_6_init_lt_axi_s_awlen,
    input  logic                                   i_aic_6_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_6_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_6_init_lt_axi_s_awqos,
    output logic                                   o_aic_6_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_6_init_lt_axi_s_awsize,
    input  logic                                   i_aic_6_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_6_init_lt_axi_s_bid,
    input  logic                                   i_aic_6_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_6_init_lt_axi_s_bresp,
    output logic                                   o_aic_6_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_6_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_6_init_lt_axi_s_rid,
    output logic                                   o_aic_6_init_lt_axi_s_rlast,
    input  logic                                   i_aic_6_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_6_init_lt_axi_s_rresp,
    output logic                                   o_aic_6_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_6_init_lt_axi_s_wdata,
    input  logic                                   i_aic_6_init_lt_axi_s_wlast,
    output logic                                   o_aic_6_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_6_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_6_init_lt_axi_s_wvalid,
    output logic                                   o_aic_6_pwr_idle_val,
    output logic                                   o_aic_6_pwr_idle_ack,
    input  logic                                   i_aic_6_pwr_idle_req,
    input  wire                                    i_aic_6_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_6_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_6_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_6_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_6_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_6_targ_lt_axi_m_arlen,
    output logic                                   o_aic_6_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_6_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_6_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_6_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_6_targ_lt_axi_m_arsize,
    output logic                                   o_aic_6_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_6_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_6_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_6_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_6_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_6_targ_lt_axi_m_awlen,
    output logic                                   o_aic_6_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_6_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_6_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_6_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_6_targ_lt_axi_m_awsize,
    output logic                                   o_aic_6_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_6_targ_lt_axi_m_bid,
    output logic                                   o_aic_6_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_6_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_6_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_6_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_6_targ_lt_axi_m_rid,
    input  logic                                   i_aic_6_targ_lt_axi_m_rlast,
    output logic                                   o_aic_6_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_6_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_6_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_6_targ_lt_axi_m_wdata,
    output logic                                   o_aic_6_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_6_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_6_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_6_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_6_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_6_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_6_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_6_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_6_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_6_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_6_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_6_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_6_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_6_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_aic_7_aon_clk,
    input  wire                                    i_aic_7_aon_rst_n,
    input  wire                                    i_aic_7_clk,
    input  wire                                    i_aic_7_clken,
    input  chip_pkg::chip_axi_addr_t               i_aic_7_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_7_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_7_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_7_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_7_init_ht_axi_s_arlen,
    input  logic                                   i_aic_7_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_7_init_ht_axi_s_arprot,
    output logic                                   o_aic_7_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_7_init_ht_axi_s_arsize,
    input  logic                                   i_aic_7_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t            o_aic_7_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_7_init_ht_axi_s_rid,
    output logic                                   o_aic_7_init_ht_axi_s_rlast,
    input  logic                                   i_aic_7_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_7_init_ht_axi_s_rresp,
    output logic                                   o_aic_7_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_7_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_7_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_7_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t   i_aic_7_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_7_init_ht_axi_s_awlen,
    input  logic                                   i_aic_7_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_7_init_ht_axi_s_awprot,
    output logic                                   o_aic_7_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_7_init_ht_axi_s_awsize,
    input  logic                                   i_aic_7_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t   o_aic_7_init_ht_axi_s_bid,
    input  logic                                   i_aic_7_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_7_init_ht_axi_s_bresp,
    output logic                                   o_aic_7_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_aic_7_init_ht_axi_s_wdata,
    input  logic                                   i_aic_7_init_ht_axi_s_wlast,
    output logic                                   o_aic_7_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t           i_aic_7_init_ht_axi_s_wstrb,
    input  logic                                   i_aic_7_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_7_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                    i_aic_7_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                    i_aic_7_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_7_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                      i_aic_7_init_lt_axi_s_arlen,
    input  logic                                   i_aic_7_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                     i_aic_7_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                      i_aic_7_init_lt_axi_s_arqos,
    output logic                                   o_aic_7_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                     i_aic_7_init_lt_axi_s_arsize,
    input  logic                                   i_aic_7_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t               i_aic_7_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                    i_aic_7_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                    i_aic_7_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t   i_aic_7_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                      i_aic_7_init_lt_axi_s_awlen,
    input  logic                                   i_aic_7_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                     i_aic_7_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                      i_aic_7_init_lt_axi_s_awqos,
    output logic                                   o_aic_7_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                     i_aic_7_init_lt_axi_s_awsize,
    input  logic                                   i_aic_7_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_7_init_lt_axi_s_bid,
    input  logic                                   i_aic_7_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                     o_aic_7_init_lt_axi_s_bresp,
    output logic                                   o_aic_7_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_7_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t   o_aic_7_init_lt_axi_s_rid,
    output logic                                   o_aic_7_init_lt_axi_s_rlast,
    input  logic                                   i_aic_7_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                     o_aic_7_init_lt_axi_s_rresp,
    output logic                                   o_aic_7_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_7_init_lt_axi_s_wdata,
    input  logic                                   i_aic_7_init_lt_axi_s_wlast,
    output logic                                   o_aic_7_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t           i_aic_7_init_lt_axi_s_wstrb,
    input  logic                                   i_aic_7_init_lt_axi_s_wvalid,
    output logic                                   o_aic_7_pwr_idle_val,
    output logic                                   o_aic_7_pwr_idle_ack,
    input  logic                                   i_aic_7_pwr_idle_req,
    input  wire                                    i_aic_7_rst_n,
    output chip_pkg::chip_axi_addr_t               o_aic_7_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_aic_7_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_aic_7_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_7_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                      o_aic_7_targ_lt_axi_m_arlen,
    output logic                                   o_aic_7_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_aic_7_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                      o_aic_7_targ_lt_axi_m_arqos,
    input  logic                                   i_aic_7_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                     o_aic_7_targ_lt_axi_m_arsize,
    output logic                                   o_aic_7_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t               o_aic_7_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_aic_7_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_aic_7_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t   o_aic_7_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                      o_aic_7_targ_lt_axi_m_awlen,
    output logic                                   o_aic_7_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_aic_7_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                      o_aic_7_targ_lt_axi_m_awqos,
    input  logic                                   i_aic_7_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                     o_aic_7_targ_lt_axi_m_awsize,
    output logic                                   o_aic_7_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_7_targ_lt_axi_m_bid,
    output logic                                   o_aic_7_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_aic_7_targ_lt_axi_m_bresp,
    input  logic                                   i_aic_7_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t            i_aic_7_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t   i_aic_7_targ_lt_axi_m_rid,
    input  logic                                   i_aic_7_targ_lt_axi_m_rlast,
    output logic                                   o_aic_7_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_aic_7_targ_lt_axi_m_rresp,
    input  logic                                   i_aic_7_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t            o_aic_7_targ_lt_axi_m_wdata,
    output logic                                   o_aic_7_targ_lt_axi_m_wlast,
    input  logic                                   i_aic_7_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t           o_aic_7_targ_lt_axi_m_wstrb,
    output logic                                   o_aic_7_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_aic_7_targ_syscfg_apb_m_paddr,
    output logic                                   o_aic_7_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_aic_7_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_aic_7_targ_syscfg_apb_m_prdata,
    input  logic                                   i_aic_7_targ_syscfg_apb_m_pready,
    output logic                                   o_aic_7_targ_syscfg_apb_m_psel,
    input  logic                                   i_aic_7_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_aic_7_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_aic_7_targ_syscfg_apb_m_pwdata,
    output logic                                   o_aic_7_targ_syscfg_apb_m_pwrite,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld,
    input  logic [686:0]                           i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld,
    output logic [108:0]                           o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld,
    input  logic [146:0]                           i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld,
    output logic [686:0]                           o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld,
    input  logic [182:0]                           i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data,
    input  logic                                   i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head,
    output logic                                   o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy,
    input  logic                                   i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail,
    input  logic                                   i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld,
    output logic [182:0]                           o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data,
    output logic                                   o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head,
    input  logic                                   i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy,
    output logic                                   o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail,
    output logic                                   o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld,
    output logic [686:0]                           o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld,
    input  logic [108:0]                           i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld,
    output logic [146:0]                           o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld,
    input  logic [686:0]                           i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld,
    output logic [182:0]                           o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data,
    output logic                                   o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head,
    input  logic                                   i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy,
    output logic                                   o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail,
    output logic                                   o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld,
    input  logic [182:0]                           i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data,
    input  logic                                   i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head,
    output logic                                   o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy,
    input  logic                                   i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail,
    input  logic                                   i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld,
    input  wire                                    i_l2_4_aon_clk,
    input  wire                                    i_l2_4_aon_rst_n,
    input  wire                                    i_l2_4_clk,
    input  wire                                    i_l2_4_clken,
    output logic                                   o_l2_4_pwr_idle_val,
    output logic                                   o_l2_4_pwr_idle_ack,
    input  logic                                   i_l2_4_pwr_idle_req,
    input  wire                                    i_l2_4_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_4_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_4_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_4_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_4_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_4_targ_ht_axi_m_arlen,
    output logic                                   o_l2_4_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_4_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_4_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_4_targ_ht_axi_m_arsize,
    output logic                                   o_l2_4_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_4_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_4_targ_ht_axi_m_rid,
    input  logic                                   i_l2_4_targ_ht_axi_m_rlast,
    output logic                                   o_l2_4_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_4_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_4_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_4_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_4_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_4_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_4_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_4_targ_ht_axi_m_awlen,
    output logic                                   o_l2_4_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_4_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_4_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_4_targ_ht_axi_m_awsize,
    output logic                                   o_l2_4_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_4_targ_ht_axi_m_bid,
    output logic                                   o_l2_4_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_4_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_4_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_4_targ_ht_axi_m_wdata,
    output logic                                   o_l2_4_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_4_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_4_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_4_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_4_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_4_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_4_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_4_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_4_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_4_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_4_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_4_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_4_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_4_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_5_aon_clk,
    input  wire                                    i_l2_5_aon_rst_n,
    input  wire                                    i_l2_5_clk,
    input  wire                                    i_l2_5_clken,
    output logic                                   o_l2_5_pwr_idle_val,
    output logic                                   o_l2_5_pwr_idle_ack,
    input  logic                                   i_l2_5_pwr_idle_req,
    input  wire                                    i_l2_5_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_5_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_5_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_5_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_5_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_5_targ_ht_axi_m_arlen,
    output logic                                   o_l2_5_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_5_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_5_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_5_targ_ht_axi_m_arsize,
    output logic                                   o_l2_5_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_5_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_5_targ_ht_axi_m_rid,
    input  logic                                   i_l2_5_targ_ht_axi_m_rlast,
    output logic                                   o_l2_5_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_5_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_5_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_5_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_5_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_5_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_5_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_5_targ_ht_axi_m_awlen,
    output logic                                   o_l2_5_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_5_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_5_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_5_targ_ht_axi_m_awsize,
    output logic                                   o_l2_5_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_5_targ_ht_axi_m_bid,
    output logic                                   o_l2_5_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_5_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_5_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_5_targ_ht_axi_m_wdata,
    output logic                                   o_l2_5_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_5_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_5_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_5_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_5_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_5_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_5_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_5_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_5_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_5_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_5_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_5_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_5_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_5_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_6_aon_clk,
    input  wire                                    i_l2_6_aon_rst_n,
    input  wire                                    i_l2_6_clk,
    input  wire                                    i_l2_6_clken,
    output logic                                   o_l2_6_pwr_idle_val,
    output logic                                   o_l2_6_pwr_idle_ack,
    input  logic                                   i_l2_6_pwr_idle_req,
    input  wire                                    i_l2_6_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_6_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_6_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_6_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_6_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_6_targ_ht_axi_m_arlen,
    output logic                                   o_l2_6_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_6_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_6_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_6_targ_ht_axi_m_arsize,
    output logic                                   o_l2_6_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_6_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_6_targ_ht_axi_m_rid,
    input  logic                                   i_l2_6_targ_ht_axi_m_rlast,
    output logic                                   o_l2_6_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_6_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_6_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_6_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_6_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_6_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_6_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_6_targ_ht_axi_m_awlen,
    output logic                                   o_l2_6_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_6_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_6_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_6_targ_ht_axi_m_awsize,
    output logic                                   o_l2_6_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_6_targ_ht_axi_m_bid,
    output logic                                   o_l2_6_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_6_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_6_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_6_targ_ht_axi_m_wdata,
    output logic                                   o_l2_6_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_6_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_6_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_6_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_6_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_6_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_6_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_6_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_6_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_6_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_6_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_6_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_6_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_6_targ_syscfg_apb_m_pwrite,
    input  wire                                    i_l2_7_aon_clk,
    input  wire                                    i_l2_7_aon_rst_n,
    input  wire                                    i_l2_7_clk,
    input  wire                                    i_l2_7_clken,
    output logic                                   o_l2_7_pwr_idle_val,
    output logic                                   o_l2_7_pwr_idle_ack,
    input  logic                                   i_l2_7_pwr_idle_req,
    input  wire                                    i_l2_7_rst_n,
    output chip_pkg::chip_axi_addr_t               o_l2_7_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                    o_l2_7_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                    o_l2_7_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_7_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                      o_l2_7_targ_ht_axi_m_arlen,
    output logic                                   o_l2_7_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                     o_l2_7_targ_ht_axi_m_arprot,
    input  logic                                   i_l2_7_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                     o_l2_7_targ_ht_axi_m_arsize,
    output logic                                   o_l2_7_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t            i_l2_7_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_7_targ_ht_axi_m_rid,
    input  logic                                   i_l2_7_targ_ht_axi_m_rlast,
    output logic                                   o_l2_7_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                     i_l2_7_targ_ht_axi_m_rresp,
    input  logic                                   i_l2_7_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t               o_l2_7_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                    o_l2_7_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                    o_l2_7_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t           o_l2_7_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                      o_l2_7_targ_ht_axi_m_awlen,
    output logic                                   o_l2_7_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                     o_l2_7_targ_ht_axi_m_awprot,
    input  logic                                   i_l2_7_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                     o_l2_7_targ_ht_axi_m_awsize,
    output logic                                   o_l2_7_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t           i_l2_7_targ_ht_axi_m_bid,
    output logic                                   o_l2_7_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                     i_l2_7_targ_ht_axi_m_bresp,
    input  logic                                   i_l2_7_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t            o_l2_7_targ_ht_axi_m_wdata,
    output logic                                   o_l2_7_targ_ht_axi_m_wlast,
    input  logic                                   i_l2_7_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t           o_l2_7_targ_ht_axi_m_wstrb,
    output logic                                   o_l2_7_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t            o_l2_7_targ_syscfg_apb_m_paddr,
    output logic                                   o_l2_7_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                 o_l2_7_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t        i_l2_7_targ_syscfg_apb_m_prdata,
    input  logic                                   i_l2_7_targ_syscfg_apb_m_pready,
    output logic                                   o_l2_7_targ_syscfg_apb_m_psel,
    input  logic                                   i_l2_7_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t        o_l2_7_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t        o_l2_7_targ_syscfg_apb_m_pwdata,
    output logic                                   o_l2_7_targ_syscfg_apb_m_pwrite,
    input  logic                                   i_l2_addr_mode_port_b0,
    input  logic                                   i_l2_addr_mode_port_b1,
    input  logic                                   i_l2_intr_mode_port_b0,
    input  logic                                   i_l2_intr_mode_port_b1,
    input  logic                                   i_lpddr_graph_addr_mode_port_b0,
    input  logic                                   i_lpddr_graph_addr_mode_port_b1,
    input  logic                                   i_lpddr_graph_intr_mode_port_b0,
    input  logic                                   i_lpddr_graph_intr_mode_port_b1,
    input  logic                                   i_lpddr_ppp_addr_mode_port_b0,
    input  logic                                   i_lpddr_ppp_addr_mode_port_b1,
    input  logic                                   i_lpddr_ppp_intr_mode_port_b0,
    input  logic                                   i_lpddr_ppp_intr_mode_port_b1,
    input  wire                                    i_noc_clk,
    input  wire                                    i_noc_rst_n,
    // DFT Interface
    input  wire           tck,
    input  wire           trst,
    input  logic          tms,
    input  logic          tdi,
    output logic          tdo_en,
    output logic          tdo,
    input  wire           test_clk,
    input  logic          test_mode,
    input  logic          edt_update,
    input  logic          scan_en,
    input  logic [30-1:0] scan_in,
    output logic [30-1:0] scan_out
);

logic [2:0] aic_4_targ_tok_ocpl_m_mcmd_ext;
assign o_aic_4_targ_tok_ocpl_m_mcmd = aic_4_targ_tok_ocpl_m_mcmd_ext[0];
logic [2:0] aic_5_targ_tok_ocpl_m_mcmd_ext;
assign o_aic_5_targ_tok_ocpl_m_mcmd = aic_5_targ_tok_ocpl_m_mcmd_ext[0];
logic [2:0] aic_6_targ_tok_ocpl_m_mcmd_ext;
assign o_aic_6_targ_tok_ocpl_m_mcmd = aic_6_targ_tok_ocpl_m_mcmd_ext[0];
logic [2:0] aic_7_targ_tok_ocpl_m_mcmd_ext;
assign o_aic_7_targ_tok_ocpl_m_mcmd = aic_7_targ_tok_ocpl_m_mcmd_ext[0];


    // -- Automatically-generated Reset Synchronizers -- //
    wire aic_4_aon_rst_n_synced;
    wire aic_5_aon_rst_n_synced;
    wire aic_6_aon_rst_n_synced;
    wire aic_7_aon_rst_n_synced;
    wire l2_4_aon_rst_n_synced;
    wire l2_5_aon_rst_n_synced;
    wire l2_6_aon_rst_n_synced;
    wire l2_7_aon_rst_n_synced;

    // AIC 4 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_aic_4_aon_rst_n_sync (
        .i_clk          (i_aic_4_aon_clk),
        .i_rst_n        (i_aic_4_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (aic_4_aon_rst_n_synced)
    );

    // AIC 5 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_aic_5_aon_rst_n_sync (
        .i_clk          (i_aic_5_aon_clk),
        .i_rst_n        (i_aic_5_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (aic_5_aon_rst_n_synced)
    );

    // AIC 6 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_aic_6_aon_rst_n_sync (
        .i_clk          (i_aic_6_aon_clk),
        .i_rst_n        (i_aic_6_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (aic_6_aon_rst_n_synced)
    );

    // AIC 7 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_aic_7_aon_rst_n_sync (
        .i_clk          (i_aic_7_aon_clk),
        .i_rst_n        (i_aic_7_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (aic_7_aon_rst_n_synced)
    );

    // L2 4 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_l2_4_aon_rst_n_sync (
        .i_clk          (i_l2_4_aon_clk),
        .i_rst_n        (i_l2_4_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (l2_4_aon_rst_n_synced)
    );

    // L2 5 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_l2_5_aon_rst_n_sync (
        .i_clk          (i_l2_5_aon_clk),
        .i_rst_n        (i_l2_5_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (l2_5_aon_rst_n_synced)
    );

    // L2 6 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_l2_6_aon_rst_n_sync (
        .i_clk          (i_l2_6_aon_clk),
        .i_rst_n        (i_l2_6_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (l2_6_aon_rst_n_synced)
    );

    // L2 7 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_l2_7_aon_rst_n_sync (
        .i_clk          (i_l2_7_aon_clk),
        .i_rst_n        (i_l2_7_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (l2_7_aon_rst_n_synced)
    );

    noc_h_north u_noc_h_north (
    .i_aic_4_aon_clk(i_aic_4_aon_clk),
    .i_aic_4_aon_rst_n(aic_4_aon_rst_n_synced),
    .i_aic_4_clk(i_aic_4_clk),
    .i_aic_4_clken(i_aic_4_clken),
    .i_aic_4_init_ht_axi_s_araddr(i_aic_4_init_ht_axi_s_araddr),
    .i_aic_4_init_ht_axi_s_arburst(i_aic_4_init_ht_axi_s_arburst),
    .i_aic_4_init_ht_axi_s_arcache(i_aic_4_init_ht_axi_s_arcache),
    .i_aic_4_init_ht_axi_s_arid(i_aic_4_init_ht_axi_s_arid),
    .i_aic_4_init_ht_axi_s_arlen(i_aic_4_init_ht_axi_s_arlen),
    .i_aic_4_init_ht_axi_s_arlock(i_aic_4_init_ht_axi_s_arlock),
    .i_aic_4_init_ht_axi_s_arprot(i_aic_4_init_ht_axi_s_arprot),
    .o_aic_4_init_ht_axi_s_arready(o_aic_4_init_ht_axi_s_arready),
    .i_aic_4_init_ht_axi_s_arsize(i_aic_4_init_ht_axi_s_arsize),
    .i_aic_4_init_ht_axi_s_arvalid(i_aic_4_init_ht_axi_s_arvalid),
    .o_aic_4_init_ht_axi_s_rdata(o_aic_4_init_ht_axi_s_rdata),
    .o_aic_4_init_ht_axi_s_rid(o_aic_4_init_ht_axi_s_rid),
    .o_aic_4_init_ht_axi_s_rlast(o_aic_4_init_ht_axi_s_rlast),
    .i_aic_4_init_ht_axi_s_rready(i_aic_4_init_ht_axi_s_rready),
    .o_aic_4_init_ht_axi_s_rresp(o_aic_4_init_ht_axi_s_rresp),
    .o_aic_4_init_ht_axi_s_rvalid(o_aic_4_init_ht_axi_s_rvalid),
    .i_aic_4_init_ht_axi_s_awaddr(i_aic_4_init_ht_axi_s_awaddr),
    .i_aic_4_init_ht_axi_s_awburst(i_aic_4_init_ht_axi_s_awburst),
    .i_aic_4_init_ht_axi_s_awcache(i_aic_4_init_ht_axi_s_awcache),
    .i_aic_4_init_ht_axi_s_awid(i_aic_4_init_ht_axi_s_awid),
    .i_aic_4_init_ht_axi_s_awlen(i_aic_4_init_ht_axi_s_awlen),
    .i_aic_4_init_ht_axi_s_awlock(i_aic_4_init_ht_axi_s_awlock),
    .i_aic_4_init_ht_axi_s_awprot(i_aic_4_init_ht_axi_s_awprot),
    .o_aic_4_init_ht_axi_s_awready(o_aic_4_init_ht_axi_s_awready),
    .i_aic_4_init_ht_axi_s_awsize(i_aic_4_init_ht_axi_s_awsize),
    .i_aic_4_init_ht_axi_s_awvalid(i_aic_4_init_ht_axi_s_awvalid),
    .o_aic_4_init_ht_axi_s_bid(o_aic_4_init_ht_axi_s_bid),
    .i_aic_4_init_ht_axi_s_bready(i_aic_4_init_ht_axi_s_bready),
    .o_aic_4_init_ht_axi_s_bresp(o_aic_4_init_ht_axi_s_bresp),
    .o_aic_4_init_ht_axi_s_bvalid(o_aic_4_init_ht_axi_s_bvalid),
    .i_aic_4_init_ht_axi_s_wdata(i_aic_4_init_ht_axi_s_wdata),
    .i_aic_4_init_ht_axi_s_wlast(i_aic_4_init_ht_axi_s_wlast),
    .o_aic_4_init_ht_axi_s_wready(o_aic_4_init_ht_axi_s_wready),
    .i_aic_4_init_ht_axi_s_wstrb(i_aic_4_init_ht_axi_s_wstrb),
    .i_aic_4_init_ht_axi_s_wvalid(i_aic_4_init_ht_axi_s_wvalid),
    .i_aic_4_init_lt_axi_s_araddr(i_aic_4_init_lt_axi_s_araddr),
    .i_aic_4_init_lt_axi_s_arburst(i_aic_4_init_lt_axi_s_arburst),
    .i_aic_4_init_lt_axi_s_arcache(i_aic_4_init_lt_axi_s_arcache),
    .i_aic_4_init_lt_axi_s_arid(i_aic_4_init_lt_axi_s_arid),
    .i_aic_4_init_lt_axi_s_arlen(i_aic_4_init_lt_axi_s_arlen),
    .i_aic_4_init_lt_axi_s_arlock(i_aic_4_init_lt_axi_s_arlock),
    .i_aic_4_init_lt_axi_s_arprot(i_aic_4_init_lt_axi_s_arprot),
    .i_aic_4_init_lt_axi_s_arqos(i_aic_4_init_lt_axi_s_arqos),
    .o_aic_4_init_lt_axi_s_arready(o_aic_4_init_lt_axi_s_arready),
    .i_aic_4_init_lt_axi_s_arsize(i_aic_4_init_lt_axi_s_arsize),
    .i_aic_4_init_lt_axi_s_arvalid(i_aic_4_init_lt_axi_s_arvalid),
    .i_aic_4_init_lt_axi_s_awaddr(i_aic_4_init_lt_axi_s_awaddr),
    .i_aic_4_init_lt_axi_s_awburst(i_aic_4_init_lt_axi_s_awburst),
    .i_aic_4_init_lt_axi_s_awcache(i_aic_4_init_lt_axi_s_awcache),
    .i_aic_4_init_lt_axi_s_awid(i_aic_4_init_lt_axi_s_awid),
    .i_aic_4_init_lt_axi_s_awlen(i_aic_4_init_lt_axi_s_awlen),
    .i_aic_4_init_lt_axi_s_awlock(i_aic_4_init_lt_axi_s_awlock),
    .i_aic_4_init_lt_axi_s_awprot(i_aic_4_init_lt_axi_s_awprot),
    .i_aic_4_init_lt_axi_s_awqos(i_aic_4_init_lt_axi_s_awqos),
    .o_aic_4_init_lt_axi_s_awready(o_aic_4_init_lt_axi_s_awready),
    .i_aic_4_init_lt_axi_s_awsize(i_aic_4_init_lt_axi_s_awsize),
    .i_aic_4_init_lt_axi_s_awvalid(i_aic_4_init_lt_axi_s_awvalid),
    .o_aic_4_init_lt_axi_s_bid(o_aic_4_init_lt_axi_s_bid),
    .i_aic_4_init_lt_axi_s_bready(i_aic_4_init_lt_axi_s_bready),
    .o_aic_4_init_lt_axi_s_bresp(o_aic_4_init_lt_axi_s_bresp),
    .o_aic_4_init_lt_axi_s_bvalid(o_aic_4_init_lt_axi_s_bvalid),
    .o_aic_4_init_lt_axi_s_rdata(o_aic_4_init_lt_axi_s_rdata),
    .o_aic_4_init_lt_axi_s_rid(o_aic_4_init_lt_axi_s_rid),
    .o_aic_4_init_lt_axi_s_rlast(o_aic_4_init_lt_axi_s_rlast),
    .i_aic_4_init_lt_axi_s_rready(i_aic_4_init_lt_axi_s_rready),
    .o_aic_4_init_lt_axi_s_rresp(o_aic_4_init_lt_axi_s_rresp),
    .o_aic_4_init_lt_axi_s_rvalid(o_aic_4_init_lt_axi_s_rvalid),
    .i_aic_4_init_lt_axi_s_wdata(i_aic_4_init_lt_axi_s_wdata),
    .i_aic_4_init_lt_axi_s_wlast(i_aic_4_init_lt_axi_s_wlast),
    .o_aic_4_init_lt_axi_s_wready(o_aic_4_init_lt_axi_s_wready),
    .i_aic_4_init_lt_axi_s_wstrb(i_aic_4_init_lt_axi_s_wstrb),
    .i_aic_4_init_lt_axi_s_wvalid(i_aic_4_init_lt_axi_s_wvalid),
    .o_aic_4_pwr_idle_val(o_aic_4_pwr_idle_val),
    .o_aic_4_pwr_idle_ack(o_aic_4_pwr_idle_ack),
    .i_aic_4_pwr_idle_req(i_aic_4_pwr_idle_req),
    .i_aic_4_rst_n(i_aic_4_rst_n),
    .o_aic_4_targ_lt_axi_m_araddr(o_aic_4_targ_lt_axi_m_araddr),
    .o_aic_4_targ_lt_axi_m_arburst(o_aic_4_targ_lt_axi_m_arburst),
    .o_aic_4_targ_lt_axi_m_arcache(o_aic_4_targ_lt_axi_m_arcache),
    .o_aic_4_targ_lt_axi_m_arid(o_aic_4_targ_lt_axi_m_arid),
    .o_aic_4_targ_lt_axi_m_arlen(o_aic_4_targ_lt_axi_m_arlen),
    .o_aic_4_targ_lt_axi_m_arlock(o_aic_4_targ_lt_axi_m_arlock),
    .o_aic_4_targ_lt_axi_m_arprot(o_aic_4_targ_lt_axi_m_arprot),
    .o_aic_4_targ_lt_axi_m_arqos(o_aic_4_targ_lt_axi_m_arqos),
    .i_aic_4_targ_lt_axi_m_arready(i_aic_4_targ_lt_axi_m_arready),
    .o_aic_4_targ_lt_axi_m_arsize(o_aic_4_targ_lt_axi_m_arsize),
    .o_aic_4_targ_lt_axi_m_arvalid(o_aic_4_targ_lt_axi_m_arvalid),
    .o_aic_4_targ_lt_axi_m_awaddr(o_aic_4_targ_lt_axi_m_awaddr),
    .o_aic_4_targ_lt_axi_m_awburst(o_aic_4_targ_lt_axi_m_awburst),
    .o_aic_4_targ_lt_axi_m_awcache(o_aic_4_targ_lt_axi_m_awcache),
    .o_aic_4_targ_lt_axi_m_awid(o_aic_4_targ_lt_axi_m_awid),
    .o_aic_4_targ_lt_axi_m_awlen(o_aic_4_targ_lt_axi_m_awlen),
    .o_aic_4_targ_lt_axi_m_awlock(o_aic_4_targ_lt_axi_m_awlock),
    .o_aic_4_targ_lt_axi_m_awprot(o_aic_4_targ_lt_axi_m_awprot),
    .o_aic_4_targ_lt_axi_m_awqos(o_aic_4_targ_lt_axi_m_awqos),
    .i_aic_4_targ_lt_axi_m_awready(i_aic_4_targ_lt_axi_m_awready),
    .o_aic_4_targ_lt_axi_m_awsize(o_aic_4_targ_lt_axi_m_awsize),
    .o_aic_4_targ_lt_axi_m_awvalid(o_aic_4_targ_lt_axi_m_awvalid),
    .i_aic_4_targ_lt_axi_m_bid(i_aic_4_targ_lt_axi_m_bid),
    .o_aic_4_targ_lt_axi_m_bready(o_aic_4_targ_lt_axi_m_bready),
    .i_aic_4_targ_lt_axi_m_bresp(i_aic_4_targ_lt_axi_m_bresp),
    .i_aic_4_targ_lt_axi_m_bvalid(i_aic_4_targ_lt_axi_m_bvalid),
    .i_aic_4_targ_lt_axi_m_rdata(i_aic_4_targ_lt_axi_m_rdata),
    .i_aic_4_targ_lt_axi_m_rid(i_aic_4_targ_lt_axi_m_rid),
    .i_aic_4_targ_lt_axi_m_rlast(i_aic_4_targ_lt_axi_m_rlast),
    .o_aic_4_targ_lt_axi_m_rready(o_aic_4_targ_lt_axi_m_rready),
    .i_aic_4_targ_lt_axi_m_rresp(i_aic_4_targ_lt_axi_m_rresp),
    .i_aic_4_targ_lt_axi_m_rvalid(i_aic_4_targ_lt_axi_m_rvalid),
    .o_aic_4_targ_lt_axi_m_wdata(o_aic_4_targ_lt_axi_m_wdata),
    .o_aic_4_targ_lt_axi_m_wlast(o_aic_4_targ_lt_axi_m_wlast),
    .i_aic_4_targ_lt_axi_m_wready(i_aic_4_targ_lt_axi_m_wready),
    .o_aic_4_targ_lt_axi_m_wstrb(o_aic_4_targ_lt_axi_m_wstrb),
    .o_aic_4_targ_lt_axi_m_wvalid(o_aic_4_targ_lt_axi_m_wvalid),
    .o_aic_4_targ_syscfg_apb_m_paddr(o_aic_4_targ_syscfg_apb_m_paddr),
    .o_aic_4_targ_syscfg_apb_m_penable(o_aic_4_targ_syscfg_apb_m_penable),
    .o_aic_4_targ_syscfg_apb_m_pprot(o_aic_4_targ_syscfg_apb_m_pprot),
    .i_aic_4_targ_syscfg_apb_m_prdata(i_aic_4_targ_syscfg_apb_m_prdata),
    .i_aic_4_targ_syscfg_apb_m_pready(i_aic_4_targ_syscfg_apb_m_pready),
    .o_aic_4_targ_syscfg_apb_m_psel(o_aic_4_targ_syscfg_apb_m_psel),
    .i_aic_4_targ_syscfg_apb_m_pslverr(i_aic_4_targ_syscfg_apb_m_pslverr),
    .o_aic_4_targ_syscfg_apb_m_pstrb(o_aic_4_targ_syscfg_apb_m_pstrb),
    .o_aic_4_targ_syscfg_apb_m_pwdata(o_aic_4_targ_syscfg_apb_m_pwdata),
    .o_aic_4_targ_syscfg_apb_m_pwrite(o_aic_4_targ_syscfg_apb_m_pwrite),
    .i_aic_5_aon_clk(i_aic_5_aon_clk),
    .i_aic_5_aon_rst_n(aic_5_aon_rst_n_synced),
    .i_aic_5_clk(i_aic_5_clk),
    .i_aic_5_clken(i_aic_5_clken),
    .i_aic_5_init_ht_axi_s_araddr(i_aic_5_init_ht_axi_s_araddr),
    .i_aic_5_init_ht_axi_s_arburst(i_aic_5_init_ht_axi_s_arburst),
    .i_aic_5_init_ht_axi_s_arcache(i_aic_5_init_ht_axi_s_arcache),
    .i_aic_5_init_ht_axi_s_arid(i_aic_5_init_ht_axi_s_arid),
    .i_aic_5_init_ht_axi_s_arlen(i_aic_5_init_ht_axi_s_arlen),
    .i_aic_5_init_ht_axi_s_arlock(i_aic_5_init_ht_axi_s_arlock),
    .i_aic_5_init_ht_axi_s_arprot(i_aic_5_init_ht_axi_s_arprot),
    .o_aic_5_init_ht_axi_s_arready(o_aic_5_init_ht_axi_s_arready),
    .i_aic_5_init_ht_axi_s_arsize(i_aic_5_init_ht_axi_s_arsize),
    .i_aic_5_init_ht_axi_s_arvalid(i_aic_5_init_ht_axi_s_arvalid),
    .o_aic_5_init_ht_axi_s_rdata(o_aic_5_init_ht_axi_s_rdata),
    .o_aic_5_init_ht_axi_s_rid(o_aic_5_init_ht_axi_s_rid),
    .o_aic_5_init_ht_axi_s_rlast(o_aic_5_init_ht_axi_s_rlast),
    .i_aic_5_init_ht_axi_s_rready(i_aic_5_init_ht_axi_s_rready),
    .o_aic_5_init_ht_axi_s_rresp(o_aic_5_init_ht_axi_s_rresp),
    .o_aic_5_init_ht_axi_s_rvalid(o_aic_5_init_ht_axi_s_rvalid),
    .i_aic_5_init_ht_axi_s_awaddr(i_aic_5_init_ht_axi_s_awaddr),
    .i_aic_5_init_ht_axi_s_awburst(i_aic_5_init_ht_axi_s_awburst),
    .i_aic_5_init_ht_axi_s_awcache(i_aic_5_init_ht_axi_s_awcache),
    .i_aic_5_init_ht_axi_s_awid(i_aic_5_init_ht_axi_s_awid),
    .i_aic_5_init_ht_axi_s_awlen(i_aic_5_init_ht_axi_s_awlen),
    .i_aic_5_init_ht_axi_s_awlock(i_aic_5_init_ht_axi_s_awlock),
    .i_aic_5_init_ht_axi_s_awprot(i_aic_5_init_ht_axi_s_awprot),
    .o_aic_5_init_ht_axi_s_awready(o_aic_5_init_ht_axi_s_awready),
    .i_aic_5_init_ht_axi_s_awsize(i_aic_5_init_ht_axi_s_awsize),
    .i_aic_5_init_ht_axi_s_awvalid(i_aic_5_init_ht_axi_s_awvalid),
    .o_aic_5_init_ht_axi_s_bid(o_aic_5_init_ht_axi_s_bid),
    .i_aic_5_init_ht_axi_s_bready(i_aic_5_init_ht_axi_s_bready),
    .o_aic_5_init_ht_axi_s_bresp(o_aic_5_init_ht_axi_s_bresp),
    .o_aic_5_init_ht_axi_s_bvalid(o_aic_5_init_ht_axi_s_bvalid),
    .i_aic_5_init_ht_axi_s_wdata(i_aic_5_init_ht_axi_s_wdata),
    .i_aic_5_init_ht_axi_s_wlast(i_aic_5_init_ht_axi_s_wlast),
    .o_aic_5_init_ht_axi_s_wready(o_aic_5_init_ht_axi_s_wready),
    .i_aic_5_init_ht_axi_s_wstrb(i_aic_5_init_ht_axi_s_wstrb),
    .i_aic_5_init_ht_axi_s_wvalid(i_aic_5_init_ht_axi_s_wvalid),
    .i_aic_5_init_lt_axi_s_araddr(i_aic_5_init_lt_axi_s_araddr),
    .i_aic_5_init_lt_axi_s_arburst(i_aic_5_init_lt_axi_s_arburst),
    .i_aic_5_init_lt_axi_s_arcache(i_aic_5_init_lt_axi_s_arcache),
    .i_aic_5_init_lt_axi_s_arid(i_aic_5_init_lt_axi_s_arid),
    .i_aic_5_init_lt_axi_s_arlen(i_aic_5_init_lt_axi_s_arlen),
    .i_aic_5_init_lt_axi_s_arlock(i_aic_5_init_lt_axi_s_arlock),
    .i_aic_5_init_lt_axi_s_arprot(i_aic_5_init_lt_axi_s_arprot),
    .i_aic_5_init_lt_axi_s_arqos(i_aic_5_init_lt_axi_s_arqos),
    .o_aic_5_init_lt_axi_s_arready(o_aic_5_init_lt_axi_s_arready),
    .i_aic_5_init_lt_axi_s_arsize(i_aic_5_init_lt_axi_s_arsize),
    .i_aic_5_init_lt_axi_s_arvalid(i_aic_5_init_lt_axi_s_arvalid),
    .i_aic_5_init_lt_axi_s_awaddr(i_aic_5_init_lt_axi_s_awaddr),
    .i_aic_5_init_lt_axi_s_awburst(i_aic_5_init_lt_axi_s_awburst),
    .i_aic_5_init_lt_axi_s_awcache(i_aic_5_init_lt_axi_s_awcache),
    .i_aic_5_init_lt_axi_s_awid(i_aic_5_init_lt_axi_s_awid),
    .i_aic_5_init_lt_axi_s_awlen(i_aic_5_init_lt_axi_s_awlen),
    .i_aic_5_init_lt_axi_s_awlock(i_aic_5_init_lt_axi_s_awlock),
    .i_aic_5_init_lt_axi_s_awprot(i_aic_5_init_lt_axi_s_awprot),
    .i_aic_5_init_lt_axi_s_awqos(i_aic_5_init_lt_axi_s_awqos),
    .o_aic_5_init_lt_axi_s_awready(o_aic_5_init_lt_axi_s_awready),
    .i_aic_5_init_lt_axi_s_awsize(i_aic_5_init_lt_axi_s_awsize),
    .i_aic_5_init_lt_axi_s_awvalid(i_aic_5_init_lt_axi_s_awvalid),
    .o_aic_5_init_lt_axi_s_bid(o_aic_5_init_lt_axi_s_bid),
    .i_aic_5_init_lt_axi_s_bready(i_aic_5_init_lt_axi_s_bready),
    .o_aic_5_init_lt_axi_s_bresp(o_aic_5_init_lt_axi_s_bresp),
    .o_aic_5_init_lt_axi_s_bvalid(o_aic_5_init_lt_axi_s_bvalid),
    .o_aic_5_init_lt_axi_s_rdata(o_aic_5_init_lt_axi_s_rdata),
    .o_aic_5_init_lt_axi_s_rid(o_aic_5_init_lt_axi_s_rid),
    .o_aic_5_init_lt_axi_s_rlast(o_aic_5_init_lt_axi_s_rlast),
    .i_aic_5_init_lt_axi_s_rready(i_aic_5_init_lt_axi_s_rready),
    .o_aic_5_init_lt_axi_s_rresp(o_aic_5_init_lt_axi_s_rresp),
    .o_aic_5_init_lt_axi_s_rvalid(o_aic_5_init_lt_axi_s_rvalid),
    .i_aic_5_init_lt_axi_s_wdata(i_aic_5_init_lt_axi_s_wdata),
    .i_aic_5_init_lt_axi_s_wlast(i_aic_5_init_lt_axi_s_wlast),
    .o_aic_5_init_lt_axi_s_wready(o_aic_5_init_lt_axi_s_wready),
    .i_aic_5_init_lt_axi_s_wstrb(i_aic_5_init_lt_axi_s_wstrb),
    .i_aic_5_init_lt_axi_s_wvalid(i_aic_5_init_lt_axi_s_wvalid),
    .o_aic_5_pwr_idle_val(o_aic_5_pwr_idle_val),
    .o_aic_5_pwr_idle_ack(o_aic_5_pwr_idle_ack),
    .i_aic_5_pwr_idle_req(i_aic_5_pwr_idle_req),
    .i_aic_5_rst_n(i_aic_5_rst_n),
    .o_aic_5_targ_lt_axi_m_araddr(o_aic_5_targ_lt_axi_m_araddr),
    .o_aic_5_targ_lt_axi_m_arburst(o_aic_5_targ_lt_axi_m_arburst),
    .o_aic_5_targ_lt_axi_m_arcache(o_aic_5_targ_lt_axi_m_arcache),
    .o_aic_5_targ_lt_axi_m_arid(o_aic_5_targ_lt_axi_m_arid),
    .o_aic_5_targ_lt_axi_m_arlen(o_aic_5_targ_lt_axi_m_arlen),
    .o_aic_5_targ_lt_axi_m_arlock(o_aic_5_targ_lt_axi_m_arlock),
    .o_aic_5_targ_lt_axi_m_arprot(o_aic_5_targ_lt_axi_m_arprot),
    .o_aic_5_targ_lt_axi_m_arqos(o_aic_5_targ_lt_axi_m_arqos),
    .i_aic_5_targ_lt_axi_m_arready(i_aic_5_targ_lt_axi_m_arready),
    .o_aic_5_targ_lt_axi_m_arsize(o_aic_5_targ_lt_axi_m_arsize),
    .o_aic_5_targ_lt_axi_m_arvalid(o_aic_5_targ_lt_axi_m_arvalid),
    .o_aic_5_targ_lt_axi_m_awaddr(o_aic_5_targ_lt_axi_m_awaddr),
    .o_aic_5_targ_lt_axi_m_awburst(o_aic_5_targ_lt_axi_m_awburst),
    .o_aic_5_targ_lt_axi_m_awcache(o_aic_5_targ_lt_axi_m_awcache),
    .o_aic_5_targ_lt_axi_m_awid(o_aic_5_targ_lt_axi_m_awid),
    .o_aic_5_targ_lt_axi_m_awlen(o_aic_5_targ_lt_axi_m_awlen),
    .o_aic_5_targ_lt_axi_m_awlock(o_aic_5_targ_lt_axi_m_awlock),
    .o_aic_5_targ_lt_axi_m_awprot(o_aic_5_targ_lt_axi_m_awprot),
    .o_aic_5_targ_lt_axi_m_awqos(o_aic_5_targ_lt_axi_m_awqos),
    .i_aic_5_targ_lt_axi_m_awready(i_aic_5_targ_lt_axi_m_awready),
    .o_aic_5_targ_lt_axi_m_awsize(o_aic_5_targ_lt_axi_m_awsize),
    .o_aic_5_targ_lt_axi_m_awvalid(o_aic_5_targ_lt_axi_m_awvalid),
    .i_aic_5_targ_lt_axi_m_bid(i_aic_5_targ_lt_axi_m_bid),
    .o_aic_5_targ_lt_axi_m_bready(o_aic_5_targ_lt_axi_m_bready),
    .i_aic_5_targ_lt_axi_m_bresp(i_aic_5_targ_lt_axi_m_bresp),
    .i_aic_5_targ_lt_axi_m_bvalid(i_aic_5_targ_lt_axi_m_bvalid),
    .i_aic_5_targ_lt_axi_m_rdata(i_aic_5_targ_lt_axi_m_rdata),
    .i_aic_5_targ_lt_axi_m_rid(i_aic_5_targ_lt_axi_m_rid),
    .i_aic_5_targ_lt_axi_m_rlast(i_aic_5_targ_lt_axi_m_rlast),
    .o_aic_5_targ_lt_axi_m_rready(o_aic_5_targ_lt_axi_m_rready),
    .i_aic_5_targ_lt_axi_m_rresp(i_aic_5_targ_lt_axi_m_rresp),
    .i_aic_5_targ_lt_axi_m_rvalid(i_aic_5_targ_lt_axi_m_rvalid),
    .o_aic_5_targ_lt_axi_m_wdata(o_aic_5_targ_lt_axi_m_wdata),
    .o_aic_5_targ_lt_axi_m_wlast(o_aic_5_targ_lt_axi_m_wlast),
    .i_aic_5_targ_lt_axi_m_wready(i_aic_5_targ_lt_axi_m_wready),
    .o_aic_5_targ_lt_axi_m_wstrb(o_aic_5_targ_lt_axi_m_wstrb),
    .o_aic_5_targ_lt_axi_m_wvalid(o_aic_5_targ_lt_axi_m_wvalid),
    .o_aic_5_targ_syscfg_apb_m_paddr(o_aic_5_targ_syscfg_apb_m_paddr),
    .o_aic_5_targ_syscfg_apb_m_penable(o_aic_5_targ_syscfg_apb_m_penable),
    .o_aic_5_targ_syscfg_apb_m_pprot(o_aic_5_targ_syscfg_apb_m_pprot),
    .i_aic_5_targ_syscfg_apb_m_prdata(i_aic_5_targ_syscfg_apb_m_prdata),
    .i_aic_5_targ_syscfg_apb_m_pready(i_aic_5_targ_syscfg_apb_m_pready),
    .o_aic_5_targ_syscfg_apb_m_psel(o_aic_5_targ_syscfg_apb_m_psel),
    .i_aic_5_targ_syscfg_apb_m_pslverr(i_aic_5_targ_syscfg_apb_m_pslverr),
    .o_aic_5_targ_syscfg_apb_m_pstrb(o_aic_5_targ_syscfg_apb_m_pstrb),
    .o_aic_5_targ_syscfg_apb_m_pwdata(o_aic_5_targ_syscfg_apb_m_pwdata),
    .o_aic_5_targ_syscfg_apb_m_pwrite(o_aic_5_targ_syscfg_apb_m_pwrite),
    .i_aic_6_aon_clk(i_aic_6_aon_clk),
    .i_aic_6_aon_rst_n(aic_6_aon_rst_n_synced),
    .i_aic_6_clk(i_aic_6_clk),
    .i_aic_6_clken(i_aic_6_clken),
    .i_aic_6_init_ht_axi_s_araddr(i_aic_6_init_ht_axi_s_araddr),
    .i_aic_6_init_ht_axi_s_arburst(i_aic_6_init_ht_axi_s_arburst),
    .i_aic_6_init_ht_axi_s_arcache(i_aic_6_init_ht_axi_s_arcache),
    .i_aic_6_init_ht_axi_s_arid(i_aic_6_init_ht_axi_s_arid),
    .i_aic_6_init_ht_axi_s_arlen(i_aic_6_init_ht_axi_s_arlen),
    .i_aic_6_init_ht_axi_s_arlock(i_aic_6_init_ht_axi_s_arlock),
    .i_aic_6_init_ht_axi_s_arprot(i_aic_6_init_ht_axi_s_arprot),
    .o_aic_6_init_ht_axi_s_arready(o_aic_6_init_ht_axi_s_arready),
    .i_aic_6_init_ht_axi_s_arsize(i_aic_6_init_ht_axi_s_arsize),
    .i_aic_6_init_ht_axi_s_arvalid(i_aic_6_init_ht_axi_s_arvalid),
    .o_aic_6_init_ht_axi_s_rdata(o_aic_6_init_ht_axi_s_rdata),
    .o_aic_6_init_ht_axi_s_rid(o_aic_6_init_ht_axi_s_rid),
    .o_aic_6_init_ht_axi_s_rlast(o_aic_6_init_ht_axi_s_rlast),
    .i_aic_6_init_ht_axi_s_rready(i_aic_6_init_ht_axi_s_rready),
    .o_aic_6_init_ht_axi_s_rresp(o_aic_6_init_ht_axi_s_rresp),
    .o_aic_6_init_ht_axi_s_rvalid(o_aic_6_init_ht_axi_s_rvalid),
    .i_aic_6_init_ht_axi_s_awaddr(i_aic_6_init_ht_axi_s_awaddr),
    .i_aic_6_init_ht_axi_s_awburst(i_aic_6_init_ht_axi_s_awburst),
    .i_aic_6_init_ht_axi_s_awcache(i_aic_6_init_ht_axi_s_awcache),
    .i_aic_6_init_ht_axi_s_awid(i_aic_6_init_ht_axi_s_awid),
    .i_aic_6_init_ht_axi_s_awlen(i_aic_6_init_ht_axi_s_awlen),
    .i_aic_6_init_ht_axi_s_awlock(i_aic_6_init_ht_axi_s_awlock),
    .i_aic_6_init_ht_axi_s_awprot(i_aic_6_init_ht_axi_s_awprot),
    .o_aic_6_init_ht_axi_s_awready(o_aic_6_init_ht_axi_s_awready),
    .i_aic_6_init_ht_axi_s_awsize(i_aic_6_init_ht_axi_s_awsize),
    .i_aic_6_init_ht_axi_s_awvalid(i_aic_6_init_ht_axi_s_awvalid),
    .o_aic_6_init_ht_axi_s_bid(o_aic_6_init_ht_axi_s_bid),
    .i_aic_6_init_ht_axi_s_bready(i_aic_6_init_ht_axi_s_bready),
    .o_aic_6_init_ht_axi_s_bresp(o_aic_6_init_ht_axi_s_bresp),
    .o_aic_6_init_ht_axi_s_bvalid(o_aic_6_init_ht_axi_s_bvalid),
    .i_aic_6_init_ht_axi_s_wdata(i_aic_6_init_ht_axi_s_wdata),
    .i_aic_6_init_ht_axi_s_wlast(i_aic_6_init_ht_axi_s_wlast),
    .o_aic_6_init_ht_axi_s_wready(o_aic_6_init_ht_axi_s_wready),
    .i_aic_6_init_ht_axi_s_wstrb(i_aic_6_init_ht_axi_s_wstrb),
    .i_aic_6_init_ht_axi_s_wvalid(i_aic_6_init_ht_axi_s_wvalid),
    .i_aic_6_init_lt_axi_s_araddr(i_aic_6_init_lt_axi_s_araddr),
    .i_aic_6_init_lt_axi_s_arburst(i_aic_6_init_lt_axi_s_arburst),
    .i_aic_6_init_lt_axi_s_arcache(i_aic_6_init_lt_axi_s_arcache),
    .i_aic_6_init_lt_axi_s_arid(i_aic_6_init_lt_axi_s_arid),
    .i_aic_6_init_lt_axi_s_arlen(i_aic_6_init_lt_axi_s_arlen),
    .i_aic_6_init_lt_axi_s_arlock(i_aic_6_init_lt_axi_s_arlock),
    .i_aic_6_init_lt_axi_s_arprot(i_aic_6_init_lt_axi_s_arprot),
    .i_aic_6_init_lt_axi_s_arqos(i_aic_6_init_lt_axi_s_arqos),
    .o_aic_6_init_lt_axi_s_arready(o_aic_6_init_lt_axi_s_arready),
    .i_aic_6_init_lt_axi_s_arsize(i_aic_6_init_lt_axi_s_arsize),
    .i_aic_6_init_lt_axi_s_arvalid(i_aic_6_init_lt_axi_s_arvalid),
    .i_aic_6_init_lt_axi_s_awaddr(i_aic_6_init_lt_axi_s_awaddr),
    .i_aic_6_init_lt_axi_s_awburst(i_aic_6_init_lt_axi_s_awburst),
    .i_aic_6_init_lt_axi_s_awcache(i_aic_6_init_lt_axi_s_awcache),
    .i_aic_6_init_lt_axi_s_awid(i_aic_6_init_lt_axi_s_awid),
    .i_aic_6_init_lt_axi_s_awlen(i_aic_6_init_lt_axi_s_awlen),
    .i_aic_6_init_lt_axi_s_awlock(i_aic_6_init_lt_axi_s_awlock),
    .i_aic_6_init_lt_axi_s_awprot(i_aic_6_init_lt_axi_s_awprot),
    .i_aic_6_init_lt_axi_s_awqos(i_aic_6_init_lt_axi_s_awqos),
    .o_aic_6_init_lt_axi_s_awready(o_aic_6_init_lt_axi_s_awready),
    .i_aic_6_init_lt_axi_s_awsize(i_aic_6_init_lt_axi_s_awsize),
    .i_aic_6_init_lt_axi_s_awvalid(i_aic_6_init_lt_axi_s_awvalid),
    .o_aic_6_init_lt_axi_s_bid(o_aic_6_init_lt_axi_s_bid),
    .i_aic_6_init_lt_axi_s_bready(i_aic_6_init_lt_axi_s_bready),
    .o_aic_6_init_lt_axi_s_bresp(o_aic_6_init_lt_axi_s_bresp),
    .o_aic_6_init_lt_axi_s_bvalid(o_aic_6_init_lt_axi_s_bvalid),
    .o_aic_6_init_lt_axi_s_rdata(o_aic_6_init_lt_axi_s_rdata),
    .o_aic_6_init_lt_axi_s_rid(o_aic_6_init_lt_axi_s_rid),
    .o_aic_6_init_lt_axi_s_rlast(o_aic_6_init_lt_axi_s_rlast),
    .i_aic_6_init_lt_axi_s_rready(i_aic_6_init_lt_axi_s_rready),
    .o_aic_6_init_lt_axi_s_rresp(o_aic_6_init_lt_axi_s_rresp),
    .o_aic_6_init_lt_axi_s_rvalid(o_aic_6_init_lt_axi_s_rvalid),
    .i_aic_6_init_lt_axi_s_wdata(i_aic_6_init_lt_axi_s_wdata),
    .i_aic_6_init_lt_axi_s_wlast(i_aic_6_init_lt_axi_s_wlast),
    .o_aic_6_init_lt_axi_s_wready(o_aic_6_init_lt_axi_s_wready),
    .i_aic_6_init_lt_axi_s_wstrb(i_aic_6_init_lt_axi_s_wstrb),
    .i_aic_6_init_lt_axi_s_wvalid(i_aic_6_init_lt_axi_s_wvalid),
    .o_aic_6_pwr_idle_val(o_aic_6_pwr_idle_val),
    .o_aic_6_pwr_idle_ack(o_aic_6_pwr_idle_ack),
    .i_aic_6_pwr_idle_req(i_aic_6_pwr_idle_req),
    .i_aic_6_rst_n(i_aic_6_rst_n),
    .o_aic_6_targ_lt_axi_m_araddr(o_aic_6_targ_lt_axi_m_araddr),
    .o_aic_6_targ_lt_axi_m_arburst(o_aic_6_targ_lt_axi_m_arburst),
    .o_aic_6_targ_lt_axi_m_arcache(o_aic_6_targ_lt_axi_m_arcache),
    .o_aic_6_targ_lt_axi_m_arid(o_aic_6_targ_lt_axi_m_arid),
    .o_aic_6_targ_lt_axi_m_arlen(o_aic_6_targ_lt_axi_m_arlen),
    .o_aic_6_targ_lt_axi_m_arlock(o_aic_6_targ_lt_axi_m_arlock),
    .o_aic_6_targ_lt_axi_m_arprot(o_aic_6_targ_lt_axi_m_arprot),
    .o_aic_6_targ_lt_axi_m_arqos(o_aic_6_targ_lt_axi_m_arqos),
    .i_aic_6_targ_lt_axi_m_arready(i_aic_6_targ_lt_axi_m_arready),
    .o_aic_6_targ_lt_axi_m_arsize(o_aic_6_targ_lt_axi_m_arsize),
    .o_aic_6_targ_lt_axi_m_arvalid(o_aic_6_targ_lt_axi_m_arvalid),
    .o_aic_6_targ_lt_axi_m_awaddr(o_aic_6_targ_lt_axi_m_awaddr),
    .o_aic_6_targ_lt_axi_m_awburst(o_aic_6_targ_lt_axi_m_awburst),
    .o_aic_6_targ_lt_axi_m_awcache(o_aic_6_targ_lt_axi_m_awcache),
    .o_aic_6_targ_lt_axi_m_awid(o_aic_6_targ_lt_axi_m_awid),
    .o_aic_6_targ_lt_axi_m_awlen(o_aic_6_targ_lt_axi_m_awlen),
    .o_aic_6_targ_lt_axi_m_awlock(o_aic_6_targ_lt_axi_m_awlock),
    .o_aic_6_targ_lt_axi_m_awprot(o_aic_6_targ_lt_axi_m_awprot),
    .o_aic_6_targ_lt_axi_m_awqos(o_aic_6_targ_lt_axi_m_awqos),
    .i_aic_6_targ_lt_axi_m_awready(i_aic_6_targ_lt_axi_m_awready),
    .o_aic_6_targ_lt_axi_m_awsize(o_aic_6_targ_lt_axi_m_awsize),
    .o_aic_6_targ_lt_axi_m_awvalid(o_aic_6_targ_lt_axi_m_awvalid),
    .i_aic_6_targ_lt_axi_m_bid(i_aic_6_targ_lt_axi_m_bid),
    .o_aic_6_targ_lt_axi_m_bready(o_aic_6_targ_lt_axi_m_bready),
    .i_aic_6_targ_lt_axi_m_bresp(i_aic_6_targ_lt_axi_m_bresp),
    .i_aic_6_targ_lt_axi_m_bvalid(i_aic_6_targ_lt_axi_m_bvalid),
    .i_aic_6_targ_lt_axi_m_rdata(i_aic_6_targ_lt_axi_m_rdata),
    .i_aic_6_targ_lt_axi_m_rid(i_aic_6_targ_lt_axi_m_rid),
    .i_aic_6_targ_lt_axi_m_rlast(i_aic_6_targ_lt_axi_m_rlast),
    .o_aic_6_targ_lt_axi_m_rready(o_aic_6_targ_lt_axi_m_rready),
    .i_aic_6_targ_lt_axi_m_rresp(i_aic_6_targ_lt_axi_m_rresp),
    .i_aic_6_targ_lt_axi_m_rvalid(i_aic_6_targ_lt_axi_m_rvalid),
    .o_aic_6_targ_lt_axi_m_wdata(o_aic_6_targ_lt_axi_m_wdata),
    .o_aic_6_targ_lt_axi_m_wlast(o_aic_6_targ_lt_axi_m_wlast),
    .i_aic_6_targ_lt_axi_m_wready(i_aic_6_targ_lt_axi_m_wready),
    .o_aic_6_targ_lt_axi_m_wstrb(o_aic_6_targ_lt_axi_m_wstrb),
    .o_aic_6_targ_lt_axi_m_wvalid(o_aic_6_targ_lt_axi_m_wvalid),
    .o_aic_6_targ_syscfg_apb_m_paddr(o_aic_6_targ_syscfg_apb_m_paddr),
    .o_aic_6_targ_syscfg_apb_m_penable(o_aic_6_targ_syscfg_apb_m_penable),
    .o_aic_6_targ_syscfg_apb_m_pprot(o_aic_6_targ_syscfg_apb_m_pprot),
    .i_aic_6_targ_syscfg_apb_m_prdata(i_aic_6_targ_syscfg_apb_m_prdata),
    .i_aic_6_targ_syscfg_apb_m_pready(i_aic_6_targ_syscfg_apb_m_pready),
    .o_aic_6_targ_syscfg_apb_m_psel(o_aic_6_targ_syscfg_apb_m_psel),
    .i_aic_6_targ_syscfg_apb_m_pslverr(i_aic_6_targ_syscfg_apb_m_pslverr),
    .o_aic_6_targ_syscfg_apb_m_pstrb(o_aic_6_targ_syscfg_apb_m_pstrb),
    .o_aic_6_targ_syscfg_apb_m_pwdata(o_aic_6_targ_syscfg_apb_m_pwdata),
    .o_aic_6_targ_syscfg_apb_m_pwrite(o_aic_6_targ_syscfg_apb_m_pwrite),
    .i_aic_7_aon_clk(i_aic_7_aon_clk),
    .i_aic_7_aon_rst_n(aic_7_aon_rst_n_synced),
    .i_aic_7_clk(i_aic_7_clk),
    .i_aic_7_clken(i_aic_7_clken),
    .i_aic_7_init_ht_axi_s_araddr(i_aic_7_init_ht_axi_s_araddr),
    .i_aic_7_init_ht_axi_s_arburst(i_aic_7_init_ht_axi_s_arburst),
    .i_aic_7_init_ht_axi_s_arcache(i_aic_7_init_ht_axi_s_arcache),
    .i_aic_7_init_ht_axi_s_arid(i_aic_7_init_ht_axi_s_arid),
    .i_aic_7_init_ht_axi_s_arlen(i_aic_7_init_ht_axi_s_arlen),
    .i_aic_7_init_ht_axi_s_arlock(i_aic_7_init_ht_axi_s_arlock),
    .i_aic_7_init_ht_axi_s_arprot(i_aic_7_init_ht_axi_s_arprot),
    .o_aic_7_init_ht_axi_s_arready(o_aic_7_init_ht_axi_s_arready),
    .i_aic_7_init_ht_axi_s_arsize(i_aic_7_init_ht_axi_s_arsize),
    .i_aic_7_init_ht_axi_s_arvalid(i_aic_7_init_ht_axi_s_arvalid),
    .o_aic_7_init_ht_axi_s_rdata(o_aic_7_init_ht_axi_s_rdata),
    .o_aic_7_init_ht_axi_s_rid(o_aic_7_init_ht_axi_s_rid),
    .o_aic_7_init_ht_axi_s_rlast(o_aic_7_init_ht_axi_s_rlast),
    .i_aic_7_init_ht_axi_s_rready(i_aic_7_init_ht_axi_s_rready),
    .o_aic_7_init_ht_axi_s_rresp(o_aic_7_init_ht_axi_s_rresp),
    .o_aic_7_init_ht_axi_s_rvalid(o_aic_7_init_ht_axi_s_rvalid),
    .i_aic_7_init_ht_axi_s_awaddr(i_aic_7_init_ht_axi_s_awaddr),
    .i_aic_7_init_ht_axi_s_awburst(i_aic_7_init_ht_axi_s_awburst),
    .i_aic_7_init_ht_axi_s_awcache(i_aic_7_init_ht_axi_s_awcache),
    .i_aic_7_init_ht_axi_s_awid(i_aic_7_init_ht_axi_s_awid),
    .i_aic_7_init_ht_axi_s_awlen(i_aic_7_init_ht_axi_s_awlen),
    .i_aic_7_init_ht_axi_s_awlock(i_aic_7_init_ht_axi_s_awlock),
    .i_aic_7_init_ht_axi_s_awprot(i_aic_7_init_ht_axi_s_awprot),
    .o_aic_7_init_ht_axi_s_awready(o_aic_7_init_ht_axi_s_awready),
    .i_aic_7_init_ht_axi_s_awsize(i_aic_7_init_ht_axi_s_awsize),
    .i_aic_7_init_ht_axi_s_awvalid(i_aic_7_init_ht_axi_s_awvalid),
    .o_aic_7_init_ht_axi_s_bid(o_aic_7_init_ht_axi_s_bid),
    .i_aic_7_init_ht_axi_s_bready(i_aic_7_init_ht_axi_s_bready),
    .o_aic_7_init_ht_axi_s_bresp(o_aic_7_init_ht_axi_s_bresp),
    .o_aic_7_init_ht_axi_s_bvalid(o_aic_7_init_ht_axi_s_bvalid),
    .i_aic_7_init_ht_axi_s_wdata(i_aic_7_init_ht_axi_s_wdata),
    .i_aic_7_init_ht_axi_s_wlast(i_aic_7_init_ht_axi_s_wlast),
    .o_aic_7_init_ht_axi_s_wready(o_aic_7_init_ht_axi_s_wready),
    .i_aic_7_init_ht_axi_s_wstrb(i_aic_7_init_ht_axi_s_wstrb),
    .i_aic_7_init_ht_axi_s_wvalid(i_aic_7_init_ht_axi_s_wvalid),
    .i_aic_7_init_lt_axi_s_araddr(i_aic_7_init_lt_axi_s_araddr),
    .i_aic_7_init_lt_axi_s_arburst(i_aic_7_init_lt_axi_s_arburst),
    .i_aic_7_init_lt_axi_s_arcache(i_aic_7_init_lt_axi_s_arcache),
    .i_aic_7_init_lt_axi_s_arid(i_aic_7_init_lt_axi_s_arid),
    .i_aic_7_init_lt_axi_s_arlen(i_aic_7_init_lt_axi_s_arlen),
    .i_aic_7_init_lt_axi_s_arlock(i_aic_7_init_lt_axi_s_arlock),
    .i_aic_7_init_lt_axi_s_arprot(i_aic_7_init_lt_axi_s_arprot),
    .i_aic_7_init_lt_axi_s_arqos(i_aic_7_init_lt_axi_s_arqos),
    .o_aic_7_init_lt_axi_s_arready(o_aic_7_init_lt_axi_s_arready),
    .i_aic_7_init_lt_axi_s_arsize(i_aic_7_init_lt_axi_s_arsize),
    .i_aic_7_init_lt_axi_s_arvalid(i_aic_7_init_lt_axi_s_arvalid),
    .i_aic_7_init_lt_axi_s_awaddr(i_aic_7_init_lt_axi_s_awaddr),
    .i_aic_7_init_lt_axi_s_awburst(i_aic_7_init_lt_axi_s_awburst),
    .i_aic_7_init_lt_axi_s_awcache(i_aic_7_init_lt_axi_s_awcache),
    .i_aic_7_init_lt_axi_s_awid(i_aic_7_init_lt_axi_s_awid),
    .i_aic_7_init_lt_axi_s_awlen(i_aic_7_init_lt_axi_s_awlen),
    .i_aic_7_init_lt_axi_s_awlock(i_aic_7_init_lt_axi_s_awlock),
    .i_aic_7_init_lt_axi_s_awprot(i_aic_7_init_lt_axi_s_awprot),
    .i_aic_7_init_lt_axi_s_awqos(i_aic_7_init_lt_axi_s_awqos),
    .o_aic_7_init_lt_axi_s_awready(o_aic_7_init_lt_axi_s_awready),
    .i_aic_7_init_lt_axi_s_awsize(i_aic_7_init_lt_axi_s_awsize),
    .i_aic_7_init_lt_axi_s_awvalid(i_aic_7_init_lt_axi_s_awvalid),
    .o_aic_7_init_lt_axi_s_bid(o_aic_7_init_lt_axi_s_bid),
    .i_aic_7_init_lt_axi_s_bready(i_aic_7_init_lt_axi_s_bready),
    .o_aic_7_init_lt_axi_s_bresp(o_aic_7_init_lt_axi_s_bresp),
    .o_aic_7_init_lt_axi_s_bvalid(o_aic_7_init_lt_axi_s_bvalid),
    .o_aic_7_init_lt_axi_s_rdata(o_aic_7_init_lt_axi_s_rdata),
    .o_aic_7_init_lt_axi_s_rid(o_aic_7_init_lt_axi_s_rid),
    .o_aic_7_init_lt_axi_s_rlast(o_aic_7_init_lt_axi_s_rlast),
    .i_aic_7_init_lt_axi_s_rready(i_aic_7_init_lt_axi_s_rready),
    .o_aic_7_init_lt_axi_s_rresp(o_aic_7_init_lt_axi_s_rresp),
    .o_aic_7_init_lt_axi_s_rvalid(o_aic_7_init_lt_axi_s_rvalid),
    .i_aic_7_init_lt_axi_s_wdata(i_aic_7_init_lt_axi_s_wdata),
    .i_aic_7_init_lt_axi_s_wlast(i_aic_7_init_lt_axi_s_wlast),
    .o_aic_7_init_lt_axi_s_wready(o_aic_7_init_lt_axi_s_wready),
    .i_aic_7_init_lt_axi_s_wstrb(i_aic_7_init_lt_axi_s_wstrb),
    .i_aic_7_init_lt_axi_s_wvalid(i_aic_7_init_lt_axi_s_wvalid),
    .o_aic_7_pwr_idle_val(o_aic_7_pwr_idle_val),
    .o_aic_7_pwr_idle_ack(o_aic_7_pwr_idle_ack),
    .i_aic_7_pwr_idle_req(i_aic_7_pwr_idle_req),
    .i_aic_7_rst_n(i_aic_7_rst_n),
    .o_aic_7_targ_lt_axi_m_araddr(o_aic_7_targ_lt_axi_m_araddr),
    .o_aic_7_targ_lt_axi_m_arburst(o_aic_7_targ_lt_axi_m_arburst),
    .o_aic_7_targ_lt_axi_m_arcache(o_aic_7_targ_lt_axi_m_arcache),
    .o_aic_7_targ_lt_axi_m_arid(o_aic_7_targ_lt_axi_m_arid),
    .o_aic_7_targ_lt_axi_m_arlen(o_aic_7_targ_lt_axi_m_arlen),
    .o_aic_7_targ_lt_axi_m_arlock(o_aic_7_targ_lt_axi_m_arlock),
    .o_aic_7_targ_lt_axi_m_arprot(o_aic_7_targ_lt_axi_m_arprot),
    .o_aic_7_targ_lt_axi_m_arqos(o_aic_7_targ_lt_axi_m_arqos),
    .i_aic_7_targ_lt_axi_m_arready(i_aic_7_targ_lt_axi_m_arready),
    .o_aic_7_targ_lt_axi_m_arsize(o_aic_7_targ_lt_axi_m_arsize),
    .o_aic_7_targ_lt_axi_m_arvalid(o_aic_7_targ_lt_axi_m_arvalid),
    .o_aic_7_targ_lt_axi_m_awaddr(o_aic_7_targ_lt_axi_m_awaddr),
    .o_aic_7_targ_lt_axi_m_awburst(o_aic_7_targ_lt_axi_m_awburst),
    .o_aic_7_targ_lt_axi_m_awcache(o_aic_7_targ_lt_axi_m_awcache),
    .o_aic_7_targ_lt_axi_m_awid(o_aic_7_targ_lt_axi_m_awid),
    .o_aic_7_targ_lt_axi_m_awlen(o_aic_7_targ_lt_axi_m_awlen),
    .o_aic_7_targ_lt_axi_m_awlock(o_aic_7_targ_lt_axi_m_awlock),
    .o_aic_7_targ_lt_axi_m_awprot(o_aic_7_targ_lt_axi_m_awprot),
    .o_aic_7_targ_lt_axi_m_awqos(o_aic_7_targ_lt_axi_m_awqos),
    .i_aic_7_targ_lt_axi_m_awready(i_aic_7_targ_lt_axi_m_awready),
    .o_aic_7_targ_lt_axi_m_awsize(o_aic_7_targ_lt_axi_m_awsize),
    .o_aic_7_targ_lt_axi_m_awvalid(o_aic_7_targ_lt_axi_m_awvalid),
    .i_aic_7_targ_lt_axi_m_bid(i_aic_7_targ_lt_axi_m_bid),
    .o_aic_7_targ_lt_axi_m_bready(o_aic_7_targ_lt_axi_m_bready),
    .i_aic_7_targ_lt_axi_m_bresp(i_aic_7_targ_lt_axi_m_bresp),
    .i_aic_7_targ_lt_axi_m_bvalid(i_aic_7_targ_lt_axi_m_bvalid),
    .i_aic_7_targ_lt_axi_m_rdata(i_aic_7_targ_lt_axi_m_rdata),
    .i_aic_7_targ_lt_axi_m_rid(i_aic_7_targ_lt_axi_m_rid),
    .i_aic_7_targ_lt_axi_m_rlast(i_aic_7_targ_lt_axi_m_rlast),
    .o_aic_7_targ_lt_axi_m_rready(o_aic_7_targ_lt_axi_m_rready),
    .i_aic_7_targ_lt_axi_m_rresp(i_aic_7_targ_lt_axi_m_rresp),
    .i_aic_7_targ_lt_axi_m_rvalid(i_aic_7_targ_lt_axi_m_rvalid),
    .o_aic_7_targ_lt_axi_m_wdata(o_aic_7_targ_lt_axi_m_wdata),
    .o_aic_7_targ_lt_axi_m_wlast(o_aic_7_targ_lt_axi_m_wlast),
    .i_aic_7_targ_lt_axi_m_wready(i_aic_7_targ_lt_axi_m_wready),
    .o_aic_7_targ_lt_axi_m_wstrb(o_aic_7_targ_lt_axi_m_wstrb),
    .o_aic_7_targ_lt_axi_m_wvalid(o_aic_7_targ_lt_axi_m_wvalid),
    .o_aic_7_targ_syscfg_apb_m_paddr(o_aic_7_targ_syscfg_apb_m_paddr),
    .o_aic_7_targ_syscfg_apb_m_penable(o_aic_7_targ_syscfg_apb_m_penable),
    .o_aic_7_targ_syscfg_apb_m_pprot(o_aic_7_targ_syscfg_apb_m_pprot),
    .i_aic_7_targ_syscfg_apb_m_prdata(i_aic_7_targ_syscfg_apb_m_prdata),
    .i_aic_7_targ_syscfg_apb_m_pready(i_aic_7_targ_syscfg_apb_m_pready),
    .o_aic_7_targ_syscfg_apb_m_psel(o_aic_7_targ_syscfg_apb_m_psel),
    .i_aic_7_targ_syscfg_apb_m_pslverr(i_aic_7_targ_syscfg_apb_m_pslverr),
    .o_aic_7_targ_syscfg_apb_m_pstrb(o_aic_7_targ_syscfg_apb_m_pstrb),
    .o_aic_7_targ_syscfg_apb_m_pwdata(o_aic_7_targ_syscfg_apb_m_pwdata),
    .o_aic_7_targ_syscfg_apb_m_pwrite(o_aic_7_targ_syscfg_apb_m_pwrite),
    .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data),
    .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head),
    .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy(o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail),
    .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld(i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld),
    .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld(o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data),
    .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head),
    .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy(o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail),
    .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld(i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld),
    .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld(o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data),
    .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head),
    .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy(o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail),
    .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld(i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld),
    .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld(o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data),
    .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head),
    .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy(o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail),
    .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld(i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld),
    .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld(o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data),
    .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head),
    .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy(o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail),
    .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld(i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld),
    .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld(o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data),
    .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head),
    .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy(o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail),
    .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld(i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld),
    .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld(o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data),
    .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head),
    .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy(o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail),
    .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld(i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld),
    .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld(o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data),
    .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head),
    .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy(o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail),
    .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld(i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld),
    .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld(o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data),
    .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head),
    .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy(o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail),
    .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld(i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld),
    .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld(o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data),
    .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head),
    .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy(o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail),
    .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld(i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld),
    .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld(o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data),
    .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head),
    .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy(o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail),
    .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld(i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld),
    .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld(o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data),
    .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head),
    .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy(o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy),
    .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail),
    .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld(i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld),
    .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data),
    .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head),
    .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy(i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld(o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data),
    .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head),
    .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy(o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy),
    .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail),
    .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld(i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld),
    .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data),
    .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head),
    .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy(i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail),
    .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld(o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data),
    .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head),
    .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy(i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail),
    .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld(o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld),
    .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld(i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data),
    .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head),
    .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy(i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail),
    .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld(o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld),
    .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld(i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data),
    .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head),
    .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy(i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail),
    .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld(o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld),
    .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld(i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data),
    .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head),
    .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy(i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail),
    .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld(o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld),
    .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld(i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data),
    .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head),
    .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy(i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail),
    .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld(o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld),
    .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld(i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data),
    .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head),
    .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy(i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail),
    .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld(o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld),
    .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld(i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data),
    .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head),
    .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy(i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail),
    .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld(o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld),
    .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld(i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data),
    .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head),
    .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy(i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail),
    .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld(o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld),
    .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld(i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data),
    .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head),
    .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy(i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail),
    .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld(o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld),
    .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld(i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data),
    .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head),
    .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy(i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail),
    .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld(o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld),
    .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld(i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data),
    .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head),
    .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy(i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail),
    .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld(o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld),
    .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld(i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data),
    .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head),
    .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy(i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy),
    .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail),
    .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld(o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld),
    .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data),
    .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head),
    .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy(o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld(i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data),
    .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head),
    .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy(i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy),
    .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail),
    .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld(o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld),
    .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data),
    .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head),
    .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy(o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy),
    .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail),
    .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld(i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld),
    .i_l2_4_aon_clk(i_l2_4_aon_clk),
    .i_l2_4_aon_rst_n(l2_4_aon_rst_n_synced),
    .i_l2_4_clk(i_l2_4_clk),
    .i_l2_4_clken(i_l2_4_clken),
    .o_l2_4_pwr_idle_val(o_l2_4_pwr_idle_val),
    .o_l2_4_pwr_idle_ack(o_l2_4_pwr_idle_ack),
    .i_l2_4_pwr_idle_req(i_l2_4_pwr_idle_req),
    .i_l2_4_rst_n(i_l2_4_rst_n),
    .o_l2_4_targ_ht_axi_m_araddr(o_l2_4_targ_ht_axi_m_araddr),
    .o_l2_4_targ_ht_axi_m_arburst(o_l2_4_targ_ht_axi_m_arburst),
    .o_l2_4_targ_ht_axi_m_arcache(o_l2_4_targ_ht_axi_m_arcache),
    .o_l2_4_targ_ht_axi_m_arid(o_l2_4_targ_ht_axi_m_arid),
    .o_l2_4_targ_ht_axi_m_arlen(o_l2_4_targ_ht_axi_m_arlen),
    .o_l2_4_targ_ht_axi_m_arlock(o_l2_4_targ_ht_axi_m_arlock),
    .o_l2_4_targ_ht_axi_m_arprot(o_l2_4_targ_ht_axi_m_arprot),
    .i_l2_4_targ_ht_axi_m_arready(i_l2_4_targ_ht_axi_m_arready),
    .o_l2_4_targ_ht_axi_m_arsize(o_l2_4_targ_ht_axi_m_arsize),
    .o_l2_4_targ_ht_axi_m_arvalid(o_l2_4_targ_ht_axi_m_arvalid),
    .i_l2_4_targ_ht_axi_m_rdata(i_l2_4_targ_ht_axi_m_rdata),
    .i_l2_4_targ_ht_axi_m_rid(i_l2_4_targ_ht_axi_m_rid),
    .i_l2_4_targ_ht_axi_m_rlast(i_l2_4_targ_ht_axi_m_rlast),
    .o_l2_4_targ_ht_axi_m_rready(o_l2_4_targ_ht_axi_m_rready),
    .i_l2_4_targ_ht_axi_m_rresp(i_l2_4_targ_ht_axi_m_rresp),
    .i_l2_4_targ_ht_axi_m_rvalid(i_l2_4_targ_ht_axi_m_rvalid),
    .o_l2_4_targ_ht_axi_m_awaddr(o_l2_4_targ_ht_axi_m_awaddr),
    .o_l2_4_targ_ht_axi_m_awburst(o_l2_4_targ_ht_axi_m_awburst),
    .o_l2_4_targ_ht_axi_m_awcache(o_l2_4_targ_ht_axi_m_awcache),
    .o_l2_4_targ_ht_axi_m_awid(o_l2_4_targ_ht_axi_m_awid),
    .o_l2_4_targ_ht_axi_m_awlen(o_l2_4_targ_ht_axi_m_awlen),
    .o_l2_4_targ_ht_axi_m_awlock(o_l2_4_targ_ht_axi_m_awlock),
    .o_l2_4_targ_ht_axi_m_awprot(o_l2_4_targ_ht_axi_m_awprot),
    .i_l2_4_targ_ht_axi_m_awready(i_l2_4_targ_ht_axi_m_awready),
    .o_l2_4_targ_ht_axi_m_awsize(o_l2_4_targ_ht_axi_m_awsize),
    .o_l2_4_targ_ht_axi_m_awvalid(o_l2_4_targ_ht_axi_m_awvalid),
    .i_l2_4_targ_ht_axi_m_bid(i_l2_4_targ_ht_axi_m_bid),
    .o_l2_4_targ_ht_axi_m_bready(o_l2_4_targ_ht_axi_m_bready),
    .i_l2_4_targ_ht_axi_m_bresp(i_l2_4_targ_ht_axi_m_bresp),
    .i_l2_4_targ_ht_axi_m_bvalid(i_l2_4_targ_ht_axi_m_bvalid),
    .o_l2_4_targ_ht_axi_m_wdata(o_l2_4_targ_ht_axi_m_wdata),
    .o_l2_4_targ_ht_axi_m_wlast(o_l2_4_targ_ht_axi_m_wlast),
    .i_l2_4_targ_ht_axi_m_wready(i_l2_4_targ_ht_axi_m_wready),
    .o_l2_4_targ_ht_axi_m_wstrb(o_l2_4_targ_ht_axi_m_wstrb),
    .o_l2_4_targ_ht_axi_m_wvalid(o_l2_4_targ_ht_axi_m_wvalid),
    .o_l2_4_targ_syscfg_apb_m_paddr(o_l2_4_targ_syscfg_apb_m_paddr),
    .o_l2_4_targ_syscfg_apb_m_penable(o_l2_4_targ_syscfg_apb_m_penable),
    .o_l2_4_targ_syscfg_apb_m_pprot(o_l2_4_targ_syscfg_apb_m_pprot),
    .i_l2_4_targ_syscfg_apb_m_prdata(i_l2_4_targ_syscfg_apb_m_prdata),
    .i_l2_4_targ_syscfg_apb_m_pready(i_l2_4_targ_syscfg_apb_m_pready),
    .o_l2_4_targ_syscfg_apb_m_psel(o_l2_4_targ_syscfg_apb_m_psel),
    .i_l2_4_targ_syscfg_apb_m_pslverr(i_l2_4_targ_syscfg_apb_m_pslverr),
    .o_l2_4_targ_syscfg_apb_m_pstrb(o_l2_4_targ_syscfg_apb_m_pstrb),
    .o_l2_4_targ_syscfg_apb_m_pwdata(o_l2_4_targ_syscfg_apb_m_pwdata),
    .o_l2_4_targ_syscfg_apb_m_pwrite(o_l2_4_targ_syscfg_apb_m_pwrite),
    .i_l2_5_aon_clk(i_l2_5_aon_clk),
    .i_l2_5_aon_rst_n(l2_5_aon_rst_n_synced),
    .i_l2_5_clk(i_l2_5_clk),
    .i_l2_5_clken(i_l2_5_clken),
    .o_l2_5_pwr_idle_val(o_l2_5_pwr_idle_val),
    .o_l2_5_pwr_idle_ack(o_l2_5_pwr_idle_ack),
    .i_l2_5_pwr_idle_req(i_l2_5_pwr_idle_req),
    .i_l2_5_rst_n(i_l2_5_rst_n),
    .o_l2_5_targ_ht_axi_m_araddr(o_l2_5_targ_ht_axi_m_araddr),
    .o_l2_5_targ_ht_axi_m_arburst(o_l2_5_targ_ht_axi_m_arburst),
    .o_l2_5_targ_ht_axi_m_arcache(o_l2_5_targ_ht_axi_m_arcache),
    .o_l2_5_targ_ht_axi_m_arid(o_l2_5_targ_ht_axi_m_arid),
    .o_l2_5_targ_ht_axi_m_arlen(o_l2_5_targ_ht_axi_m_arlen),
    .o_l2_5_targ_ht_axi_m_arlock(o_l2_5_targ_ht_axi_m_arlock),
    .o_l2_5_targ_ht_axi_m_arprot(o_l2_5_targ_ht_axi_m_arprot),
    .i_l2_5_targ_ht_axi_m_arready(i_l2_5_targ_ht_axi_m_arready),
    .o_l2_5_targ_ht_axi_m_arsize(o_l2_5_targ_ht_axi_m_arsize),
    .o_l2_5_targ_ht_axi_m_arvalid(o_l2_5_targ_ht_axi_m_arvalid),
    .i_l2_5_targ_ht_axi_m_rdata(i_l2_5_targ_ht_axi_m_rdata),
    .i_l2_5_targ_ht_axi_m_rid(i_l2_5_targ_ht_axi_m_rid),
    .i_l2_5_targ_ht_axi_m_rlast(i_l2_5_targ_ht_axi_m_rlast),
    .o_l2_5_targ_ht_axi_m_rready(o_l2_5_targ_ht_axi_m_rready),
    .i_l2_5_targ_ht_axi_m_rresp(i_l2_5_targ_ht_axi_m_rresp),
    .i_l2_5_targ_ht_axi_m_rvalid(i_l2_5_targ_ht_axi_m_rvalid),
    .o_l2_5_targ_ht_axi_m_awaddr(o_l2_5_targ_ht_axi_m_awaddr),
    .o_l2_5_targ_ht_axi_m_awburst(o_l2_5_targ_ht_axi_m_awburst),
    .o_l2_5_targ_ht_axi_m_awcache(o_l2_5_targ_ht_axi_m_awcache),
    .o_l2_5_targ_ht_axi_m_awid(o_l2_5_targ_ht_axi_m_awid),
    .o_l2_5_targ_ht_axi_m_awlen(o_l2_5_targ_ht_axi_m_awlen),
    .o_l2_5_targ_ht_axi_m_awlock(o_l2_5_targ_ht_axi_m_awlock),
    .o_l2_5_targ_ht_axi_m_awprot(o_l2_5_targ_ht_axi_m_awprot),
    .i_l2_5_targ_ht_axi_m_awready(i_l2_5_targ_ht_axi_m_awready),
    .o_l2_5_targ_ht_axi_m_awsize(o_l2_5_targ_ht_axi_m_awsize),
    .o_l2_5_targ_ht_axi_m_awvalid(o_l2_5_targ_ht_axi_m_awvalid),
    .i_l2_5_targ_ht_axi_m_bid(i_l2_5_targ_ht_axi_m_bid),
    .o_l2_5_targ_ht_axi_m_bready(o_l2_5_targ_ht_axi_m_bready),
    .i_l2_5_targ_ht_axi_m_bresp(i_l2_5_targ_ht_axi_m_bresp),
    .i_l2_5_targ_ht_axi_m_bvalid(i_l2_5_targ_ht_axi_m_bvalid),
    .o_l2_5_targ_ht_axi_m_wdata(o_l2_5_targ_ht_axi_m_wdata),
    .o_l2_5_targ_ht_axi_m_wlast(o_l2_5_targ_ht_axi_m_wlast),
    .i_l2_5_targ_ht_axi_m_wready(i_l2_5_targ_ht_axi_m_wready),
    .o_l2_5_targ_ht_axi_m_wstrb(o_l2_5_targ_ht_axi_m_wstrb),
    .o_l2_5_targ_ht_axi_m_wvalid(o_l2_5_targ_ht_axi_m_wvalid),
    .o_l2_5_targ_syscfg_apb_m_paddr(o_l2_5_targ_syscfg_apb_m_paddr),
    .o_l2_5_targ_syscfg_apb_m_penable(o_l2_5_targ_syscfg_apb_m_penable),
    .o_l2_5_targ_syscfg_apb_m_pprot(o_l2_5_targ_syscfg_apb_m_pprot),
    .i_l2_5_targ_syscfg_apb_m_prdata(i_l2_5_targ_syscfg_apb_m_prdata),
    .i_l2_5_targ_syscfg_apb_m_pready(i_l2_5_targ_syscfg_apb_m_pready),
    .o_l2_5_targ_syscfg_apb_m_psel(o_l2_5_targ_syscfg_apb_m_psel),
    .i_l2_5_targ_syscfg_apb_m_pslverr(i_l2_5_targ_syscfg_apb_m_pslverr),
    .o_l2_5_targ_syscfg_apb_m_pstrb(o_l2_5_targ_syscfg_apb_m_pstrb),
    .o_l2_5_targ_syscfg_apb_m_pwdata(o_l2_5_targ_syscfg_apb_m_pwdata),
    .o_l2_5_targ_syscfg_apb_m_pwrite(o_l2_5_targ_syscfg_apb_m_pwrite),
    .i_l2_6_aon_clk(i_l2_6_aon_clk),
    .i_l2_6_aon_rst_n(l2_6_aon_rst_n_synced),
    .i_l2_6_clk(i_l2_6_clk),
    .i_l2_6_clken(i_l2_6_clken),
    .o_l2_6_pwr_idle_val(o_l2_6_pwr_idle_val),
    .o_l2_6_pwr_idle_ack(o_l2_6_pwr_idle_ack),
    .i_l2_6_pwr_idle_req(i_l2_6_pwr_idle_req),
    .i_l2_6_rst_n(i_l2_6_rst_n),
    .o_l2_6_targ_ht_axi_m_araddr(o_l2_6_targ_ht_axi_m_araddr),
    .o_l2_6_targ_ht_axi_m_arburst(o_l2_6_targ_ht_axi_m_arburst),
    .o_l2_6_targ_ht_axi_m_arcache(o_l2_6_targ_ht_axi_m_arcache),
    .o_l2_6_targ_ht_axi_m_arid(o_l2_6_targ_ht_axi_m_arid),
    .o_l2_6_targ_ht_axi_m_arlen(o_l2_6_targ_ht_axi_m_arlen),
    .o_l2_6_targ_ht_axi_m_arlock(o_l2_6_targ_ht_axi_m_arlock),
    .o_l2_6_targ_ht_axi_m_arprot(o_l2_6_targ_ht_axi_m_arprot),
    .i_l2_6_targ_ht_axi_m_arready(i_l2_6_targ_ht_axi_m_arready),
    .o_l2_6_targ_ht_axi_m_arsize(o_l2_6_targ_ht_axi_m_arsize),
    .o_l2_6_targ_ht_axi_m_arvalid(o_l2_6_targ_ht_axi_m_arvalid),
    .i_l2_6_targ_ht_axi_m_rdata(i_l2_6_targ_ht_axi_m_rdata),
    .i_l2_6_targ_ht_axi_m_rid(i_l2_6_targ_ht_axi_m_rid),
    .i_l2_6_targ_ht_axi_m_rlast(i_l2_6_targ_ht_axi_m_rlast),
    .o_l2_6_targ_ht_axi_m_rready(o_l2_6_targ_ht_axi_m_rready),
    .i_l2_6_targ_ht_axi_m_rresp(i_l2_6_targ_ht_axi_m_rresp),
    .i_l2_6_targ_ht_axi_m_rvalid(i_l2_6_targ_ht_axi_m_rvalid),
    .o_l2_6_targ_ht_axi_m_awaddr(o_l2_6_targ_ht_axi_m_awaddr),
    .o_l2_6_targ_ht_axi_m_awburst(o_l2_6_targ_ht_axi_m_awburst),
    .o_l2_6_targ_ht_axi_m_awcache(o_l2_6_targ_ht_axi_m_awcache),
    .o_l2_6_targ_ht_axi_m_awid(o_l2_6_targ_ht_axi_m_awid),
    .o_l2_6_targ_ht_axi_m_awlen(o_l2_6_targ_ht_axi_m_awlen),
    .o_l2_6_targ_ht_axi_m_awlock(o_l2_6_targ_ht_axi_m_awlock),
    .o_l2_6_targ_ht_axi_m_awprot(o_l2_6_targ_ht_axi_m_awprot),
    .i_l2_6_targ_ht_axi_m_awready(i_l2_6_targ_ht_axi_m_awready),
    .o_l2_6_targ_ht_axi_m_awsize(o_l2_6_targ_ht_axi_m_awsize),
    .o_l2_6_targ_ht_axi_m_awvalid(o_l2_6_targ_ht_axi_m_awvalid),
    .i_l2_6_targ_ht_axi_m_bid(i_l2_6_targ_ht_axi_m_bid),
    .o_l2_6_targ_ht_axi_m_bready(o_l2_6_targ_ht_axi_m_bready),
    .i_l2_6_targ_ht_axi_m_bresp(i_l2_6_targ_ht_axi_m_bresp),
    .i_l2_6_targ_ht_axi_m_bvalid(i_l2_6_targ_ht_axi_m_bvalid),
    .o_l2_6_targ_ht_axi_m_wdata(o_l2_6_targ_ht_axi_m_wdata),
    .o_l2_6_targ_ht_axi_m_wlast(o_l2_6_targ_ht_axi_m_wlast),
    .i_l2_6_targ_ht_axi_m_wready(i_l2_6_targ_ht_axi_m_wready),
    .o_l2_6_targ_ht_axi_m_wstrb(o_l2_6_targ_ht_axi_m_wstrb),
    .o_l2_6_targ_ht_axi_m_wvalid(o_l2_6_targ_ht_axi_m_wvalid),
    .o_l2_6_targ_syscfg_apb_m_paddr(o_l2_6_targ_syscfg_apb_m_paddr),
    .o_l2_6_targ_syscfg_apb_m_penable(o_l2_6_targ_syscfg_apb_m_penable),
    .o_l2_6_targ_syscfg_apb_m_pprot(o_l2_6_targ_syscfg_apb_m_pprot),
    .i_l2_6_targ_syscfg_apb_m_prdata(i_l2_6_targ_syscfg_apb_m_prdata),
    .i_l2_6_targ_syscfg_apb_m_pready(i_l2_6_targ_syscfg_apb_m_pready),
    .o_l2_6_targ_syscfg_apb_m_psel(o_l2_6_targ_syscfg_apb_m_psel),
    .i_l2_6_targ_syscfg_apb_m_pslverr(i_l2_6_targ_syscfg_apb_m_pslverr),
    .o_l2_6_targ_syscfg_apb_m_pstrb(o_l2_6_targ_syscfg_apb_m_pstrb),
    .o_l2_6_targ_syscfg_apb_m_pwdata(o_l2_6_targ_syscfg_apb_m_pwdata),
    .o_l2_6_targ_syscfg_apb_m_pwrite(o_l2_6_targ_syscfg_apb_m_pwrite),
    .i_l2_7_aon_clk(i_l2_7_aon_clk),
    .i_l2_7_aon_rst_n(l2_7_aon_rst_n_synced),
    .i_l2_7_clk(i_l2_7_clk),
    .i_l2_7_clken(i_l2_7_clken),
    .o_l2_7_pwr_idle_val(o_l2_7_pwr_idle_val),
    .o_l2_7_pwr_idle_ack(o_l2_7_pwr_idle_ack),
    .i_l2_7_pwr_idle_req(i_l2_7_pwr_idle_req),
    .i_l2_7_rst_n(i_l2_7_rst_n),
    .o_l2_7_targ_ht_axi_m_araddr(o_l2_7_targ_ht_axi_m_araddr),
    .o_l2_7_targ_ht_axi_m_arburst(o_l2_7_targ_ht_axi_m_arburst),
    .o_l2_7_targ_ht_axi_m_arcache(o_l2_7_targ_ht_axi_m_arcache),
    .o_l2_7_targ_ht_axi_m_arid(o_l2_7_targ_ht_axi_m_arid),
    .o_l2_7_targ_ht_axi_m_arlen(o_l2_7_targ_ht_axi_m_arlen),
    .o_l2_7_targ_ht_axi_m_arlock(o_l2_7_targ_ht_axi_m_arlock),
    .o_l2_7_targ_ht_axi_m_arprot(o_l2_7_targ_ht_axi_m_arprot),
    .i_l2_7_targ_ht_axi_m_arready(i_l2_7_targ_ht_axi_m_arready),
    .o_l2_7_targ_ht_axi_m_arsize(o_l2_7_targ_ht_axi_m_arsize),
    .o_l2_7_targ_ht_axi_m_arvalid(o_l2_7_targ_ht_axi_m_arvalid),
    .i_l2_7_targ_ht_axi_m_rdata(i_l2_7_targ_ht_axi_m_rdata),
    .i_l2_7_targ_ht_axi_m_rid(i_l2_7_targ_ht_axi_m_rid),
    .i_l2_7_targ_ht_axi_m_rlast(i_l2_7_targ_ht_axi_m_rlast),
    .o_l2_7_targ_ht_axi_m_rready(o_l2_7_targ_ht_axi_m_rready),
    .i_l2_7_targ_ht_axi_m_rresp(i_l2_7_targ_ht_axi_m_rresp),
    .i_l2_7_targ_ht_axi_m_rvalid(i_l2_7_targ_ht_axi_m_rvalid),
    .o_l2_7_targ_ht_axi_m_awaddr(o_l2_7_targ_ht_axi_m_awaddr),
    .o_l2_7_targ_ht_axi_m_awburst(o_l2_7_targ_ht_axi_m_awburst),
    .o_l2_7_targ_ht_axi_m_awcache(o_l2_7_targ_ht_axi_m_awcache),
    .o_l2_7_targ_ht_axi_m_awid(o_l2_7_targ_ht_axi_m_awid),
    .o_l2_7_targ_ht_axi_m_awlen(o_l2_7_targ_ht_axi_m_awlen),
    .o_l2_7_targ_ht_axi_m_awlock(o_l2_7_targ_ht_axi_m_awlock),
    .o_l2_7_targ_ht_axi_m_awprot(o_l2_7_targ_ht_axi_m_awprot),
    .i_l2_7_targ_ht_axi_m_awready(i_l2_7_targ_ht_axi_m_awready),
    .o_l2_7_targ_ht_axi_m_awsize(o_l2_7_targ_ht_axi_m_awsize),
    .o_l2_7_targ_ht_axi_m_awvalid(o_l2_7_targ_ht_axi_m_awvalid),
    .i_l2_7_targ_ht_axi_m_bid(i_l2_7_targ_ht_axi_m_bid),
    .o_l2_7_targ_ht_axi_m_bready(o_l2_7_targ_ht_axi_m_bready),
    .i_l2_7_targ_ht_axi_m_bresp(i_l2_7_targ_ht_axi_m_bresp),
    .i_l2_7_targ_ht_axi_m_bvalid(i_l2_7_targ_ht_axi_m_bvalid),
    .o_l2_7_targ_ht_axi_m_wdata(o_l2_7_targ_ht_axi_m_wdata),
    .o_l2_7_targ_ht_axi_m_wlast(o_l2_7_targ_ht_axi_m_wlast),
    .i_l2_7_targ_ht_axi_m_wready(i_l2_7_targ_ht_axi_m_wready),
    .o_l2_7_targ_ht_axi_m_wstrb(o_l2_7_targ_ht_axi_m_wstrb),
    .o_l2_7_targ_ht_axi_m_wvalid(o_l2_7_targ_ht_axi_m_wvalid),
    .o_l2_7_targ_syscfg_apb_m_paddr(o_l2_7_targ_syscfg_apb_m_paddr),
    .o_l2_7_targ_syscfg_apb_m_penable(o_l2_7_targ_syscfg_apb_m_penable),
    .o_l2_7_targ_syscfg_apb_m_pprot(o_l2_7_targ_syscfg_apb_m_pprot),
    .i_l2_7_targ_syscfg_apb_m_prdata(i_l2_7_targ_syscfg_apb_m_prdata),
    .i_l2_7_targ_syscfg_apb_m_pready(i_l2_7_targ_syscfg_apb_m_pready),
    .o_l2_7_targ_syscfg_apb_m_psel(o_l2_7_targ_syscfg_apb_m_psel),
    .i_l2_7_targ_syscfg_apb_m_pslverr(i_l2_7_targ_syscfg_apb_m_pslverr),
    .o_l2_7_targ_syscfg_apb_m_pstrb(o_l2_7_targ_syscfg_apb_m_pstrb),
    .o_l2_7_targ_syscfg_apb_m_pwdata(o_l2_7_targ_syscfg_apb_m_pwdata),
    .o_l2_7_targ_syscfg_apb_m_pwrite(o_l2_7_targ_syscfg_apb_m_pwrite),
    .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .i_noc_clk(i_noc_clk),
    .i_noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
);

noc_tok_h_north u_noc_tok_h_north (
  .i_aic_4_clk(i_aic_4_clk),
  .i_aic_4_clken(i_aic_4_clken),
  .i_aic_4_init_tok_ocpl_s_maddr(i_aic_4_init_tok_ocpl_s_maddr),
  .i_aic_4_init_tok_ocpl_s_mcmd({{ 2'b0, i_aic_4_init_tok_ocpl_s_mcmd }}),
  .i_aic_4_init_tok_ocpl_s_mdata(i_aic_4_init_tok_ocpl_s_mdata),
  .o_aic_4_init_tok_ocpl_s_scmdaccept(o_aic_4_init_tok_ocpl_s_scmdaccept),
  .o_aic_4_pwr_tok_idle_val(o_aic_4_pwr_tok_idle_val),
  .o_aic_4_pwr_tok_idle_ack(o_aic_4_pwr_tok_idle_ack),
  .i_aic_4_pwr_tok_idle_req(i_aic_4_pwr_tok_idle_req),
  .i_aic_4_rst_n(i_aic_4_rst_n),
  .o_aic_4_targ_tok_ocpl_m_maddr(o_aic_4_targ_tok_ocpl_m_maddr),
  .o_aic_4_targ_tok_ocpl_m_mcmd(aic_4_targ_tok_ocpl_m_mcmd_ext),
  .o_aic_4_targ_tok_ocpl_m_mdata(o_aic_4_targ_tok_ocpl_m_mdata),
  .i_aic_4_targ_tok_ocpl_m_scmdaccept(i_aic_4_targ_tok_ocpl_m_scmdaccept),
  .i_aic_5_clk(i_aic_5_clk),
  .i_aic_5_clken(i_aic_5_clken),
  .i_aic_5_init_tok_ocpl_s_maddr(i_aic_5_init_tok_ocpl_s_maddr),
  .i_aic_5_init_tok_ocpl_s_mcmd({{ 2'b0, i_aic_5_init_tok_ocpl_s_mcmd }}),
  .i_aic_5_init_tok_ocpl_s_mdata(i_aic_5_init_tok_ocpl_s_mdata),
  .o_aic_5_init_tok_ocpl_s_scmdaccept(o_aic_5_init_tok_ocpl_s_scmdaccept),
  .o_aic_5_pwr_tok_idle_val(o_aic_5_pwr_tok_idle_val),
  .o_aic_5_pwr_tok_idle_ack(o_aic_5_pwr_tok_idle_ack),
  .i_aic_5_pwr_tok_idle_req(i_aic_5_pwr_tok_idle_req),
  .i_aic_5_rst_n(i_aic_5_rst_n),
  .o_aic_5_targ_tok_ocpl_m_maddr(o_aic_5_targ_tok_ocpl_m_maddr),
  .o_aic_5_targ_tok_ocpl_m_mcmd(aic_5_targ_tok_ocpl_m_mcmd_ext),
  .o_aic_5_targ_tok_ocpl_m_mdata(o_aic_5_targ_tok_ocpl_m_mdata),
  .i_aic_5_targ_tok_ocpl_m_scmdaccept(i_aic_5_targ_tok_ocpl_m_scmdaccept),
  .i_aic_6_clk(i_aic_6_clk),
  .i_aic_6_clken(i_aic_6_clken),
  .i_aic_6_init_tok_ocpl_s_maddr(i_aic_6_init_tok_ocpl_s_maddr),
  .i_aic_6_init_tok_ocpl_s_mcmd({{ 2'b0, i_aic_6_init_tok_ocpl_s_mcmd }}),
  .i_aic_6_init_tok_ocpl_s_mdata(i_aic_6_init_tok_ocpl_s_mdata),
  .o_aic_6_init_tok_ocpl_s_scmdaccept(o_aic_6_init_tok_ocpl_s_scmdaccept),
  .o_aic_6_pwr_tok_idle_val(o_aic_6_pwr_tok_idle_val),
  .o_aic_6_pwr_tok_idle_ack(o_aic_6_pwr_tok_idle_ack),
  .i_aic_6_pwr_tok_idle_req(i_aic_6_pwr_tok_idle_req),
  .i_aic_6_rst_n(i_aic_6_rst_n),
  .o_aic_6_targ_tok_ocpl_m_maddr(o_aic_6_targ_tok_ocpl_m_maddr),
  .o_aic_6_targ_tok_ocpl_m_mcmd(aic_6_targ_tok_ocpl_m_mcmd_ext),
  .o_aic_6_targ_tok_ocpl_m_mdata(o_aic_6_targ_tok_ocpl_m_mdata),
  .i_aic_6_targ_tok_ocpl_m_scmdaccept(i_aic_6_targ_tok_ocpl_m_scmdaccept),
  .i_aic_7_clk(i_aic_7_clk),
  .i_aic_7_clken(i_aic_7_clken),
  .i_aic_7_init_tok_ocpl_s_maddr(i_aic_7_init_tok_ocpl_s_maddr),
  .i_aic_7_init_tok_ocpl_s_mcmd({{ 2'b0, i_aic_7_init_tok_ocpl_s_mcmd }}),
  .i_aic_7_init_tok_ocpl_s_mdata(i_aic_7_init_tok_ocpl_s_mdata),
  .o_aic_7_init_tok_ocpl_s_scmdaccept(o_aic_7_init_tok_ocpl_s_scmdaccept),
  .o_aic_7_pwr_tok_idle_val(o_aic_7_pwr_tok_idle_val),
  .o_aic_7_pwr_tok_idle_ack(o_aic_7_pwr_tok_idle_ack),
  .i_aic_7_pwr_tok_idle_req(i_aic_7_pwr_tok_idle_req),
  .i_aic_7_rst_n(i_aic_7_rst_n),
  .o_aic_7_targ_tok_ocpl_m_maddr(o_aic_7_targ_tok_ocpl_m_maddr),
  .o_aic_7_targ_tok_ocpl_m_mcmd(aic_7_targ_tok_ocpl_m_mcmd_ext),
  .o_aic_7_targ_tok_ocpl_m_mdata(o_aic_7_targ_tok_ocpl_m_mdata),
  .i_aic_7_targ_tok_ocpl_m_scmdaccept(i_aic_7_targ_tok_ocpl_m_scmdaccept),
  .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data),
  .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head),
  .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy),
  .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail),
  .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld),
  .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data),
  .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head),
  .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy),
  .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail),
  .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld),
  .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data),
  .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head),
  .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy),
  .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail),
  .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld),
  .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data),
  .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head),
  .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy),
  .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail),
  .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld),
  .i_noc_clk(i_noc_clk),
  .i_noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en)
);
endmodule
