`ifndef GUARD_SOC_MGMT_MEMORY_MAP_APB_TEST_SV
`define GUARD_SOC_MGMT_MEMORY_MAP_APB_TEST_SV
// Extends from AI CORE soc_mgmt base test class
class soc_mgmt_memory_map_apb_test extends soc_mgmt_base_test;

  /** UVM Component Utility macro */
  `uvm_component_utils(soc_mgmt_memory_map_apb_test)
  
  bit [36-1:0] apb_addr_intr[$];
  
  int  apb_write_addr;
  int  apb_write_data;
  int loop_strt;
  int loop_len;

  apb_master_wr_rd_sequence apb_wr_rd_seq;

  // soc_mgmt user Inteface Handle
  virtual soc_mgmt_if soc_mgmt_if;

  /** Class Constructor */
  function new(string name = "soc_mgmt_memory_map_apb_test", uvm_component parent=null);
    super.new(name,parent);
  endfunction: new

  // Build Phase
  virtual function void build_phase(uvm_phase phase);
    `uvm_info("Build phase", "Entered...", UVM_LOW)
    super.build_phase(phase);


    /** Factory override of the master transaction object */
    set_type_override_by_type (svt_axi_master_transaction::get_type(), cust_svt_axi_master_transaction::get_type());

    `uvm_info("build_phase", "Loaded cust_svt_axi_system_configuration ", UVM_LOW)

    // random selection of slave response normal or zero delay sequence
    apb_wr_rd_seq	= apb_master_wr_rd_sequence::type_id::create("apb_wr_rd_seq");

    // Recieve soc_mgmt user interface handle
    uvm_config_db#(virtual soc_mgmt_if)::get(
        uvm_root::get(), "uvm_test_top", "soc_mgmt_if", soc_mgmt_if);

    `uvm_info("build_phase", "Exiting...", UVM_LOW)
  endfunction: build_phase

  virtual task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    
    `uvm_info("base_test:run_phase", "Entered...", UVM_LOW)

    
    if ($value$plusargs ("LOOP_STRT=%d", loop_strt))
      `uvm_info("SOC_MGMT_APB",$sformatf("value of loop_start is %d",loop_strt ), UVM_LOW)
    else loop_strt=0;

    if ($value$plusargs ("LOOP_LEN=%d", loop_len))
      `uvm_info("SOC_MGMT_APB",$sformatf("value of loop_len is  %d",loop_len ), UVM_LOW)
    else loop_len=2;
    
    `uvm_info("SOC_MGMT_APB",$sformatf("value of loop_start is %0d and loop_len is %d",loop_strt, loop_len ), UVM_LOW)

    // Address and data
    `uvm_info("SOC_MGMT_APB_LP",$sformatf("Entered into running phase"), UVM_LOW)
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_CLOCK_GEN_CSR_ST_ADDR);
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_CLOCK_GEN_CSR_END_ADDR - 8);
    
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_RESET_GEN_CSR_ST_ADDR);
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_RESET_GEN_CSR_END_ADDR - 8);
    
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_NOC_AO_CSR_ST_ADDR);
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_NOC_AO_CSR_END_ADDR - 8);
    
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_MISC_AO_CSR_ST_ADDR);
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_MISC_AO_CSR_END_ADDR - 8);
    
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_DLM_CSR_ST_ADDR);
    apb_addr_intr.push_back(soc_mgmt_common_pkg::SYS_CFG_SOC_MGMT_AO_CSR_DLM_CSR_END_ADDR - 8);


    @(posedge soc_mgmt_if.o_ao_rst_n);
    `uvm_info("SOC_MGMT_APB",$sformatf("introducing delay .. "), UVM_LOW)
    #100;
    `uvm_info("SOC_MGMT_APB",$sformatf("after delay .. "), UVM_LOW)

    for (int i =loop_strt;i<loop_len;i++) begin
        apb_wr_rd_seq.randomize() with {
        cfg_addr        == apb_addr_intr[i]; // pctl_ao_csr_reg_ppmu_reset_control
        cfg_data        == 'hFFFF_FFFF;
        };
        // Start the sequence on the respective sequencer
       apb_wr_rd_seq.start(env.apb_master_env.master.sequencer);  //apb_master_env.master.sequencer.apb_master_wr_rd_sequence
       `uvm_info("SOC_MGMT_AXI",$sformatf("sequence ended for addr %0h",apb_addr_intr[i] ), UVM_LOW)
    end

    `uvm_info("base_test:run_phase", "Exiting...", UVM_LOW)
    phase.drop_objection(this);
  endtask

endclass:soc_mgmt_memory_map_apb_test

`endif // GUARD_SOC_MGMT_MEMORY_MAP_APB_TEST_SV
