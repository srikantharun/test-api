`ifndef TEST_PKG_SV
`define TEST_PKG_SV

package test_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import axe_uvm_resource_allocator_pkg::*;

  `include "test.svh"

endpackage : test_pkg

`endif // TEST_PKG_SV
