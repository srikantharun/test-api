// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: Andrew Dickson <andrew.dickson@axelera.ai>

/// Generic PVT Probe Wrapper IP containing the instance of the PVT Probe
/// Used for compilation only.

module tu_tem0501ar01_ln05lpe_4007002 #(
)
(
  // Probe VSS
  inout logic AVSS_TS  , 
  // Probe GND
  inout logic AVSS_GD  , 
  // Probe IBias
  inout logic IBIAS_TS , 
  // Probe VSense
  inout logic VSENSE_TS
);

endmodule
