module axe_ax65_cluster
  import apu_pkg::*;
#(
    parameter int unsigned CORE_WIDTH = 6,
    parameter int unsigned MAX_CORE_WIDTH = 8,
    parameter int unsigned BHT_WIDTH = 7,
    parameter int unsigned DCACHE_WIDTH = 16,
    parameter int unsigned ICACHE_WIDTH = 8,
    parameter int unsigned L2_WIDTH = 4,
    parameter int unsigned L2C_BANK_WIDTH = 4,
    parameter int unsigned L2C_BANK_DATA_WIDTH = 8,
    parameter int unsigned L2C_BANK_TAG_WIDTH = 64,
    parameter int unsigned SINK_WIDTH = 6,
    parameter int unsigned SOURCE_WIDTH = 5,
    parameter int unsigned CTRL_IN_WIDTH = 9,
    parameter int unsigned CTRL_OUT_WIDTH = 1
) (
    /// Slow ref clock
    input wire i_mtime_clk,
    input wire i_por_rst_n,
    /// Fast core clocks
    input wire [CORE_WIDTH - 1:0] i_cores_clk,
    input wire [CORE_WIDTH - 1:0] i_cores_rst_n,
    /// Fast AXI clock
    input wire i_aclk,
    input wire i_arst_n,
    /// Fast l2 clock
    input wire i_l2c_clk,
    input wire i_l2c_rst_n,

    //////////////////////////////////////////////
    /// COREs sigs
    //////////////////////////////////////////////
    input  axe_tcl_sram_pkg::impl_inp_t [CORE_WIDTH - 1:0] i_cores_ctrl,
    output axe_tcl_sram_pkg::impl_oup_t [CORE_WIDTH - 1:0] o_cores_ctrl,
    input logic [CORE_WIDTH - 1:0] i_cores_disable_init,
    input logic [CORE_WIDTH - 1:0][63:0] i_cores_hart_id,
    input logic [CORE_WIDTH - 1:0] i_cores_meip,
    input logic [CORE_WIDTH - 1:0] i_cores_msip,
    input logic [CORE_WIDTH - 1:0] i_cores_nmi,
    input logic [CORE_WIDTH - 1:0][47:0] i_cores_reset_vector,
    input logic [CORE_WIDTH - 1:0] i_cores_seip,
    output logic [CORE_WIDTH - 1:0] o_cores_wfi_mode,
    /// Debug sigs
    input logic [CORE_WIDTH - 1:0] i_cores_debugint,
    input logic [CORE_WIDTH - 1:0] i_cores_resethaltreq,
    output logic [CORE_WIDTH - 1:0] o_cores_hart_unavail,
    output logic [CORE_WIDTH - 1:0] o_cores_hart_under_reset,

    //////////////////////////////////////////////
    /// AXIs sigs
    //////////////////////////////////////////////
    // IOCP
    input ax65_axi_lt_s_aw_t i_iocp_axi_s_aw,
    output logic o_iocp_axi_s_awready,
    input logic i_iocp_axi_s_awvalid,
    input ax65_axi_lt_w_t i_iocp_axi_s_w,
    output logic o_iocp_axi_s_wready,
    input logic i_iocp_axi_s_wvalid,
    output ax65_axi_lt_s_b_t o_iocp_axi_s_b,
    input logic i_iocp_axi_s_bready,
    output logic o_iocp_axi_s_bvalid,
    input ax65_axi_lt_s_ar_t i_iocp_axi_s_ar,
    output logic o_iocp_axi_s_arready,
    input logic i_iocp_axi_s_arvalid,
    output ax65_axi_lt_s_r_t o_iocp_axi_s_r,
    input logic i_iocp_axi_s_rready,
    output logic o_iocp_axi_s_rvalid,
    // MEM
    output ax65_axi_mt_m_aw_t o_mem_axi_m_aw,
    input logic i_mem_axi_m_awready,
    output logic o_mem_axi_m_awvalid,
    output apu_axi_mt_w_t o_mem_axi_m_w,
    input logic i_mem_axi_m_wready,
    output logic o_mem_axi_m_wvalid,
    input ax65_axi_mt_m_b_t i_mem_axi_m_b,
    output logic o_mem_axi_m_bready,
    input logic i_mem_axi_m_bvalid,
    output ax65_axi_mt_m_ar_t o_mem_axi_m_ar,
    input logic i_mem_axi_m_arready,
    output logic o_mem_axi_m_arvalid,
    input ax65_axi_mt_m_r_t i_mem_axi_m_r,
    output logic o_mem_axi_m_rready,
    input logic i_mem_axi_m_rvalid,
    // MMIO
    output apu_axi_lt_m_aw_t o_mmio_axi_m_aw,
    input logic i_mmio_axi_m_awready,
    output logic o_mmio_axi_m_awvalid,
    output apu_axi_lt_w_t o_mmio_axi_m_w,
    input logic i_mmio_axi_m_wready,
    output logic o_mmio_axi_m_wvalid,
    input apu_axi_lt_m_b_t i_mmio_axi_m_b,
    output logic o_mmio_axi_m_bready,
    input logic i_mmio_axi_m_bvalid,
    output apu_axi_lt_m_ar_t o_mmio_axi_m_ar,
    input logic i_mmio_axi_m_arready,
    output logic o_mmio_axi_m_arvalid,
    input apu_axi_lt_m_r_t i_mmio_axi_m_r,
    output logic o_mmio_axi_m_rready,
    input logic i_mmio_axi_m_rvalid,

    //////////////////////////////////////////////
    /// L2 sigs
    //////////////////////////////////////////////
    input  axe_tcl_sram_pkg::impl_inp_t i_l2c_ctrl,
    output axe_tcl_sram_pkg::impl_oup_t o_l2c_ctrl,
    input logic i_l2c_disable_init,
    output logic o_l2c_err_int,

    //////////////////////////////////////////////
    /// Misc sigs
    //////////////////////////////////////////////
    output logic [APU_AIC_WIDTH - 1:0] o_aic_mtip,
    input  logic [APU_AIC_WIDTH - 1:0] i_aic_stoptime,
    input logic i_test_mode
);

  logic [CORE_WIDTH + APU_AIC_WIDTH - 1:0] all_cores_mtip;
  logic [CORE_WIDTH + APU_AIC_WIDTH - 1:0] all_cores_stoptime;
  logic [CORE_WIDTH - 1:0] cores_mtip;
  logic [CORE_WIDTH - 1:0] cores_stoptime;
  logic [CORE_WIDTH - 1:0] cores_wfi_mode;

  always_comb o_aic_mtip = all_cores_mtip[CORE_WIDTH + APU_AIC_WIDTH - 1:CORE_WIDTH];
  always_comb cores_mtip = all_cores_mtip[CORE_WIDTH - 1:0];
  always_comb o_cores_wfi_mode = cores_wfi_mode;

  always_comb all_cores_stoptime[CORE_WIDTH + APU_AIC_WIDTH - 1:CORE_WIDTH] = i_aic_stoptime;
  always_comb all_cores_stoptime[CORE_WIDTH - 1:0] = cores_stoptime;

  logic [CORE_WIDTH - 1:0] cores_coherent_state;
  logic [CORE_WIDTH - 1:0] cores_coherent_enable;
  logic [CORE_WIDTH - 1:0][39:0] cores_dcu_a_address;
  logic [CORE_WIDTH - 1:0] cores_dcu_a_corrupt;
  logic [CORE_WIDTH - 1:0][255:0] cores_dcu_a_data;
  logic [CORE_WIDTH - 1:0][31:0] cores_dcu_a_mask;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_a_opcode;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_a_param;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_a_size;
  logic [CORE_WIDTH - 1:0][SOURCE_WIDTH - 1:0] cores_dcu_a_source;
  logic [CORE_WIDTH - 1:0][11:0] cores_dcu_a_user;
  logic [CORE_WIDTH - 1:0] cores_dcu_a_ready;
  logic [CORE_WIDTH - 1:0] cores_dcu_a_valid;
  logic [CORE_WIDTH - 1:0][39:0] cores_dcu_b_address;
  logic [CORE_WIDTH - 1:0] cores_dcu_b_corrupt;
  logic [CORE_WIDTH - 1:0][255:0] cores_dcu_b_data;
  logic [CORE_WIDTH - 1:0][31:0] cores_dcu_b_mask;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_b_opcode;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_b_param;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_b_size;
  logic [CORE_WIDTH - 1:0][SOURCE_WIDTH - 1:0] cores_dcu_b_source;
  logic [CORE_WIDTH - 1:0] cores_dcu_b_ready;
  logic [CORE_WIDTH - 1:0] cores_dcu_b_valid;
  logic [CORE_WIDTH - 1:0][39:0] cores_dcu_c_address;
  logic [CORE_WIDTH - 1:0] cores_dcu_c_corrupt;
  logic [CORE_WIDTH - 1:0][255:0] cores_dcu_c_data;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_c_opcode;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_c_param;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_c_size;
  logic [CORE_WIDTH - 1:0][SOURCE_WIDTH - 1:0] cores_dcu_c_source;
  logic [CORE_WIDTH - 1:0][7:0] cores_dcu_c_user;
  logic [CORE_WIDTH - 1:0] cores_dcu_c_ready;
  logic [CORE_WIDTH - 1:0] cores_dcu_c_valid;
  logic [CORE_WIDTH - 1:0] cores_dcu_d_corrupt;
  logic [CORE_WIDTH - 1:0][255:0] cores_dcu_d_data;
  logic [CORE_WIDTH - 1:0] cores_dcu_d_denied;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_d_opcode;
  logic [CORE_WIDTH - 1:0][1:0] cores_dcu_d_param;
  logic [CORE_WIDTH - 1:0][2:0] cores_dcu_d_size;
  logic [CORE_WIDTH - 1:0][SINK_WIDTH - 1:0] cores_dcu_d_sink;
  logic [CORE_WIDTH - 1:0][SOURCE_WIDTH - 1:0] cores_dcu_d_source;
  logic [CORE_WIDTH - 1:0][5:0] cores_dcu_d_user;
  logic [CORE_WIDTH - 1:0] cores_dcu_d_ready;
  logic [CORE_WIDTH - 1:0] cores_dcu_d_valid;
  logic [CORE_WIDTH - 1:0][SINK_WIDTH - 1:0] cores_dcu_e_sink;
  logic [CORE_WIDTH - 1:0] cores_dcu_e_ready;
  logic [CORE_WIDTH - 1:0] cores_dcu_e_valid;
  logic [CORE_WIDTH - 1:0][39:0] cores_icu_a_address;
  logic [CORE_WIDTH - 1:0] cores_icu_a_corrupt;
  logic [CORE_WIDTH - 1:0][255:0] cores_icu_a_data;
  logic [CORE_WIDTH - 1:0][31:0] cores_icu_a_mask;
  logic [CORE_WIDTH - 1:0][2:0] cores_icu_a_opcode;
  logic [CORE_WIDTH - 1:0][2:0] cores_icu_a_param;
  logic [CORE_WIDTH - 1:0][2:0] cores_icu_a_size;
  logic [CORE_WIDTH - 1:0][SOURCE_WIDTH - 1:0] cores_icu_a_source;
  logic [CORE_WIDTH - 1:0][11:0] cores_icu_a_user;
  logic [CORE_WIDTH - 1:0] cores_icu_a_ready;
  logic [CORE_WIDTH - 1:0] cores_icu_a_valid;
  logic [CORE_WIDTH - 1:0] cores_icu_d_corrupt;
  logic [CORE_WIDTH - 1:0][255:0] cores_icu_d_data;
  logic [CORE_WIDTH - 1:0] cores_icu_d_denied;
  logic [CORE_WIDTH - 1:0][2:0] cores_icu_d_opcode;
  logic [CORE_WIDTH - 1:0][1:0] cores_icu_d_param;
  logic [CORE_WIDTH - 1:0][2:0] cores_icu_d_size;
  logic [CORE_WIDTH - 1:0][SINK_WIDTH - 1:0] cores_icu_d_sink;
  logic [CORE_WIDTH - 1:0][SOURCE_WIDTH - 1:0] cores_icu_d_source;
  logic [CORE_WIDTH - 1:0][5:0] cores_icu_d_user;
  logic [CORE_WIDTH - 1:0] cores_icu_d_ready;
  logic [CORE_WIDTH - 1:0] cores_icu_d_valid;
  logic [CORE_WIDTH - 1:0][39:0] cores_mpipe_axi_araddr;
  logic [CORE_WIDTH - 1:0][1:0] cores_mpipe_axi_arburst;
  logic [CORE_WIDTH - 1:0][3:0] cores_mpipe_axi_arcache;
  logic [CORE_WIDTH - 1:0][4:0] cores_mpipe_axi_arid;
  logic [CORE_WIDTH - 1:0][7:0] cores_mpipe_axi_arlen;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_arlock;
  logic [CORE_WIDTH - 1:0][2:0] cores_mpipe_axi_arprot;
  logic [CORE_WIDTH - 1:0][2:0] cores_mpipe_axi_arsize;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_arready;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_arvalid;
  logic [CORE_WIDTH - 1:0][39:0] cores_mpipe_axi_awaddr;
  logic [CORE_WIDTH - 1:0][1:0] cores_mpipe_axi_awburst;
  logic [CORE_WIDTH - 1:0][3:0] cores_mpipe_axi_awcache;
  logic [CORE_WIDTH - 1:0][4:0] cores_mpipe_axi_awid;
  logic [CORE_WIDTH - 1:0][7:0] cores_mpipe_axi_awlen;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_awlock;
  logic [CORE_WIDTH - 1:0][2:0] cores_mpipe_axi_awprot;
  logic [CORE_WIDTH - 1:0][2:0] cores_mpipe_axi_awsize;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_awready;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_awvalid;
  logic [CORE_WIDTH - 1:0][4:0] cores_mpipe_axi_bid;
  logic [CORE_WIDTH - 1:0][1:0] cores_mpipe_axi_bresp;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_bready;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_bvalid;
  logic [CORE_WIDTH - 1:0][63:0] cores_mpipe_axi_rdata;
  logic [CORE_WIDTH - 1:0][4:0] cores_mpipe_axi_rid;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_rlast;
  logic [CORE_WIDTH - 1:0][1:0] cores_mpipe_axi_rresp;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_rready;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_rvalid;
  logic [CORE_WIDTH - 1:0][63:0] cores_mpipe_axi_wdata;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_wlast;
  logic [CORE_WIDTH - 1:0][(64 / 8) - 1:0] cores_mpipe_axi_wstrb;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_wready;
  logic [CORE_WIDTH - 1:0] cores_mpipe_axi_wvalid;

  // DS_CORES
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_coherent_enable;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_coherent_state;
  logic [MAX_CORE_WIDTH - 1:0][((40) - 1):0] ds_cores_m0_a_address;
  logic [MAX_CORE_WIDTH - 1:0][0:0] ds_cores_m0_a_corrupt;
  logic [MAX_CORE_WIDTH - 1:0][((256) - 1):0] ds_cores_m0_a_data;
  logic [MAX_CORE_WIDTH - 1:0][(256) / 8 - 1:0] ds_cores_m0_a_mask;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_a_opcode;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_a_param;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_a_size;
  logic [MAX_CORE_WIDTH - 1:0][(SOURCE_WIDTH - 1):0] ds_cores_m0_a_source;
  logic [MAX_CORE_WIDTH - 1:0][11:0] ds_cores_m0_a_user;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_a_valid;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_b_ready;
  logic [MAX_CORE_WIDTH - 1:0][((40) - 1):0] ds_cores_m0_c_address;
  logic [MAX_CORE_WIDTH - 1:0][0:0] ds_cores_m0_c_corrupt;
  logic [MAX_CORE_WIDTH - 1:0][((256) - 1):0] ds_cores_m0_c_data;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_c_opcode;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_c_param;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_c_size;
  logic [MAX_CORE_WIDTH - 1:0][(SOURCE_WIDTH - 1):0] ds_cores_m0_c_source;
  logic [MAX_CORE_WIDTH - 1:0][7:0] ds_cores_m0_c_user;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_c_valid;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_d_ready;
  logic [MAX_CORE_WIDTH - 1:0][(SINK_WIDTH - 1):0] ds_cores_m0_e_sink;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_e_valid;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_a_ready;
  logic [MAX_CORE_WIDTH - 1:0][((40) - 1):0] ds_cores_m0_b_address;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_b_corrupt;
  logic [MAX_CORE_WIDTH - 1:0][((256) - 1):0] ds_cores_m0_b_data;
  logic [MAX_CORE_WIDTH - 1:0][((256) / 8) - 1:0] ds_cores_m0_b_mask;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_b_opcode;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_b_param;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_b_size;
  logic [MAX_CORE_WIDTH - 1:0][(SOURCE_WIDTH - 1):0] ds_cores_m0_b_source;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_b_valid;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_c_ready;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_d_corrupt;
  logic [MAX_CORE_WIDTH - 1:0][((256) - 1):0] ds_cores_m0_d_data;
  logic [MAX_CORE_WIDTH - 1:0][0:0] ds_cores_m0_d_denied;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_d_opcode;
  logic [MAX_CORE_WIDTH - 1:0][1:0] ds_cores_m0_d_param;
  logic [MAX_CORE_WIDTH - 1:0][(SINK_WIDTH - 1):0] ds_cores_m0_d_sink;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m0_d_size;
  logic [MAX_CORE_WIDTH - 1:0][(SOURCE_WIDTH - 1):0] ds_cores_m0_d_source;
  logic [MAX_CORE_WIDTH - 1:0][5:0] ds_cores_m0_d_user;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_d_valid;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m0_e_ready;
  logic [MAX_CORE_WIDTH - 1:0][39:0] ds_cores_m1_axi_araddr;
  logic [MAX_CORE_WIDTH - 1:0][1:0] ds_cores_m1_axi_arburst;
  logic [MAX_CORE_WIDTH - 1:0][3:0] ds_cores_m1_axi_arcache;
  logic [MAX_CORE_WIDTH - 1:0][4:0] ds_cores_m1_axi_arid;
  logic [MAX_CORE_WIDTH - 1:0][7:0] ds_cores_m1_axi_arlen;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_arlock;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m1_axi_arprot;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m1_axi_arsize;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_arready;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_arvalid;
  logic [MAX_CORE_WIDTH - 1:0][39:0] ds_cores_m1_axi_awaddr;
  logic [MAX_CORE_WIDTH - 1:0][1:0] ds_cores_m1_axi_awburst;
  logic [MAX_CORE_WIDTH - 1:0][3:0] ds_cores_m1_axi_awcache;
  logic [MAX_CORE_WIDTH - 1:0][4:0] ds_cores_m1_axi_awid;
  logic [MAX_CORE_WIDTH - 1:0][7:0] ds_cores_m1_axi_awlen;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_awlock;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m1_axi_awprot;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m1_axi_awsize;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_awready;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_awvalid;
  logic [MAX_CORE_WIDTH - 1:0][4:0] ds_cores_m1_axi_bid;
  logic [MAX_CORE_WIDTH - 1:0][1:0] ds_cores_m1_axi_bresp;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_bready;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_bvalid;
  logic [MAX_CORE_WIDTH - 1:0][63:0] ds_cores_m1_axi_rdata;
  logic [MAX_CORE_WIDTH - 1:0][4:0] ds_cores_m1_axi_rid;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_rlast;
  logic [MAX_CORE_WIDTH - 1:0][1:0] ds_cores_m1_axi_rresp;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_rready;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_rvalid;
  logic [MAX_CORE_WIDTH - 1:0][63:0] ds_cores_m1_axi_wdata;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_wlast;
  logic [MAX_CORE_WIDTH - 1:0][(64 / 8) -1:0] ds_cores_m1_axi_wstrb;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_wready;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m1_axi_wvalid;
  logic [MAX_CORE_WIDTH - 1:0][((40) - 1):0] ds_cores_m2_a_address;
  logic [MAX_CORE_WIDTH - 1:0][0:0] ds_cores_m2_a_corrupt;
  logic [MAX_CORE_WIDTH - 1:0][((256) - 1):0] ds_cores_m2_a_data;
  logic [MAX_CORE_WIDTH - 1:0][(256) / 8 - 1:0] ds_cores_m2_a_mask;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m2_a_opcode;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m2_a_param;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m2_a_size;
  logic [MAX_CORE_WIDTH - 1:0][(SOURCE_WIDTH - 1):0] ds_cores_m2_a_source;
  logic [MAX_CORE_WIDTH - 1:0][11:0] ds_cores_m2_a_user;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m2_a_valid;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m2_d_ready;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m2_a_ready;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m2_d_corrupt;
  logic [MAX_CORE_WIDTH - 1:0][((256) - 1):0] ds_cores_m2_d_data;
  logic [MAX_CORE_WIDTH - 1:0][0:0] ds_cores_m2_d_denied;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m2_d_opcode;
  logic [MAX_CORE_WIDTH - 1:0][1:0] ds_cores_m2_d_param;
  logic [MAX_CORE_WIDTH - 1:0][(SINK_WIDTH - 1):0] ds_cores_m2_d_sink;
  logic [MAX_CORE_WIDTH - 1:0][2:0] ds_cores_m2_d_size;
  logic [MAX_CORE_WIDTH - 1:0][(SOURCE_WIDTH - 1):0] ds_cores_m2_d_source;
  logic [MAX_CORE_WIDTH - 1:0][5:0] ds_cores_m2_d_user;
  logic [MAX_CORE_WIDTH - 1:0] ds_cores_m2_d_valid;

  apu_axi_lt_m_ar_t plmt_axi_ar;
  logic plmt_axi_arready;
  logic plmt_axi_arvalid;
  apu_axi_lt_m_aw_t plmt_axi_aw;
  logic plmt_axi_awready;
  logic plmt_axi_awvalid;
  apu_axi_lt_m_b_t plmt_axi_b;
  logic plmt_axi_bready;
  logic plmt_axi_bvalid;
  apu_axi_lt_m_r_t plmt_axi_r;
  logic plmt_axi_rready;
  logic plmt_axi_rvalid;
  apu_axi_lt_w_t plmt_axi_w;
  logic plmt_axi_wready;
  logic plmt_axi_wvalid;

  /// Fast core clocks
  wire [CORE_WIDTH - 1:0] cores_clk;
  wire [CORE_WIDTH - 1:0] cores_dcu_clk;
  /// Enable sigs for apu_core_p
  logic [CORE_WIDTH - 1:0] cores_clk_enable;
  logic [CORE_WIDTH - 1:0] cores_dcu_clk_enable;
  /// Fast l2c clock
  wire l2c_clk;
  /// Div2 l2c clock
  wire l2c_banks_clk;
  wire l2c_banks_clk_en;

  apu_cluster_power_management_unit #(
    .CORE_WIDTH(CORE_WIDTH),
    .SYNC_STAGES(3),
    .PIPELINE_STAGES(1)
  ) u_apu_pmu (
    /// Fast core clocks
    .i_cores_clk(i_cores_clk),
    .i_cores_rst_n(i_cores_rst_n),
    /// Fast l2c clock
    .i_l2c_clk(i_l2c_clk),
    .i_l2c_rst_n(i_l2c_rst_n),

    /// Fast core clocks
    .o_cores_clk(cores_clk),
    .o_cores_dcu_clk(cores_dcu_clk),
    /// Enable sigs for apu_core_p
    .o_cores_clk_enable(cores_clk_enable),
    .o_cores_dcu_clk_enable(cores_dcu_clk_enable),
    /// Fast l2c clock
    .o_l2c_clk(l2c_clk),
    /// Div2 l2c clock
    .o_l2c_banks_clk(l2c_banks_clk),
    .o_l2c_banks_clk_en(l2c_banks_clk_en),

    /// DFT
    .i_test_en('0),

    /// internal state
    .i_cores_wfi_mode(cores_wfi_mode),
    .i_cores_debugint(i_cores_debugint),
    .i_cores_nmi(i_cores_nmi),
    .i_cores_meip(i_cores_meip),
    .i_cores_seip(i_cores_seip),
    .i_cores_msip(i_cores_msip),
    .i_cores_mtip(cores_mtip),
    .i_cores_coherent_state(cores_coherent_state),
    .i_cores_coherent_enable(cores_coherent_enable)
  );

  for (genvar i = 0; unsigned'(i) < CORE_WIDTH; i++) begin: g_cores
    apu_core_p u_core_p (
      .i_clk(i_cores_clk[i]),
      .i_rst_n(i_cores_rst_n[i]),

      // Core clocks management
      .i_core_clk_enable(cores_clk_enable[i]),
      .i_core_dcu_clk_enable(cores_dcu_clk_enable[i]),

      // JTAG
      .ijtag_tck('0),
      .ijtag_reset('0),
      .ijtag_sel('0),
      .ijtag_ue('0),
      .ijtag_se('0),
      .ijtag_ce('0),
      .ijtag_si('0),
      .ijtag_so(),
      // DFT
      .test_clk('0),
      .test_mode('0),
      .edt_update('0),
      .scan_en('0),
      .scan_in('0),
      .scan_out(),
      // BIST
      .bisr_clk('0),
      .bisr_reset('0),
      .bisr_shift_en('0),
      .bisr_si('0),
      .bisr_so(),

      //////////////////////////////////////////////
      /// CORE sigs
      //////////////////////////////////////////////
      .i_coherent_state(cores_coherent_state[i]),
      .o_coherent_enable(cores_coherent_enable[i]),
      .o_wfi_mode(cores_wfi_mode[i]),
      .o_dcu_a_address(cores_dcu_a_address[i]),
      .o_dcu_a_corrupt(cores_dcu_a_corrupt[i]),
      .o_dcu_a_data(cores_dcu_a_data[i]),
      .o_dcu_a_mask(cores_dcu_a_mask[i]),
      .o_dcu_a_opcode(cores_dcu_a_opcode[i]),
      .o_dcu_a_param(cores_dcu_a_param[i]),
      .o_dcu_a_size(cores_dcu_a_size[i]),
      .o_dcu_a_source(cores_dcu_a_source[i]),
      .o_dcu_a_user(cores_dcu_a_user[i]),
      .i_dcu_a_ready(cores_dcu_a_ready[i]),
      .o_dcu_a_valid(cores_dcu_a_valid[i]),
      .i_dcu_b_address(cores_dcu_b_address[i]),
      .i_dcu_b_corrupt(cores_dcu_b_corrupt[i]),
      .i_dcu_b_data(cores_dcu_b_data[i]),
      .i_dcu_b_mask(cores_dcu_b_mask[i]),
      .i_dcu_b_opcode(cores_dcu_b_opcode[i]),
      .i_dcu_b_param(cores_dcu_b_param[i]),
      .i_dcu_b_size(cores_dcu_b_size[i]),
      .i_dcu_b_source(cores_dcu_b_source[i]),
      .o_dcu_b_ready(cores_dcu_b_ready[i]),
      .i_dcu_b_valid(cores_dcu_b_valid[i]),
      .o_dcu_c_address(cores_dcu_c_address[i]),
      .o_dcu_c_corrupt(cores_dcu_c_corrupt[i]),
      .o_dcu_c_data(cores_dcu_c_data[i]),
      .o_dcu_c_opcode(cores_dcu_c_opcode[i]),
      .o_dcu_c_param(cores_dcu_c_param[i]),
      .o_dcu_c_size(cores_dcu_c_size[i]),
      .o_dcu_c_source(cores_dcu_c_source[i]),
      .o_dcu_c_user(cores_dcu_c_user[i]),
      .i_dcu_c_ready(cores_dcu_c_ready[i]),
      .o_dcu_c_valid(cores_dcu_c_valid[i]),
      .i_dcu_d_corrupt(cores_dcu_d_corrupt[i]),
      .i_dcu_d_data(cores_dcu_d_data[i]),
      .i_dcu_d_denied(cores_dcu_d_denied[i]),
      .i_dcu_d_opcode(cores_dcu_d_opcode[i]),
      .i_dcu_d_param(cores_dcu_d_param[i]),
      .i_dcu_d_size(cores_dcu_d_size[i]),
      .i_dcu_d_sink(cores_dcu_d_sink[i]),
      .i_dcu_d_source(cores_dcu_d_source[i]),
      .i_dcu_d_user(cores_dcu_d_user[i]),
      .o_dcu_d_ready(cores_dcu_d_ready[i]),
      .i_dcu_d_valid(cores_dcu_d_valid[i]),
      .o_dcu_e_sink(cores_dcu_e_sink[i]),
      .i_dcu_e_ready(cores_dcu_e_ready[i]),
      .o_dcu_e_valid(cores_dcu_e_valid[i]),
      .o_icu_a_address(cores_icu_a_address[i]),
      .o_icu_a_corrupt(cores_icu_a_corrupt[i]),
      .o_icu_a_data(cores_icu_a_data[i]),
      .o_icu_a_mask(cores_icu_a_mask[i]),
      .o_icu_a_opcode(cores_icu_a_opcode[i]),
      .o_icu_a_param(cores_icu_a_param[i]),
      .o_icu_a_size(cores_icu_a_size[i]),
      .o_icu_a_source(cores_icu_a_source[i]),
      .o_icu_a_user(cores_icu_a_user[i]),
      .i_icu_a_ready(cores_icu_a_ready[i]),
      .o_icu_a_valid(cores_icu_a_valid[i]),
      .i_icu_d_corrupt(cores_icu_d_corrupt[i]),
      .i_icu_d_data(cores_icu_d_data[i]),
      .i_icu_d_denied(cores_icu_d_denied[i]),
      .i_icu_d_opcode(cores_icu_d_opcode[i]),
      .i_icu_d_param(cores_icu_d_param[i]),
      .i_icu_d_size(cores_icu_d_size[i]),
      .i_icu_d_sink(cores_icu_d_sink[i]),
      .i_icu_d_source(cores_icu_d_source[i]),
      .i_icu_d_user(cores_icu_d_user[i]),
      .o_icu_d_ready(cores_icu_d_ready[i]),
      .i_icu_d_valid(cores_icu_d_valid[i]),
      .o_mpipe_axi_m_araddr(cores_mpipe_axi_araddr[i]),
      .o_mpipe_axi_m_arburst(cores_mpipe_axi_arburst[i]),
      .o_mpipe_axi_m_arcache(cores_mpipe_axi_arcache[i]),
      .o_mpipe_axi_m_arid(cores_mpipe_axi_arid[i]),
      .o_mpipe_axi_m_arlen(cores_mpipe_axi_arlen[i]),
      .o_mpipe_axi_m_arlock(cores_mpipe_axi_arlock[i]),
      .o_mpipe_axi_m_arprot(cores_mpipe_axi_arprot[i]),
      .o_mpipe_axi_m_arsize(cores_mpipe_axi_arsize[i]),
      .i_mpipe_axi_m_arready(cores_mpipe_axi_arready[i]),
      .o_mpipe_axi_m_arvalid(cores_mpipe_axi_arvalid[i]),
      .o_mpipe_axi_m_awaddr(cores_mpipe_axi_awaddr[i]),
      .o_mpipe_axi_m_awburst(cores_mpipe_axi_awburst[i]),
      .o_mpipe_axi_m_awcache(cores_mpipe_axi_awcache[i]),
      .o_mpipe_axi_m_awid(cores_mpipe_axi_awid[i]),
      .o_mpipe_axi_m_awlen(cores_mpipe_axi_awlen[i]),
      .o_mpipe_axi_m_awlock(cores_mpipe_axi_awlock[i]),
      .o_mpipe_axi_m_awprot(cores_mpipe_axi_awprot[i]),
      .o_mpipe_axi_m_awsize(cores_mpipe_axi_awsize[i]),
      .i_mpipe_axi_m_awready(cores_mpipe_axi_awready[i]),
      .o_mpipe_axi_m_awvalid(cores_mpipe_axi_awvalid[i]),
      .i_mpipe_axi_m_bid(cores_mpipe_axi_bid[i]),
      .i_mpipe_axi_m_bresp(cores_mpipe_axi_bresp[i]),
      .o_mpipe_axi_m_bready(cores_mpipe_axi_bready[i]),
      .i_mpipe_axi_m_bvalid(cores_mpipe_axi_bvalid[i]),
      .i_mpipe_axi_m_rdata(cores_mpipe_axi_rdata[i]),
      .i_mpipe_axi_m_rid(cores_mpipe_axi_rid[i]),
      .i_mpipe_axi_m_rlast(cores_mpipe_axi_rlast[i]),
      .i_mpipe_axi_m_rresp(cores_mpipe_axi_rresp[i]),
      .o_mpipe_axi_m_rready(cores_mpipe_axi_rready[i]),
      .i_mpipe_axi_m_rvalid(cores_mpipe_axi_rvalid[i]),
      .o_mpipe_axi_m_wdata(cores_mpipe_axi_wdata[i]),
      .o_mpipe_axi_m_wlast(cores_mpipe_axi_wlast[i]),
      .o_mpipe_axi_m_wstrb(cores_mpipe_axi_wstrb[i]),
      .i_mpipe_axi_m_wready(cores_mpipe_axi_wready[i]),
      .o_mpipe_axi_m_wvalid(cores_mpipe_axi_wvalid[i]),
      .i_dcache_disable_init(i_cores_disable_init[i]),
      .i_icache_disable_init(i_cores_disable_init[i]),
      .i_debugint(i_cores_debugint[i]),
      .i_hart_id(i_cores_hart_id[i]),
      .o_hart_unavail(o_cores_hart_unavail[i]),
      .o_hart_under_reset(o_cores_hart_under_reset[i]),
      .i_meip(i_cores_meip[i]),
      .i_msip(i_cores_msip[i]),
      .i_mtip(cores_mtip[i]),
      .i_nmi(i_cores_nmi[i]),
      .i_reset_vector(i_cores_reset_vector[i]),
      .i_resethaltreq(i_cores_resethaltreq[i]),
      .i_seip(i_cores_seip[i]),
      .o_stoptime(cores_stoptime[i]),
      .i_core_ctrl(i_cores_ctrl[i]),
      .o_core_ctrl(o_cores_ctrl[i])
    );
  end: g_cores

  ax65_bridge_wrapper #(
    .CORE_WIDTH(CORE_WIDTH),
    .MAX_CORE_WIDTH(MAX_CORE_WIDTH),
    .SINK_WIDTH(SINK_WIDTH),
    .SOURCE_WIDTH(SOURCE_WIDTH)
  ) u_bridge_wrapper (
    .i_aclk,
    .i_test_mode,
    .i_us_cores_clk(cores_clk),
    .i_us_cores_rst_n(i_cores_rst_n),
    .i_us_cores_dcu_clk(cores_dcu_clk),
    .i_us_cores_l2_clk({CORE_WIDTH{l2c_clk}}),
    .i_us_cores_l2_rst_n({CORE_WIDTH{i_l2c_rst_n}}),
    .i_us_cores_coherent_enable(cores_coherent_enable),
    .o_us_cores_coherent_state(cores_coherent_state),
    .i_us_cores_dcu_a_address(cores_dcu_a_address),
    .i_us_cores_dcu_a_corrupt(cores_dcu_a_corrupt),
    .i_us_cores_dcu_a_data(cores_dcu_a_data),
    .i_us_cores_dcu_a_mask(cores_dcu_a_mask),
    .i_us_cores_dcu_a_opcode(cores_dcu_a_opcode),
    .i_us_cores_dcu_a_param(cores_dcu_a_param),
    .i_us_cores_dcu_a_size(cores_dcu_a_size),
    .i_us_cores_dcu_a_source(cores_dcu_a_source),
    .i_us_cores_dcu_a_user(cores_dcu_a_user),
    .o_us_cores_dcu_a_ready(cores_dcu_a_ready),
    .i_us_cores_dcu_a_valid(cores_dcu_a_valid),
    .o_us_cores_dcu_b_address(cores_dcu_b_address),
    .o_us_cores_dcu_b_corrupt(cores_dcu_b_corrupt),
    .o_us_cores_dcu_b_data(cores_dcu_b_data),
    .o_us_cores_dcu_b_mask(cores_dcu_b_mask),
    .o_us_cores_dcu_b_opcode(cores_dcu_b_opcode),
    .o_us_cores_dcu_b_param(cores_dcu_b_param),
    .o_us_cores_dcu_b_size(cores_dcu_b_size),
    .o_us_cores_dcu_b_source(cores_dcu_b_source),
    .i_us_cores_dcu_b_ready(cores_dcu_b_ready),
    .o_us_cores_dcu_b_valid(cores_dcu_b_valid),
    .i_us_cores_dcu_c_address(cores_dcu_c_address),
    .i_us_cores_dcu_c_corrupt(cores_dcu_c_corrupt),
    .i_us_cores_dcu_c_data(cores_dcu_c_data),
    .i_us_cores_dcu_c_opcode(cores_dcu_c_opcode),
    .i_us_cores_dcu_c_param(cores_dcu_c_param),
    .i_us_cores_dcu_c_size(cores_dcu_c_size),
    .i_us_cores_dcu_c_source(cores_dcu_c_source),
    .i_us_cores_dcu_c_user(cores_dcu_c_user),
    .o_us_cores_dcu_c_ready(cores_dcu_c_ready),
    .i_us_cores_dcu_c_valid(cores_dcu_c_valid),
    .o_us_cores_dcu_d_corrupt(cores_dcu_d_corrupt),
    .o_us_cores_dcu_d_data(cores_dcu_d_data),
    .o_us_cores_dcu_d_denied(cores_dcu_d_denied),
    .o_us_cores_dcu_d_opcode(cores_dcu_d_opcode),
    .o_us_cores_dcu_d_param(cores_dcu_d_param),
    .o_us_cores_dcu_d_size(cores_dcu_d_size),
    .o_us_cores_dcu_d_sink(cores_dcu_d_sink),
    .o_us_cores_dcu_d_source(cores_dcu_d_source),
    .o_us_cores_dcu_d_user(cores_dcu_d_user),
    .i_us_cores_dcu_d_ready(cores_dcu_d_ready),
    .o_us_cores_dcu_d_valid(cores_dcu_d_valid),
    .i_us_cores_dcu_e_sink(cores_dcu_e_sink),
    .o_us_cores_dcu_e_ready(cores_dcu_e_ready),
    .i_us_cores_dcu_e_valid(cores_dcu_e_valid),
    .i_us_cores_icu_a_address(cores_icu_a_address),
    .i_us_cores_icu_a_corrupt(cores_icu_a_corrupt),
    .i_us_cores_icu_a_data(cores_icu_a_data),
    .i_us_cores_icu_a_mask(cores_icu_a_mask),
    .i_us_cores_icu_a_opcode(cores_icu_a_opcode),
    .i_us_cores_icu_a_param(cores_icu_a_param),
    .i_us_cores_icu_a_size(cores_icu_a_size),
    .i_us_cores_icu_a_source(cores_icu_a_source),
    .i_us_cores_icu_a_user(cores_icu_a_user),
    .o_us_cores_icu_a_ready(cores_icu_a_ready),
    .i_us_cores_icu_a_valid(cores_icu_a_valid),
    .o_us_cores_icu_d_corrupt(cores_icu_d_corrupt),
    .o_us_cores_icu_d_data(cores_icu_d_data),
    .o_us_cores_icu_d_denied(cores_icu_d_denied),
    .o_us_cores_icu_d_opcode(cores_icu_d_opcode),
    .o_us_cores_icu_d_param(cores_icu_d_param),
    .o_us_cores_icu_d_size(cores_icu_d_size),
    .o_us_cores_icu_d_sink(cores_icu_d_sink),
    .o_us_cores_icu_d_source(cores_icu_d_source),
    .o_us_cores_icu_d_user(cores_icu_d_user),
    .i_us_cores_icu_d_ready(cores_icu_d_ready),
    .o_us_cores_icu_d_valid(cores_icu_d_valid),
    .i_us_cores_mpipe_axi_s_araddr(cores_mpipe_axi_araddr),
    .i_us_cores_mpipe_axi_s_arburst(cores_mpipe_axi_arburst),
    .i_us_cores_mpipe_axi_s_arcache(cores_mpipe_axi_arcache),
    .i_us_cores_mpipe_axi_s_arid(cores_mpipe_axi_arid),
    .i_us_cores_mpipe_axi_s_arlen(cores_mpipe_axi_arlen),
    .i_us_cores_mpipe_axi_s_arlock(cores_mpipe_axi_arlock),
    .i_us_cores_mpipe_axi_s_arprot(cores_mpipe_axi_arprot),
    .i_us_cores_mpipe_axi_s_arsize(cores_mpipe_axi_arsize),
    .o_us_cores_mpipe_axi_s_arready(cores_mpipe_axi_arready),
    .i_us_cores_mpipe_axi_s_arvalid(cores_mpipe_axi_arvalid),
    .i_us_cores_mpipe_axi_s_awaddr(cores_mpipe_axi_awaddr),
    .i_us_cores_mpipe_axi_s_awburst(cores_mpipe_axi_awburst),
    .i_us_cores_mpipe_axi_s_awcache(cores_mpipe_axi_awcache),
    .i_us_cores_mpipe_axi_s_awid(cores_mpipe_axi_awid),
    .i_us_cores_mpipe_axi_s_awlen(cores_mpipe_axi_awlen),
    .i_us_cores_mpipe_axi_s_awlock(cores_mpipe_axi_awlock),
    .i_us_cores_mpipe_axi_s_awprot(cores_mpipe_axi_awprot),
    .i_us_cores_mpipe_axi_s_awsize(cores_mpipe_axi_awsize),
    .o_us_cores_mpipe_axi_s_awready(cores_mpipe_axi_awready),
    .i_us_cores_mpipe_axi_s_awvalid(cores_mpipe_axi_awvalid),
    .o_us_cores_mpipe_axi_s_bid(cores_mpipe_axi_bid),
    .o_us_cores_mpipe_axi_s_bresp(cores_mpipe_axi_bresp),
    .i_us_cores_mpipe_axi_s_bready(cores_mpipe_axi_bready),
    .o_us_cores_mpipe_axi_s_bvalid(cores_mpipe_axi_bvalid),
    .o_us_cores_mpipe_axi_s_rdata(cores_mpipe_axi_rdata),
    .o_us_cores_mpipe_axi_s_rid(cores_mpipe_axi_rid),
    .o_us_cores_mpipe_axi_s_rlast(cores_mpipe_axi_rlast),
    .o_us_cores_mpipe_axi_s_rresp(cores_mpipe_axi_rresp),
    .i_us_cores_mpipe_axi_s_rready(cores_mpipe_axi_rready),
    .o_us_cores_mpipe_axi_s_rvalid(cores_mpipe_axi_rvalid),
    .i_us_cores_mpipe_axi_s_wdata(cores_mpipe_axi_wdata),
    .i_us_cores_mpipe_axi_s_wlast(cores_mpipe_axi_wlast),
    .i_us_cores_mpipe_axi_s_wstrb(cores_mpipe_axi_wstrb),
    .o_us_cores_mpipe_axi_s_wready(cores_mpipe_axi_wready),
    .i_us_cores_mpipe_axi_s_wvalid(cores_mpipe_axi_wvalid),
    .o_ds_cores_coherent_enable(ds_cores_coherent_enable),
    .i_ds_cores_coherent_state(ds_cores_coherent_state),
    .o_ds_cores_m0_a_address(ds_cores_m0_a_address),
    .o_ds_cores_m0_a_corrupt(ds_cores_m0_a_corrupt),
    .o_ds_cores_m0_a_data(ds_cores_m0_a_data),
    .o_ds_cores_m0_a_mask(ds_cores_m0_a_mask),
    .o_ds_cores_m0_a_opcode(ds_cores_m0_a_opcode),
    .o_ds_cores_m0_a_param(ds_cores_m0_a_param),
    .o_ds_cores_m0_a_size(ds_cores_m0_a_size),
    .o_ds_cores_m0_a_source(ds_cores_m0_a_source),
    .o_ds_cores_m0_a_user(ds_cores_m0_a_user),
    .i_ds_cores_m0_a_ready(ds_cores_m0_a_ready),
    .o_ds_cores_m0_a_valid(ds_cores_m0_a_valid),
    .i_ds_cores_m0_b_address(ds_cores_m0_b_address),
    .i_ds_cores_m0_b_corrupt(ds_cores_m0_b_corrupt),
    .i_ds_cores_m0_b_data(ds_cores_m0_b_data),
    .i_ds_cores_m0_b_mask(ds_cores_m0_b_mask),
    .i_ds_cores_m0_b_opcode(ds_cores_m0_b_opcode),
    .i_ds_cores_m0_b_param(ds_cores_m0_b_param),
    .i_ds_cores_m0_b_size(ds_cores_m0_b_size),
    .i_ds_cores_m0_b_source(ds_cores_m0_b_source),
    .o_ds_cores_m0_b_ready(ds_cores_m0_b_ready),
    .i_ds_cores_m0_b_valid(ds_cores_m0_b_valid),
    .o_ds_cores_m0_c_address(ds_cores_m0_c_address),
    .o_ds_cores_m0_c_corrupt(ds_cores_m0_c_corrupt),
    .o_ds_cores_m0_c_data(ds_cores_m0_c_data),
    .o_ds_cores_m0_c_opcode(ds_cores_m0_c_opcode),
    .o_ds_cores_m0_c_param(ds_cores_m0_c_param),
    .o_ds_cores_m0_c_size(ds_cores_m0_c_size),
    .o_ds_cores_m0_c_source(ds_cores_m0_c_source),
    .o_ds_cores_m0_c_user(ds_cores_m0_c_user),
    .i_ds_cores_m0_c_ready(ds_cores_m0_c_ready),
    .o_ds_cores_m0_c_valid(ds_cores_m0_c_valid),
    .i_ds_cores_m0_d_corrupt(ds_cores_m0_d_corrupt),
    .i_ds_cores_m0_d_data(ds_cores_m0_d_data),
    .i_ds_cores_m0_d_denied(ds_cores_m0_d_denied),
    .i_ds_cores_m0_d_opcode(ds_cores_m0_d_opcode),
    .i_ds_cores_m0_d_param(ds_cores_m0_d_param),
    .i_ds_cores_m0_d_size(ds_cores_m0_d_size),
    .i_ds_cores_m0_d_sink(ds_cores_m0_d_sink),
    .i_ds_cores_m0_d_source(ds_cores_m0_d_source),
    .i_ds_cores_m0_d_user(ds_cores_m0_d_user),
    .o_ds_cores_m0_d_ready(ds_cores_m0_d_ready),
    .i_ds_cores_m0_d_valid(ds_cores_m0_d_valid),
    .o_ds_cores_m0_e_sink(ds_cores_m0_e_sink),
    .i_ds_cores_m0_e_ready(ds_cores_m0_e_ready),
    .o_ds_cores_m0_e_valid(ds_cores_m0_e_valid),
    .o_ds_cores_m1_axi_m_araddr(ds_cores_m1_axi_araddr),
    .o_ds_cores_m1_axi_m_arburst(ds_cores_m1_axi_arburst),
    .o_ds_cores_m1_axi_m_arcache(ds_cores_m1_axi_arcache),
    .o_ds_cores_m1_axi_m_arid(ds_cores_m1_axi_arid),
    .o_ds_cores_m1_axi_m_arlen(ds_cores_m1_axi_arlen),
    .o_ds_cores_m1_axi_m_arlock(ds_cores_m1_axi_arlock),
    .o_ds_cores_m1_axi_m_arprot(ds_cores_m1_axi_arprot),
    .o_ds_cores_m1_axi_m_arsize(ds_cores_m1_axi_arsize),
    .i_ds_cores_m1_axi_m_arready(ds_cores_m1_axi_arready),
    .o_ds_cores_m1_axi_m_arvalid(ds_cores_m1_axi_arvalid),
    .o_ds_cores_m1_axi_m_awaddr(ds_cores_m1_axi_awaddr),
    .o_ds_cores_m1_axi_m_awburst(ds_cores_m1_axi_awburst),
    .o_ds_cores_m1_axi_m_awcache(ds_cores_m1_axi_awcache),
    .o_ds_cores_m1_axi_m_awid(ds_cores_m1_axi_awid),
    .o_ds_cores_m1_axi_m_awlen(ds_cores_m1_axi_awlen),
    .o_ds_cores_m1_axi_m_awlock(ds_cores_m1_axi_awlock),
    .o_ds_cores_m1_axi_m_awprot(ds_cores_m1_axi_awprot),
    .o_ds_cores_m1_axi_m_awsize(ds_cores_m1_axi_awsize),
    .i_ds_cores_m1_axi_m_awready(ds_cores_m1_axi_awready),
    .o_ds_cores_m1_axi_m_awvalid(ds_cores_m1_axi_awvalid),
    .i_ds_cores_m1_axi_m_bid(ds_cores_m1_axi_bid),
    .i_ds_cores_m1_axi_m_bresp(ds_cores_m1_axi_bresp),
    .o_ds_cores_m1_axi_m_bready(ds_cores_m1_axi_bready),
    .o_ds_cores_m1_axi_m_bvalid(ds_cores_m1_axi_bvalid),
    .i_ds_cores_m1_axi_m_rdata(ds_cores_m1_axi_rdata),
    .i_ds_cores_m1_axi_m_rid(ds_cores_m1_axi_rid),
    .i_ds_cores_m1_axi_m_rlast(ds_cores_m1_axi_rlast),
    .i_ds_cores_m1_axi_m_rresp(ds_cores_m1_axi_rresp),
    .o_ds_cores_m1_axi_m_rready(ds_cores_m1_axi_rready),
    .o_ds_cores_m1_axi_m_rvalid(ds_cores_m1_axi_rvalid),
    .o_ds_cores_m1_axi_m_wdata(ds_cores_m1_axi_wdata),
    .o_ds_cores_m1_axi_m_wlast(ds_cores_m1_axi_wlast),
    .o_ds_cores_m1_axi_m_wstrb(ds_cores_m1_axi_wstrb),
    .i_ds_cores_m1_axi_m_wready(ds_cores_m1_axi_wready),
    .o_ds_cores_m1_axi_m_wvalid(ds_cores_m1_axi_wvalid),
    .o_ds_cores_m2_a_address(ds_cores_m2_a_address),
    .o_ds_cores_m2_a_corrupt(ds_cores_m2_a_corrupt),
    .o_ds_cores_m2_a_data(ds_cores_m2_a_data),
    .o_ds_cores_m2_a_mask(ds_cores_m2_a_mask),
    .o_ds_cores_m2_a_opcode(ds_cores_m2_a_opcode),
    .o_ds_cores_m2_a_param(ds_cores_m2_a_param),
    .o_ds_cores_m2_a_size(ds_cores_m2_a_size),
    .o_ds_cores_m2_a_source(ds_cores_m2_a_source),
    .o_ds_cores_m2_a_user(ds_cores_m2_a_user),
    .i_ds_cores_m2_a_ready(ds_cores_m2_a_ready),
    .o_ds_cores_m2_a_valid(ds_cores_m2_a_valid),
    .i_ds_cores_m2_d_corrupt(ds_cores_m2_d_corrupt),
    .i_ds_cores_m2_d_data(ds_cores_m2_d_data),
    .i_ds_cores_m2_d_denied(ds_cores_m2_d_denied),
    .i_ds_cores_m2_d_opcode(ds_cores_m2_d_opcode),
    .i_ds_cores_m2_d_param(ds_cores_m2_d_param),
    .i_ds_cores_m2_d_size(ds_cores_m2_d_size),
    .i_ds_cores_m2_d_sink(ds_cores_m2_d_sink),
    .i_ds_cores_m2_d_source(ds_cores_m2_d_source),
    .i_ds_cores_m2_d_user(ds_cores_m2_d_user),
    .o_ds_cores_m2_d_ready(ds_cores_m2_d_ready),
    .i_ds_cores_m2_d_valid(ds_cores_m2_d_valid)
  );

  apu_l2c_p u_l2c_p (
    .i_clk(l2c_clk),
    .i_rst_n(i_l2c_rst_n),
    .i_aclk,
    .i_arst_n,
    .i_l2c_banks_clk(l2c_banks_clk),
    .i_l2c_banks_clk_en(l2c_banks_clk_en),

    // JTAG
    .ijtag_tck('0),
    .ijtag_reset('0),
    .ijtag_sel('0),
    .ijtag_ue('0),
    .ijtag_se('0),
    .ijtag_ce('0),
    .ijtag_si('0),
    .ijtag_so(),
    // DFT
    .test_clk('0),
    .test_mode('0),
    .edt_update('0),
    .scan_en('0),
    .scan_in('0),
    .scan_out(),
    // BIST
    .bisr_clk('0),
    .bisr_reset('0),
    .bisr_shift_en('0),
    .bisr_si('0),
    .bisr_so(),

    //////////////////////////////////////////////
    /// CORES sigs
    //////////////////////////////////////////////
    .i_core0_coherent_enable(ds_cores_coherent_enable[0]),
    .o_core0_coherent_state(ds_cores_coherent_state[0]),
    .i_core0_m0_a_address(ds_cores_m0_a_address[0]),
    .i_core0_m0_a_corrupt(ds_cores_m0_a_corrupt[0]),
    .i_core0_m0_a_data(ds_cores_m0_a_data[0]),
    .i_core0_m0_a_mask(ds_cores_m0_a_mask[0]),
    .i_core0_m0_a_opcode(ds_cores_m0_a_opcode[0]),
    .i_core0_m0_a_param(ds_cores_m0_a_param[0]),
    .i_core0_m0_a_size(ds_cores_m0_a_size[0]),
    .i_core0_m0_a_source(ds_cores_m0_a_source[0]),
    .i_core0_m0_a_user(ds_cores_m0_a_user[0]),
    .o_core0_m0_a_ready(ds_cores_m0_a_ready[0]),
    .i_core0_m0_a_valid(ds_cores_m0_a_valid[0]),
    .o_core0_m0_b_address(ds_cores_m0_b_address[0]),
    .o_core0_m0_b_corrupt(ds_cores_m0_b_corrupt[0]),
    .o_core0_m0_b_data(ds_cores_m0_b_data[0]),
    .o_core0_m0_b_mask(ds_cores_m0_b_mask[0]),
    .o_core0_m0_b_opcode(ds_cores_m0_b_opcode[0]),
    .o_core0_m0_b_param(ds_cores_m0_b_param[0]),
    .o_core0_m0_b_size(ds_cores_m0_b_size[0]),
    .o_core0_m0_b_source(ds_cores_m0_b_source[0]),
    .i_core0_m0_b_ready(ds_cores_m0_b_ready[0]),
    .o_core0_m0_b_valid(ds_cores_m0_b_valid[0]),
    .i_core0_m0_c_address(ds_cores_m0_c_address[0]),
    .i_core0_m0_c_corrupt(ds_cores_m0_c_corrupt[0]),
    .i_core0_m0_c_data(ds_cores_m0_c_data[0]),
    .i_core0_m0_c_opcode(ds_cores_m0_c_opcode[0]),
    .i_core0_m0_c_param(ds_cores_m0_c_param[0]),
    .i_core0_m0_c_size(ds_cores_m0_c_size[0]),
    .i_core0_m0_c_source(ds_cores_m0_c_source[0]),
    .i_core0_m0_c_user(ds_cores_m0_c_user[0]),
    .o_core0_m0_c_ready(ds_cores_m0_c_ready[0]),
    .i_core0_m0_c_valid(ds_cores_m0_c_valid[0]),
    .o_core0_m0_d_corrupt(ds_cores_m0_d_corrupt[0]),
    .o_core0_m0_d_data(ds_cores_m0_d_data[0]),
    .o_core0_m0_d_denied(ds_cores_m0_d_denied[0]),
    .o_core0_m0_d_opcode(ds_cores_m0_d_opcode[0]),
    .o_core0_m0_d_param(ds_cores_m0_d_param[0]),
    .o_core0_m0_d_size(ds_cores_m0_d_size[0]),
    .o_core0_m0_d_sink(ds_cores_m0_d_sink[0]),
    .o_core0_m0_d_source(ds_cores_m0_d_source[0]),
    .o_core0_m0_d_user(ds_cores_m0_d_user[0]),
    .i_core0_m0_d_ready(ds_cores_m0_d_ready[0]),
    .o_core0_m0_d_valid(ds_cores_m0_d_valid[0]),
    .i_core0_m0_e_sink(ds_cores_m0_e_sink[0]),
    .o_core0_m0_e_ready(ds_cores_m0_e_ready[0]),
    .i_core0_m0_e_valid(ds_cores_m0_e_valid[0]),
    .i_core0_m1_axi_s_araddr(ds_cores_m1_axi_araddr[0]),
    .i_core0_m1_axi_s_arburst(ds_cores_m1_axi_arburst[0]),
    .i_core0_m1_axi_s_arcache(ds_cores_m1_axi_arcache[0]),
    .i_core0_m1_axi_s_arid(ds_cores_m1_axi_arid[0]),
    .i_core0_m1_axi_s_arlen(ds_cores_m1_axi_arlen[0]),
    .i_core0_m1_axi_s_arlock(ds_cores_m1_axi_arlock[0]),
    .i_core0_m1_axi_s_arprot(ds_cores_m1_axi_arprot[0]),
    .i_core0_m1_axi_s_arsize(ds_cores_m1_axi_arsize[0]),
    .o_core0_m1_axi_s_arready(ds_cores_m1_axi_arready[0]),
    .i_core0_m1_axi_s_arvalid(ds_cores_m1_axi_arvalid[0]),
    .i_core0_m1_axi_s_awaddr(ds_cores_m1_axi_awaddr[0]),
    .i_core0_m1_axi_s_awburst(ds_cores_m1_axi_awburst[0]),
    .i_core0_m1_axi_s_awcache(ds_cores_m1_axi_awcache[0]),
    .i_core0_m1_axi_s_awid(ds_cores_m1_axi_awid[0]),
    .i_core0_m1_axi_s_awlen(ds_cores_m1_axi_awlen[0]),
    .i_core0_m1_axi_s_awlock(ds_cores_m1_axi_awlock[0]),
    .i_core0_m1_axi_s_awprot(ds_cores_m1_axi_awprot[0]),
    .i_core0_m1_axi_s_awsize(ds_cores_m1_axi_awsize[0]),
    .o_core0_m1_axi_s_awready(ds_cores_m1_axi_awready[0]),
    .i_core0_m1_axi_s_awvalid(ds_cores_m1_axi_awvalid[0]),
    .o_core0_m1_axi_s_bid(ds_cores_m1_axi_bid[0]),
    .o_core0_m1_axi_s_bresp(ds_cores_m1_axi_bresp[0]),
    .i_core0_m1_axi_s_bready(ds_cores_m1_axi_bready[0]),
    .o_core0_m1_axi_s_bvalid(ds_cores_m1_axi_bvalid[0]),
    .o_core0_m1_axi_s_rdata(ds_cores_m1_axi_rdata[0]),
    .o_core0_m1_axi_s_rid(ds_cores_m1_axi_rid[0]),
    .o_core0_m1_axi_s_rlast(ds_cores_m1_axi_rlast[0]),
    .o_core0_m1_axi_s_rresp(ds_cores_m1_axi_rresp[0]),
    .i_core0_m1_axi_s_rready(ds_cores_m1_axi_rready[0]),
    .o_core0_m1_axi_s_rvalid(ds_cores_m1_axi_rvalid[0]),
    .i_core0_m1_axi_s_wdata(ds_cores_m1_axi_wdata[0]),
    .i_core0_m1_axi_s_wlast(ds_cores_m1_axi_wlast[0]),
    .i_core0_m1_axi_s_wstrb(ds_cores_m1_axi_wstrb[0]),
    .o_core0_m1_axi_s_wready(ds_cores_m1_axi_wready[0]),
    .i_core0_m1_axi_s_wvalid(ds_cores_m1_axi_wvalid[0]),
    .i_core0_m2_a_address(ds_cores_m2_a_address[0]),
    .i_core0_m2_a_corrupt(ds_cores_m2_a_corrupt[0]),
    .i_core0_m2_a_data(ds_cores_m2_a_data[0]),
    .i_core0_m2_a_mask(ds_cores_m2_a_mask[0]),
    .i_core0_m2_a_opcode(ds_cores_m2_a_opcode[0]),
    .i_core0_m2_a_param(ds_cores_m2_a_param[0]),
    .i_core0_m2_a_size(ds_cores_m2_a_size[0]),
    .i_core0_m2_a_source(ds_cores_m2_a_source[0]),
    .i_core0_m2_a_user(ds_cores_m2_a_user[0]),
    .o_core0_m2_a_ready(ds_cores_m2_a_ready[0]),
    .i_core0_m2_a_valid(ds_cores_m2_a_valid[0]),
    .o_core0_m2_d_corrupt(ds_cores_m2_d_corrupt[0]),
    .o_core0_m2_d_data(ds_cores_m2_d_data[0]),
    .o_core0_m2_d_denied(ds_cores_m2_d_denied[0]),
    .o_core0_m2_d_opcode(ds_cores_m2_d_opcode[0]),
    .o_core0_m2_d_param(ds_cores_m2_d_param[0]),
    .o_core0_m2_d_size(ds_cores_m2_d_size[0]),
    .o_core0_m2_d_sink(ds_cores_m2_d_sink[0]),
    .o_core0_m2_d_source(ds_cores_m2_d_source[0]),
    .o_core0_m2_d_user(ds_cores_m2_d_user[0]),
    .i_core0_m2_d_ready(ds_cores_m2_d_ready[0]),
    .o_core0_m2_d_valid(ds_cores_m2_d_valid[0]),

    .i_core1_coherent_enable(ds_cores_coherent_enable[1]),
    .o_core1_coherent_state(ds_cores_coherent_state[1]),
    .i_core1_m0_a_address(ds_cores_m0_a_address[1]),
    .i_core1_m0_a_corrupt(ds_cores_m0_a_corrupt[1]),
    .i_core1_m0_a_data(ds_cores_m0_a_data[1]),
    .i_core1_m0_a_mask(ds_cores_m0_a_mask[1]),
    .i_core1_m0_a_opcode(ds_cores_m0_a_opcode[1]),
    .i_core1_m0_a_param(ds_cores_m0_a_param[1]),
    .i_core1_m0_a_size(ds_cores_m0_a_size[1]),
    .i_core1_m0_a_source(ds_cores_m0_a_source[1]),
    .i_core1_m0_a_user(ds_cores_m0_a_user[1]),
    .o_core1_m0_a_ready(ds_cores_m0_a_ready[1]),
    .i_core1_m0_a_valid(ds_cores_m0_a_valid[1]),
    .o_core1_m0_b_address(ds_cores_m0_b_address[1]),
    .o_core1_m0_b_corrupt(ds_cores_m0_b_corrupt[1]),
    .o_core1_m0_b_data(ds_cores_m0_b_data[1]),
    .o_core1_m0_b_mask(ds_cores_m0_b_mask[1]),
    .o_core1_m0_b_opcode(ds_cores_m0_b_opcode[1]),
    .o_core1_m0_b_param(ds_cores_m0_b_param[1]),
    .o_core1_m0_b_size(ds_cores_m0_b_size[1]),
    .o_core1_m0_b_source(ds_cores_m0_b_source[1]),
    .i_core1_m0_b_ready(ds_cores_m0_b_ready[1]),
    .o_core1_m0_b_valid(ds_cores_m0_b_valid[1]),
    .i_core1_m0_c_address(ds_cores_m0_c_address[1]),
    .i_core1_m0_c_corrupt(ds_cores_m0_c_corrupt[1]),
    .i_core1_m0_c_data(ds_cores_m0_c_data[1]),
    .i_core1_m0_c_opcode(ds_cores_m0_c_opcode[1]),
    .i_core1_m0_c_param(ds_cores_m0_c_param[1]),
    .i_core1_m0_c_size(ds_cores_m0_c_size[1]),
    .i_core1_m0_c_source(ds_cores_m0_c_source[1]),
    .i_core1_m0_c_user(ds_cores_m0_c_user[1]),
    .o_core1_m0_c_ready(ds_cores_m0_c_ready[1]),
    .i_core1_m0_c_valid(ds_cores_m0_c_valid[1]),
    .o_core1_m0_d_corrupt(ds_cores_m0_d_corrupt[1]),
    .o_core1_m0_d_data(ds_cores_m0_d_data[1]),
    .o_core1_m0_d_denied(ds_cores_m0_d_denied[1]),
    .o_core1_m0_d_opcode(ds_cores_m0_d_opcode[1]),
    .o_core1_m0_d_param(ds_cores_m0_d_param[1]),
    .o_core1_m0_d_size(ds_cores_m0_d_size[1]),
    .o_core1_m0_d_sink(ds_cores_m0_d_sink[1]),
    .o_core1_m0_d_source(ds_cores_m0_d_source[1]),
    .o_core1_m0_d_user(ds_cores_m0_d_user[1]),
    .i_core1_m0_d_ready(ds_cores_m0_d_ready[1]),
    .o_core1_m0_d_valid(ds_cores_m0_d_valid[1]),
    .i_core1_m0_e_sink(ds_cores_m0_e_sink[1]),
    .o_core1_m0_e_ready(ds_cores_m0_e_ready[1]),
    .i_core1_m0_e_valid(ds_cores_m0_e_valid[1]),
    .i_core1_m1_axi_s_araddr(ds_cores_m1_axi_araddr[1]),
    .i_core1_m1_axi_s_arburst(ds_cores_m1_axi_arburst[1]),
    .i_core1_m1_axi_s_arcache(ds_cores_m1_axi_arcache[1]),
    .i_core1_m1_axi_s_arid(ds_cores_m1_axi_arid[1]),
    .i_core1_m1_axi_s_arlen(ds_cores_m1_axi_arlen[1]),
    .i_core1_m1_axi_s_arlock(ds_cores_m1_axi_arlock[1]),
    .i_core1_m1_axi_s_arprot(ds_cores_m1_axi_arprot[1]),
    .i_core1_m1_axi_s_arsize(ds_cores_m1_axi_arsize[1]),
    .o_core1_m1_axi_s_arready(ds_cores_m1_axi_arready[1]),
    .i_core1_m1_axi_s_arvalid(ds_cores_m1_axi_arvalid[1]),
    .i_core1_m1_axi_s_awaddr(ds_cores_m1_axi_awaddr[1]),
    .i_core1_m1_axi_s_awburst(ds_cores_m1_axi_awburst[1]),
    .i_core1_m1_axi_s_awcache(ds_cores_m1_axi_awcache[1]),
    .i_core1_m1_axi_s_awid(ds_cores_m1_axi_awid[1]),
    .i_core1_m1_axi_s_awlen(ds_cores_m1_axi_awlen[1]),
    .i_core1_m1_axi_s_awlock(ds_cores_m1_axi_awlock[1]),
    .i_core1_m1_axi_s_awprot(ds_cores_m1_axi_awprot[1]),
    .i_core1_m1_axi_s_awsize(ds_cores_m1_axi_awsize[1]),
    .o_core1_m1_axi_s_awready(ds_cores_m1_axi_awready[1]),
    .i_core1_m1_axi_s_awvalid(ds_cores_m1_axi_awvalid[1]),
    .o_core1_m1_axi_s_bid(ds_cores_m1_axi_bid[1]),
    .o_core1_m1_axi_s_bresp(ds_cores_m1_axi_bresp[1]),
    .i_core1_m1_axi_s_bready(ds_cores_m1_axi_bready[1]),
    .o_core1_m1_axi_s_bvalid(ds_cores_m1_axi_bvalid[1]),
    .o_core1_m1_axi_s_rdata(ds_cores_m1_axi_rdata[1]),
    .o_core1_m1_axi_s_rid(ds_cores_m1_axi_rid[1]),
    .o_core1_m1_axi_s_rlast(ds_cores_m1_axi_rlast[1]),
    .o_core1_m1_axi_s_rresp(ds_cores_m1_axi_rresp[1]),
    .i_core1_m1_axi_s_rready(ds_cores_m1_axi_rready[1]),
    .o_core1_m1_axi_s_rvalid(ds_cores_m1_axi_rvalid[1]),
    .i_core1_m1_axi_s_wdata(ds_cores_m1_axi_wdata[1]),
    .i_core1_m1_axi_s_wlast(ds_cores_m1_axi_wlast[1]),
    .i_core1_m1_axi_s_wstrb(ds_cores_m1_axi_wstrb[1]),
    .o_core1_m1_axi_s_wready(ds_cores_m1_axi_wready[1]),
    .i_core1_m1_axi_s_wvalid(ds_cores_m1_axi_wvalid[1]),
    .i_core1_m2_a_address(ds_cores_m2_a_address[1]),
    .i_core1_m2_a_corrupt(ds_cores_m2_a_corrupt[1]),
    .i_core1_m2_a_data(ds_cores_m2_a_data[1]),
    .i_core1_m2_a_mask(ds_cores_m2_a_mask[1]),
    .i_core1_m2_a_opcode(ds_cores_m2_a_opcode[1]),
    .i_core1_m2_a_param(ds_cores_m2_a_param[1]),
    .i_core1_m2_a_size(ds_cores_m2_a_size[1]),
    .i_core1_m2_a_source(ds_cores_m2_a_source[1]),
    .i_core1_m2_a_user(ds_cores_m2_a_user[1]),
    .o_core1_m2_a_ready(ds_cores_m2_a_ready[1]),
    .i_core1_m2_a_valid(ds_cores_m2_a_valid[1]),
    .o_core1_m2_d_corrupt(ds_cores_m2_d_corrupt[1]),
    .o_core1_m2_d_data(ds_cores_m2_d_data[1]),
    .o_core1_m2_d_denied(ds_cores_m2_d_denied[1]),
    .o_core1_m2_d_opcode(ds_cores_m2_d_opcode[1]),
    .o_core1_m2_d_param(ds_cores_m2_d_param[1]),
    .o_core1_m2_d_size(ds_cores_m2_d_size[1]),
    .o_core1_m2_d_sink(ds_cores_m2_d_sink[1]),
    .o_core1_m2_d_source(ds_cores_m2_d_source[1]),
    .o_core1_m2_d_user(ds_cores_m2_d_user[1]),
    .i_core1_m2_d_ready(ds_cores_m2_d_ready[1]),
    .o_core1_m2_d_valid(ds_cores_m2_d_valid[1]),

    .i_core2_coherent_enable(ds_cores_coherent_enable[2]),
    .o_core2_coherent_state(ds_cores_coherent_state[2]),
    .i_core2_m0_a_address(ds_cores_m0_a_address[2]),
    .i_core2_m0_a_corrupt(ds_cores_m0_a_corrupt[2]),
    .i_core2_m0_a_data(ds_cores_m0_a_data[2]),
    .i_core2_m0_a_mask(ds_cores_m0_a_mask[2]),
    .i_core2_m0_a_opcode(ds_cores_m0_a_opcode[2]),
    .i_core2_m0_a_param(ds_cores_m0_a_param[2]),
    .i_core2_m0_a_size(ds_cores_m0_a_size[2]),
    .i_core2_m0_a_source(ds_cores_m0_a_source[2]),
    .i_core2_m0_a_user(ds_cores_m0_a_user[2]),
    .o_core2_m0_a_ready(ds_cores_m0_a_ready[2]),
    .i_core2_m0_a_valid(ds_cores_m0_a_valid[2]),
    .o_core2_m0_b_address(ds_cores_m0_b_address[2]),
    .o_core2_m0_b_corrupt(ds_cores_m0_b_corrupt[2]),
    .o_core2_m0_b_data(ds_cores_m0_b_data[2]),
    .o_core2_m0_b_mask(ds_cores_m0_b_mask[2]),
    .o_core2_m0_b_opcode(ds_cores_m0_b_opcode[2]),
    .o_core2_m0_b_param(ds_cores_m0_b_param[2]),
    .o_core2_m0_b_size(ds_cores_m0_b_size[2]),
    .o_core2_m0_b_source(ds_cores_m0_b_source[2]),
    .i_core2_m0_b_ready(ds_cores_m0_b_ready[2]),
    .o_core2_m0_b_valid(ds_cores_m0_b_valid[2]),
    .i_core2_m0_c_address(ds_cores_m0_c_address[2]),
    .i_core2_m0_c_corrupt(ds_cores_m0_c_corrupt[2]),
    .i_core2_m0_c_data(ds_cores_m0_c_data[2]),
    .i_core2_m0_c_opcode(ds_cores_m0_c_opcode[2]),
    .i_core2_m0_c_param(ds_cores_m0_c_param[2]),
    .i_core2_m0_c_size(ds_cores_m0_c_size[2]),
    .i_core2_m0_c_source(ds_cores_m0_c_source[2]),
    .i_core2_m0_c_user(ds_cores_m0_c_user[2]),
    .o_core2_m0_c_ready(ds_cores_m0_c_ready[2]),
    .i_core2_m0_c_valid(ds_cores_m0_c_valid[2]),
    .o_core2_m0_d_corrupt(ds_cores_m0_d_corrupt[2]),
    .o_core2_m0_d_data(ds_cores_m0_d_data[2]),
    .o_core2_m0_d_denied(ds_cores_m0_d_denied[2]),
    .o_core2_m0_d_opcode(ds_cores_m0_d_opcode[2]),
    .o_core2_m0_d_param(ds_cores_m0_d_param[2]),
    .o_core2_m0_d_size(ds_cores_m0_d_size[2]),
    .o_core2_m0_d_sink(ds_cores_m0_d_sink[2]),
    .o_core2_m0_d_source(ds_cores_m0_d_source[2]),
    .o_core2_m0_d_user(ds_cores_m0_d_user[2]),
    .i_core2_m0_d_ready(ds_cores_m0_d_ready[2]),
    .o_core2_m0_d_valid(ds_cores_m0_d_valid[2]),
    .i_core2_m0_e_sink(ds_cores_m0_e_sink[2]),
    .o_core2_m0_e_ready(ds_cores_m0_e_ready[2]),
    .i_core2_m0_e_valid(ds_cores_m0_e_valid[2]),
    .i_core2_m1_axi_s_araddr(ds_cores_m1_axi_araddr[2]),
    .i_core2_m1_axi_s_arburst(ds_cores_m1_axi_arburst[2]),
    .i_core2_m1_axi_s_arcache(ds_cores_m1_axi_arcache[2]),
    .i_core2_m1_axi_s_arid(ds_cores_m1_axi_arid[2]),
    .i_core2_m1_axi_s_arlen(ds_cores_m1_axi_arlen[2]),
    .i_core2_m1_axi_s_arlock(ds_cores_m1_axi_arlock[2]),
    .i_core2_m1_axi_s_arprot(ds_cores_m1_axi_arprot[2]),
    .i_core2_m1_axi_s_arsize(ds_cores_m1_axi_arsize[2]),
    .o_core2_m1_axi_s_arready(ds_cores_m1_axi_arready[2]),
    .i_core2_m1_axi_s_arvalid(ds_cores_m1_axi_arvalid[2]),
    .i_core2_m1_axi_s_awaddr(ds_cores_m1_axi_awaddr[2]),
    .i_core2_m1_axi_s_awburst(ds_cores_m1_axi_awburst[2]),
    .i_core2_m1_axi_s_awcache(ds_cores_m1_axi_awcache[2]),
    .i_core2_m1_axi_s_awid(ds_cores_m1_axi_awid[2]),
    .i_core2_m1_axi_s_awlen(ds_cores_m1_axi_awlen[2]),
    .i_core2_m1_axi_s_awlock(ds_cores_m1_axi_awlock[2]),
    .i_core2_m1_axi_s_awprot(ds_cores_m1_axi_awprot[2]),
    .i_core2_m1_axi_s_awsize(ds_cores_m1_axi_awsize[2]),
    .o_core2_m1_axi_s_awready(ds_cores_m1_axi_awready[2]),
    .i_core2_m1_axi_s_awvalid(ds_cores_m1_axi_awvalid[2]),
    .o_core2_m1_axi_s_bid(ds_cores_m1_axi_bid[2]),
    .o_core2_m1_axi_s_bresp(ds_cores_m1_axi_bresp[2]),
    .i_core2_m1_axi_s_bready(ds_cores_m1_axi_bready[2]),
    .o_core2_m1_axi_s_bvalid(ds_cores_m1_axi_bvalid[2]),
    .o_core2_m1_axi_s_rdata(ds_cores_m1_axi_rdata[2]),
    .o_core2_m1_axi_s_rid(ds_cores_m1_axi_rid[2]),
    .o_core2_m1_axi_s_rlast(ds_cores_m1_axi_rlast[2]),
    .o_core2_m1_axi_s_rresp(ds_cores_m1_axi_rresp[2]),
    .i_core2_m1_axi_s_rready(ds_cores_m1_axi_rready[2]),
    .o_core2_m1_axi_s_rvalid(ds_cores_m1_axi_rvalid[2]),
    .i_core2_m1_axi_s_wdata(ds_cores_m1_axi_wdata[2]),
    .i_core2_m1_axi_s_wlast(ds_cores_m1_axi_wlast[2]),
    .i_core2_m1_axi_s_wstrb(ds_cores_m1_axi_wstrb[2]),
    .o_core2_m1_axi_s_wready(ds_cores_m1_axi_wready[2]),
    .i_core2_m1_axi_s_wvalid(ds_cores_m1_axi_wvalid[2]),
    .i_core2_m2_a_address(ds_cores_m2_a_address[2]),
    .i_core2_m2_a_corrupt(ds_cores_m2_a_corrupt[2]),
    .i_core2_m2_a_data(ds_cores_m2_a_data[2]),
    .i_core2_m2_a_mask(ds_cores_m2_a_mask[2]),
    .i_core2_m2_a_opcode(ds_cores_m2_a_opcode[2]),
    .i_core2_m2_a_param(ds_cores_m2_a_param[2]),
    .i_core2_m2_a_size(ds_cores_m2_a_size[2]),
    .i_core2_m2_a_source(ds_cores_m2_a_source[2]),
    .i_core2_m2_a_user(ds_cores_m2_a_user[2]),
    .o_core2_m2_a_ready(ds_cores_m2_a_ready[2]),
    .i_core2_m2_a_valid(ds_cores_m2_a_valid[2]),
    .o_core2_m2_d_corrupt(ds_cores_m2_d_corrupt[2]),
    .o_core2_m2_d_data(ds_cores_m2_d_data[2]),
    .o_core2_m2_d_denied(ds_cores_m2_d_denied[2]),
    .o_core2_m2_d_opcode(ds_cores_m2_d_opcode[2]),
    .o_core2_m2_d_param(ds_cores_m2_d_param[2]),
    .o_core2_m2_d_size(ds_cores_m2_d_size[2]),
    .o_core2_m2_d_sink(ds_cores_m2_d_sink[2]),
    .o_core2_m2_d_source(ds_cores_m2_d_source[2]),
    .o_core2_m2_d_user(ds_cores_m2_d_user[2]),
    .i_core2_m2_d_ready(ds_cores_m2_d_ready[2]),
    .o_core2_m2_d_valid(ds_cores_m2_d_valid[2]),

    .i_core3_coherent_enable(ds_cores_coherent_enable[3]),
    .o_core3_coherent_state(ds_cores_coherent_state[3]),
    .i_core3_m0_a_address(ds_cores_m0_a_address[3]),
    .i_core3_m0_a_corrupt(ds_cores_m0_a_corrupt[3]),
    .i_core3_m0_a_data(ds_cores_m0_a_data[3]),
    .i_core3_m0_a_mask(ds_cores_m0_a_mask[3]),
    .i_core3_m0_a_opcode(ds_cores_m0_a_opcode[3]),
    .i_core3_m0_a_param(ds_cores_m0_a_param[3]),
    .i_core3_m0_a_size(ds_cores_m0_a_size[3]),
    .i_core3_m0_a_source(ds_cores_m0_a_source[3]),
    .i_core3_m0_a_user(ds_cores_m0_a_user[3]),
    .o_core3_m0_a_ready(ds_cores_m0_a_ready[3]),
    .i_core3_m0_a_valid(ds_cores_m0_a_valid[3]),
    .o_core3_m0_b_address(ds_cores_m0_b_address[3]),
    .o_core3_m0_b_corrupt(ds_cores_m0_b_corrupt[3]),
    .o_core3_m0_b_data(ds_cores_m0_b_data[3]),
    .o_core3_m0_b_mask(ds_cores_m0_b_mask[3]),
    .o_core3_m0_b_opcode(ds_cores_m0_b_opcode[3]),
    .o_core3_m0_b_param(ds_cores_m0_b_param[3]),
    .o_core3_m0_b_size(ds_cores_m0_b_size[3]),
    .o_core3_m0_b_source(ds_cores_m0_b_source[3]),
    .i_core3_m0_b_ready(ds_cores_m0_b_ready[3]),
    .o_core3_m0_b_valid(ds_cores_m0_b_valid[3]),
    .i_core3_m0_c_address(ds_cores_m0_c_address[3]),
    .i_core3_m0_c_corrupt(ds_cores_m0_c_corrupt[3]),
    .i_core3_m0_c_data(ds_cores_m0_c_data[3]),
    .i_core3_m0_c_opcode(ds_cores_m0_c_opcode[3]),
    .i_core3_m0_c_param(ds_cores_m0_c_param[3]),
    .i_core3_m0_c_size(ds_cores_m0_c_size[3]),
    .i_core3_m0_c_source(ds_cores_m0_c_source[3]),
    .i_core3_m0_c_user(ds_cores_m0_c_user[3]),
    .o_core3_m0_c_ready(ds_cores_m0_c_ready[3]),
    .i_core3_m0_c_valid(ds_cores_m0_c_valid[3]),
    .o_core3_m0_d_corrupt(ds_cores_m0_d_corrupt[3]),
    .o_core3_m0_d_data(ds_cores_m0_d_data[3]),
    .o_core3_m0_d_denied(ds_cores_m0_d_denied[3]),
    .o_core3_m0_d_opcode(ds_cores_m0_d_opcode[3]),
    .o_core3_m0_d_param(ds_cores_m0_d_param[3]),
    .o_core3_m0_d_size(ds_cores_m0_d_size[3]),
    .o_core3_m0_d_sink(ds_cores_m0_d_sink[3]),
    .o_core3_m0_d_source(ds_cores_m0_d_source[3]),
    .o_core3_m0_d_user(ds_cores_m0_d_user[3]),
    .i_core3_m0_d_ready(ds_cores_m0_d_ready[3]),
    .o_core3_m0_d_valid(ds_cores_m0_d_valid[3]),
    .i_core3_m0_e_sink(ds_cores_m0_e_sink[3]),
    .o_core3_m0_e_ready(ds_cores_m0_e_ready[3]),
    .i_core3_m0_e_valid(ds_cores_m0_e_valid[3]),
    .i_core3_m1_axi_s_araddr(ds_cores_m1_axi_araddr[3]),
    .i_core3_m1_axi_s_arburst(ds_cores_m1_axi_arburst[3]),
    .i_core3_m1_axi_s_arcache(ds_cores_m1_axi_arcache[3]),
    .i_core3_m1_axi_s_arid(ds_cores_m1_axi_arid[3]),
    .i_core3_m1_axi_s_arlen(ds_cores_m1_axi_arlen[3]),
    .i_core3_m1_axi_s_arlock(ds_cores_m1_axi_arlock[3]),
    .i_core3_m1_axi_s_arprot(ds_cores_m1_axi_arprot[3]),
    .i_core3_m1_axi_s_arsize(ds_cores_m1_axi_arsize[3]),
    .o_core3_m1_axi_s_arready(ds_cores_m1_axi_arready[3]),
    .i_core3_m1_axi_s_arvalid(ds_cores_m1_axi_arvalid[3]),
    .i_core3_m1_axi_s_awaddr(ds_cores_m1_axi_awaddr[3]),
    .i_core3_m1_axi_s_awburst(ds_cores_m1_axi_awburst[3]),
    .i_core3_m1_axi_s_awcache(ds_cores_m1_axi_awcache[3]),
    .i_core3_m1_axi_s_awid(ds_cores_m1_axi_awid[3]),
    .i_core3_m1_axi_s_awlen(ds_cores_m1_axi_awlen[3]),
    .i_core3_m1_axi_s_awlock(ds_cores_m1_axi_awlock[3]),
    .i_core3_m1_axi_s_awprot(ds_cores_m1_axi_awprot[3]),
    .i_core3_m1_axi_s_awsize(ds_cores_m1_axi_awsize[3]),
    .o_core3_m1_axi_s_awready(ds_cores_m1_axi_awready[3]),
    .i_core3_m1_axi_s_awvalid(ds_cores_m1_axi_awvalid[3]),
    .o_core3_m1_axi_s_bid(ds_cores_m1_axi_bid[3]),
    .o_core3_m1_axi_s_bresp(ds_cores_m1_axi_bresp[3]),
    .i_core3_m1_axi_s_bready(ds_cores_m1_axi_bready[3]),
    .o_core3_m1_axi_s_bvalid(ds_cores_m1_axi_bvalid[3]),
    .o_core3_m1_axi_s_rdata(ds_cores_m1_axi_rdata[3]),
    .o_core3_m1_axi_s_rid(ds_cores_m1_axi_rid[3]),
    .o_core3_m1_axi_s_rlast(ds_cores_m1_axi_rlast[3]),
    .o_core3_m1_axi_s_rresp(ds_cores_m1_axi_rresp[3]),
    .i_core3_m1_axi_s_rready(ds_cores_m1_axi_rready[3]),
    .o_core3_m1_axi_s_rvalid(ds_cores_m1_axi_rvalid[3]),
    .i_core3_m1_axi_s_wdata(ds_cores_m1_axi_wdata[3]),
    .i_core3_m1_axi_s_wlast(ds_cores_m1_axi_wlast[3]),
    .i_core3_m1_axi_s_wstrb(ds_cores_m1_axi_wstrb[3]),
    .o_core3_m1_axi_s_wready(ds_cores_m1_axi_wready[3]),
    .i_core3_m1_axi_s_wvalid(ds_cores_m1_axi_wvalid[3]),
    .i_core3_m2_a_address(ds_cores_m2_a_address[3]),
    .i_core3_m2_a_corrupt(ds_cores_m2_a_corrupt[3]),
    .i_core3_m2_a_data(ds_cores_m2_a_data[3]),
    .i_core3_m2_a_mask(ds_cores_m2_a_mask[3]),
    .i_core3_m2_a_opcode(ds_cores_m2_a_opcode[3]),
    .i_core3_m2_a_param(ds_cores_m2_a_param[3]),
    .i_core3_m2_a_size(ds_cores_m2_a_size[3]),
    .i_core3_m2_a_source(ds_cores_m2_a_source[3]),
    .i_core3_m2_a_user(ds_cores_m2_a_user[3]),
    .o_core3_m2_a_ready(ds_cores_m2_a_ready[3]),
    .i_core3_m2_a_valid(ds_cores_m2_a_valid[3]),
    .o_core3_m2_d_corrupt(ds_cores_m2_d_corrupt[3]),
    .o_core3_m2_d_data(ds_cores_m2_d_data[3]),
    .o_core3_m2_d_denied(ds_cores_m2_d_denied[3]),
    .o_core3_m2_d_opcode(ds_cores_m2_d_opcode[3]),
    .o_core3_m2_d_param(ds_cores_m2_d_param[3]),
    .o_core3_m2_d_size(ds_cores_m2_d_size[3]),
    .o_core3_m2_d_sink(ds_cores_m2_d_sink[3]),
    .o_core3_m2_d_source(ds_cores_m2_d_source[3]),
    .o_core3_m2_d_user(ds_cores_m2_d_user[3]),
    .i_core3_m2_d_ready(ds_cores_m2_d_ready[3]),
    .o_core3_m2_d_valid(ds_cores_m2_d_valid[3]),

    .i_core4_coherent_enable(ds_cores_coherent_enable[4]),
    .o_core4_coherent_state(ds_cores_coherent_state[4]),
    .i_core4_m0_a_address(ds_cores_m0_a_address[4]),
    .i_core4_m0_a_corrupt(ds_cores_m0_a_corrupt[4]),
    .i_core4_m0_a_data(ds_cores_m0_a_data[4]),
    .i_core4_m0_a_mask(ds_cores_m0_a_mask[4]),
    .i_core4_m0_a_opcode(ds_cores_m0_a_opcode[4]),
    .i_core4_m0_a_param(ds_cores_m0_a_param[4]),
    .i_core4_m0_a_size(ds_cores_m0_a_size[4]),
    .i_core4_m0_a_source(ds_cores_m0_a_source[4]),
    .i_core4_m0_a_user(ds_cores_m0_a_user[4]),
    .o_core4_m0_a_ready(ds_cores_m0_a_ready[4]),
    .i_core4_m0_a_valid(ds_cores_m0_a_valid[4]),
    .o_core4_m0_b_address(ds_cores_m0_b_address[4]),
    .o_core4_m0_b_corrupt(ds_cores_m0_b_corrupt[4]),
    .o_core4_m0_b_data(ds_cores_m0_b_data[4]),
    .o_core4_m0_b_mask(ds_cores_m0_b_mask[4]),
    .o_core4_m0_b_opcode(ds_cores_m0_b_opcode[4]),
    .o_core4_m0_b_param(ds_cores_m0_b_param[4]),
    .o_core4_m0_b_size(ds_cores_m0_b_size[4]),
    .o_core4_m0_b_source(ds_cores_m0_b_source[4]),
    .i_core4_m0_b_ready(ds_cores_m0_b_ready[4]),
    .o_core4_m0_b_valid(ds_cores_m0_b_valid[4]),
    .i_core4_m0_c_address(ds_cores_m0_c_address[4]),
    .i_core4_m0_c_corrupt(ds_cores_m0_c_corrupt[4]),
    .i_core4_m0_c_data(ds_cores_m0_c_data[4]),
    .i_core4_m0_c_opcode(ds_cores_m0_c_opcode[4]),
    .i_core4_m0_c_param(ds_cores_m0_c_param[4]),
    .i_core4_m0_c_size(ds_cores_m0_c_size[4]),
    .i_core4_m0_c_source(ds_cores_m0_c_source[4]),
    .i_core4_m0_c_user(ds_cores_m0_c_user[4]),
    .o_core4_m0_c_ready(ds_cores_m0_c_ready[4]),
    .i_core4_m0_c_valid(ds_cores_m0_c_valid[4]),
    .o_core4_m0_d_corrupt(ds_cores_m0_d_corrupt[4]),
    .o_core4_m0_d_data(ds_cores_m0_d_data[4]),
    .o_core4_m0_d_denied(ds_cores_m0_d_denied[4]),
    .o_core4_m0_d_opcode(ds_cores_m0_d_opcode[4]),
    .o_core4_m0_d_param(ds_cores_m0_d_param[4]),
    .o_core4_m0_d_size(ds_cores_m0_d_size[4]),
    .o_core4_m0_d_sink(ds_cores_m0_d_sink[4]),
    .o_core4_m0_d_source(ds_cores_m0_d_source[4]),
    .o_core4_m0_d_user(ds_cores_m0_d_user[4]),
    .i_core4_m0_d_ready(ds_cores_m0_d_ready[4]),
    .o_core4_m0_d_valid(ds_cores_m0_d_valid[4]),
    .i_core4_m0_e_sink(ds_cores_m0_e_sink[4]),
    .o_core4_m0_e_ready(ds_cores_m0_e_ready[4]),
    .i_core4_m0_e_valid(ds_cores_m0_e_valid[4]),
    .i_core4_m1_axi_s_araddr(ds_cores_m1_axi_araddr[4]),
    .i_core4_m1_axi_s_arburst(ds_cores_m1_axi_arburst[4]),
    .i_core4_m1_axi_s_arcache(ds_cores_m1_axi_arcache[4]),
    .i_core4_m1_axi_s_arid(ds_cores_m1_axi_arid[4]),
    .i_core4_m1_axi_s_arlen(ds_cores_m1_axi_arlen[4]),
    .i_core4_m1_axi_s_arlock(ds_cores_m1_axi_arlock[4]),
    .i_core4_m1_axi_s_arprot(ds_cores_m1_axi_arprot[4]),
    .i_core4_m1_axi_s_arsize(ds_cores_m1_axi_arsize[4]),
    .o_core4_m1_axi_s_arready(ds_cores_m1_axi_arready[4]),
    .i_core4_m1_axi_s_arvalid(ds_cores_m1_axi_arvalid[4]),
    .i_core4_m1_axi_s_awaddr(ds_cores_m1_axi_awaddr[4]),
    .i_core4_m1_axi_s_awburst(ds_cores_m1_axi_awburst[4]),
    .i_core4_m1_axi_s_awcache(ds_cores_m1_axi_awcache[4]),
    .i_core4_m1_axi_s_awid(ds_cores_m1_axi_awid[4]),
    .i_core4_m1_axi_s_awlen(ds_cores_m1_axi_awlen[4]),
    .i_core4_m1_axi_s_awlock(ds_cores_m1_axi_awlock[4]),
    .i_core4_m1_axi_s_awprot(ds_cores_m1_axi_awprot[4]),
    .i_core4_m1_axi_s_awsize(ds_cores_m1_axi_awsize[4]),
    .o_core4_m1_axi_s_awready(ds_cores_m1_axi_awready[4]),
    .i_core4_m1_axi_s_awvalid(ds_cores_m1_axi_awvalid[4]),
    .o_core4_m1_axi_s_bid(ds_cores_m1_axi_bid[4]),
    .o_core4_m1_axi_s_bresp(ds_cores_m1_axi_bresp[4]),
    .i_core4_m1_axi_s_bready(ds_cores_m1_axi_bready[4]),
    .o_core4_m1_axi_s_bvalid(ds_cores_m1_axi_bvalid[4]),
    .o_core4_m1_axi_s_rdata(ds_cores_m1_axi_rdata[4]),
    .o_core4_m1_axi_s_rid(ds_cores_m1_axi_rid[4]),
    .o_core4_m1_axi_s_rlast(ds_cores_m1_axi_rlast[4]),
    .o_core4_m1_axi_s_rresp(ds_cores_m1_axi_rresp[4]),
    .i_core4_m1_axi_s_rready(ds_cores_m1_axi_rready[4]),
    .o_core4_m1_axi_s_rvalid(ds_cores_m1_axi_rvalid[4]),
    .i_core4_m1_axi_s_wdata(ds_cores_m1_axi_wdata[4]),
    .i_core4_m1_axi_s_wlast(ds_cores_m1_axi_wlast[4]),
    .i_core4_m1_axi_s_wstrb(ds_cores_m1_axi_wstrb[4]),
    .o_core4_m1_axi_s_wready(ds_cores_m1_axi_wready[4]),
    .i_core4_m1_axi_s_wvalid(ds_cores_m1_axi_wvalid[4]),
    .i_core4_m2_a_address(ds_cores_m2_a_address[4]),
    .i_core4_m2_a_corrupt(ds_cores_m2_a_corrupt[4]),
    .i_core4_m2_a_data(ds_cores_m2_a_data[4]),
    .i_core4_m2_a_mask(ds_cores_m2_a_mask[4]),
    .i_core4_m2_a_opcode(ds_cores_m2_a_opcode[4]),
    .i_core4_m2_a_param(ds_cores_m2_a_param[4]),
    .i_core4_m2_a_size(ds_cores_m2_a_size[4]),
    .i_core4_m2_a_source(ds_cores_m2_a_source[4]),
    .i_core4_m2_a_user(ds_cores_m2_a_user[4]),
    .o_core4_m2_a_ready(ds_cores_m2_a_ready[4]),
    .i_core4_m2_a_valid(ds_cores_m2_a_valid[4]),
    .o_core4_m2_d_corrupt(ds_cores_m2_d_corrupt[4]),
    .o_core4_m2_d_data(ds_cores_m2_d_data[4]),
    .o_core4_m2_d_denied(ds_cores_m2_d_denied[4]),
    .o_core4_m2_d_opcode(ds_cores_m2_d_opcode[4]),
    .o_core4_m2_d_param(ds_cores_m2_d_param[4]),
    .o_core4_m2_d_size(ds_cores_m2_d_size[4]),
    .o_core4_m2_d_sink(ds_cores_m2_d_sink[4]),
    .o_core4_m2_d_source(ds_cores_m2_d_source[4]),
    .o_core4_m2_d_user(ds_cores_m2_d_user[4]),
    .i_core4_m2_d_ready(ds_cores_m2_d_ready[4]),
    .o_core4_m2_d_valid(ds_cores_m2_d_valid[4]),

    .i_core5_coherent_enable(ds_cores_coherent_enable[5]),
    .o_core5_coherent_state(ds_cores_coherent_state[5]),
    .i_core5_m0_a_address(ds_cores_m0_a_address[5]),
    .i_core5_m0_a_corrupt(ds_cores_m0_a_corrupt[5]),
    .i_core5_m0_a_data(ds_cores_m0_a_data[5]),
    .i_core5_m0_a_mask(ds_cores_m0_a_mask[5]),
    .i_core5_m0_a_opcode(ds_cores_m0_a_opcode[5]),
    .i_core5_m0_a_param(ds_cores_m0_a_param[5]),
    .i_core5_m0_a_size(ds_cores_m0_a_size[5]),
    .i_core5_m0_a_source(ds_cores_m0_a_source[5]),
    .i_core5_m0_a_user(ds_cores_m0_a_user[5]),
    .o_core5_m0_a_ready(ds_cores_m0_a_ready[5]),
    .i_core5_m0_a_valid(ds_cores_m0_a_valid[5]),
    .o_core5_m0_b_address(ds_cores_m0_b_address[5]),
    .o_core5_m0_b_corrupt(ds_cores_m0_b_corrupt[5]),
    .o_core5_m0_b_data(ds_cores_m0_b_data[5]),
    .o_core5_m0_b_mask(ds_cores_m0_b_mask[5]),
    .o_core5_m0_b_opcode(ds_cores_m0_b_opcode[5]),
    .o_core5_m0_b_param(ds_cores_m0_b_param[5]),
    .o_core5_m0_b_size(ds_cores_m0_b_size[5]),
    .o_core5_m0_b_source(ds_cores_m0_b_source[5]),
    .i_core5_m0_b_ready(ds_cores_m0_b_ready[5]),
    .o_core5_m0_b_valid(ds_cores_m0_b_valid[5]),
    .i_core5_m0_c_address(ds_cores_m0_c_address[5]),
    .i_core5_m0_c_corrupt(ds_cores_m0_c_corrupt[5]),
    .i_core5_m0_c_data(ds_cores_m0_c_data[5]),
    .i_core5_m0_c_opcode(ds_cores_m0_c_opcode[5]),
    .i_core5_m0_c_param(ds_cores_m0_c_param[5]),
    .i_core5_m0_c_size(ds_cores_m0_c_size[5]),
    .i_core5_m0_c_source(ds_cores_m0_c_source[5]),
    .i_core5_m0_c_user(ds_cores_m0_c_user[5]),
    .o_core5_m0_c_ready(ds_cores_m0_c_ready[5]),
    .i_core5_m0_c_valid(ds_cores_m0_c_valid[5]),
    .o_core5_m0_d_corrupt(ds_cores_m0_d_corrupt[5]),
    .o_core5_m0_d_data(ds_cores_m0_d_data[5]),
    .o_core5_m0_d_denied(ds_cores_m0_d_denied[5]),
    .o_core5_m0_d_opcode(ds_cores_m0_d_opcode[5]),
    .o_core5_m0_d_param(ds_cores_m0_d_param[5]),
    .o_core5_m0_d_size(ds_cores_m0_d_size[5]),
    .o_core5_m0_d_sink(ds_cores_m0_d_sink[5]),
    .o_core5_m0_d_source(ds_cores_m0_d_source[5]),
    .o_core5_m0_d_user(ds_cores_m0_d_user[5]),
    .i_core5_m0_d_ready(ds_cores_m0_d_ready[5]),
    .o_core5_m0_d_valid(ds_cores_m0_d_valid[5]),
    .i_core5_m0_e_sink(ds_cores_m0_e_sink[5]),
    .o_core5_m0_e_ready(ds_cores_m0_e_ready[5]),
    .i_core5_m0_e_valid(ds_cores_m0_e_valid[5]),
    .i_core5_m1_axi_s_araddr(ds_cores_m1_axi_araddr[5]),
    .i_core5_m1_axi_s_arburst(ds_cores_m1_axi_arburst[5]),
    .i_core5_m1_axi_s_arcache(ds_cores_m1_axi_arcache[5]),
    .i_core5_m1_axi_s_arid(ds_cores_m1_axi_arid[5]),
    .i_core5_m1_axi_s_arlen(ds_cores_m1_axi_arlen[5]),
    .i_core5_m1_axi_s_arlock(ds_cores_m1_axi_arlock[5]),
    .i_core5_m1_axi_s_arprot(ds_cores_m1_axi_arprot[5]),
    .i_core5_m1_axi_s_arsize(ds_cores_m1_axi_arsize[5]),
    .o_core5_m1_axi_s_arready(ds_cores_m1_axi_arready[5]),
    .i_core5_m1_axi_s_arvalid(ds_cores_m1_axi_arvalid[5]),
    .i_core5_m1_axi_s_awaddr(ds_cores_m1_axi_awaddr[5]),
    .i_core5_m1_axi_s_awburst(ds_cores_m1_axi_awburst[5]),
    .i_core5_m1_axi_s_awcache(ds_cores_m1_axi_awcache[5]),
    .i_core5_m1_axi_s_awid(ds_cores_m1_axi_awid[5]),
    .i_core5_m1_axi_s_awlen(ds_cores_m1_axi_awlen[5]),
    .i_core5_m1_axi_s_awlock(ds_cores_m1_axi_awlock[5]),
    .i_core5_m1_axi_s_awprot(ds_cores_m1_axi_awprot[5]),
    .i_core5_m1_axi_s_awsize(ds_cores_m1_axi_awsize[5]),
    .o_core5_m1_axi_s_awready(ds_cores_m1_axi_awready[5]),
    .i_core5_m1_axi_s_awvalid(ds_cores_m1_axi_awvalid[5]),
    .o_core5_m1_axi_s_bid(ds_cores_m1_axi_bid[5]),
    .o_core5_m1_axi_s_bresp(ds_cores_m1_axi_bresp[5]),
    .i_core5_m1_axi_s_bready(ds_cores_m1_axi_bready[5]),
    .o_core5_m1_axi_s_bvalid(ds_cores_m1_axi_bvalid[5]),
    .o_core5_m1_axi_s_rdata(ds_cores_m1_axi_rdata[5]),
    .o_core5_m1_axi_s_rid(ds_cores_m1_axi_rid[5]),
    .o_core5_m1_axi_s_rlast(ds_cores_m1_axi_rlast[5]),
    .o_core5_m1_axi_s_rresp(ds_cores_m1_axi_rresp[5]),
    .i_core5_m1_axi_s_rready(ds_cores_m1_axi_rready[5]),
    .o_core5_m1_axi_s_rvalid(ds_cores_m1_axi_rvalid[5]),
    .i_core5_m1_axi_s_wdata(ds_cores_m1_axi_wdata[5]),
    .i_core5_m1_axi_s_wlast(ds_cores_m1_axi_wlast[5]),
    .i_core5_m1_axi_s_wstrb(ds_cores_m1_axi_wstrb[5]),
    .o_core5_m1_axi_s_wready(ds_cores_m1_axi_wready[5]),
    .i_core5_m1_axi_s_wvalid(ds_cores_m1_axi_wvalid[5]),
    .i_core5_m2_a_address(ds_cores_m2_a_address[5]),
    .i_core5_m2_a_corrupt(ds_cores_m2_a_corrupt[5]),
    .i_core5_m2_a_data(ds_cores_m2_a_data[5]),
    .i_core5_m2_a_mask(ds_cores_m2_a_mask[5]),
    .i_core5_m2_a_opcode(ds_cores_m2_a_opcode[5]),
    .i_core5_m2_a_param(ds_cores_m2_a_param[5]),
    .i_core5_m2_a_size(ds_cores_m2_a_size[5]),
    .i_core5_m2_a_source(ds_cores_m2_a_source[5]),
    .i_core5_m2_a_user(ds_cores_m2_a_user[5]),
    .o_core5_m2_a_ready(ds_cores_m2_a_ready[5]),
    .i_core5_m2_a_valid(ds_cores_m2_a_valid[5]),
    .o_core5_m2_d_corrupt(ds_cores_m2_d_corrupt[5]),
    .o_core5_m2_d_data(ds_cores_m2_d_data[5]),
    .o_core5_m2_d_denied(ds_cores_m2_d_denied[5]),
    .o_core5_m2_d_opcode(ds_cores_m2_d_opcode[5]),
    .o_core5_m2_d_param(ds_cores_m2_d_param[5]),
    .o_core5_m2_d_size(ds_cores_m2_d_size[5]),
    .o_core5_m2_d_sink(ds_cores_m2_d_sink[5]),
    .o_core5_m2_d_source(ds_cores_m2_d_source[5]),
    .o_core5_m2_d_user(ds_cores_m2_d_user[5]),
    .i_core5_m2_d_ready(ds_cores_m2_d_ready[5]),
    .o_core5_m2_d_valid(ds_cores_m2_d_valid[5]),

    .i_core6_coherent_enable(ds_cores_coherent_enable[6]),
    .o_core6_coherent_state(ds_cores_coherent_state[6]),
    .i_core6_m0_a_address(ds_cores_m0_a_address[6]),
    .i_core6_m0_a_corrupt(ds_cores_m0_a_corrupt[6]),
    .i_core6_m0_a_data(ds_cores_m0_a_data[6]),
    .i_core6_m0_a_mask(ds_cores_m0_a_mask[6]),
    .i_core6_m0_a_opcode(ds_cores_m0_a_opcode[6]),
    .i_core6_m0_a_param(ds_cores_m0_a_param[6]),
    .i_core6_m0_a_size(ds_cores_m0_a_size[6]),
    .i_core6_m0_a_source(ds_cores_m0_a_source[6]),
    .i_core6_m0_a_user(ds_cores_m0_a_user[6]),
    .o_core6_m0_a_ready(ds_cores_m0_a_ready[6]),
    .i_core6_m0_a_valid(ds_cores_m0_a_valid[6]),
    .o_core6_m0_b_address(ds_cores_m0_b_address[6]),
    .o_core6_m0_b_corrupt(ds_cores_m0_b_corrupt[6]),
    .o_core6_m0_b_data(ds_cores_m0_b_data[6]),
    .o_core6_m0_b_mask(ds_cores_m0_b_mask[6]),
    .o_core6_m0_b_opcode(ds_cores_m0_b_opcode[6]),
    .o_core6_m0_b_param(ds_cores_m0_b_param[6]),
    .o_core6_m0_b_size(ds_cores_m0_b_size[6]),
    .o_core6_m0_b_source(ds_cores_m0_b_source[6]),
    .i_core6_m0_b_ready(ds_cores_m0_b_ready[6]),
    .o_core6_m0_b_valid(ds_cores_m0_b_valid[6]),
    .i_core6_m0_c_address(ds_cores_m0_c_address[6]),
    .i_core6_m0_c_corrupt(ds_cores_m0_c_corrupt[6]),
    .i_core6_m0_c_data(ds_cores_m0_c_data[6]),
    .i_core6_m0_c_opcode(ds_cores_m0_c_opcode[6]),
    .i_core6_m0_c_param(ds_cores_m0_c_param[6]),
    .i_core6_m0_c_size(ds_cores_m0_c_size[6]),
    .i_core6_m0_c_source(ds_cores_m0_c_source[6]),
    .i_core6_m0_c_user(ds_cores_m0_c_user[6]),
    .o_core6_m0_c_ready(ds_cores_m0_c_ready[6]),
    .i_core6_m0_c_valid(ds_cores_m0_c_valid[6]),
    .o_core6_m0_d_corrupt(ds_cores_m0_d_corrupt[6]),
    .o_core6_m0_d_data(ds_cores_m0_d_data[6]),
    .o_core6_m0_d_denied(ds_cores_m0_d_denied[6]),
    .o_core6_m0_d_opcode(ds_cores_m0_d_opcode[6]),
    .o_core6_m0_d_param(ds_cores_m0_d_param[6]),
    .o_core6_m0_d_size(ds_cores_m0_d_size[6]),
    .o_core6_m0_d_sink(ds_cores_m0_d_sink[6]),
    .o_core6_m0_d_source(ds_cores_m0_d_source[6]),
    .o_core6_m0_d_user(ds_cores_m0_d_user[6]),
    .i_core6_m0_d_ready(ds_cores_m0_d_ready[6]),
    .o_core6_m0_d_valid(ds_cores_m0_d_valid[6]),
    .i_core6_m0_e_sink(ds_cores_m0_e_sink[6]),
    .o_core6_m0_e_ready(ds_cores_m0_e_ready[6]),
    .i_core6_m0_e_valid(ds_cores_m0_e_valid[6]),
    .i_core6_m1_axi_s_araddr(ds_cores_m1_axi_araddr[6]),
    .i_core6_m1_axi_s_arburst(ds_cores_m1_axi_arburst[6]),
    .i_core6_m1_axi_s_arcache(ds_cores_m1_axi_arcache[6]),
    .i_core6_m1_axi_s_arid(ds_cores_m1_axi_arid[6]),
    .i_core6_m1_axi_s_arlen(ds_cores_m1_axi_arlen[6]),
    .i_core6_m1_axi_s_arlock(ds_cores_m1_axi_arlock[6]),
    .i_core6_m1_axi_s_arprot(ds_cores_m1_axi_arprot[6]),
    .i_core6_m1_axi_s_arsize(ds_cores_m1_axi_arsize[6]),
    .o_core6_m1_axi_s_arready(ds_cores_m1_axi_arready[6]),
    .i_core6_m1_axi_s_arvalid(ds_cores_m1_axi_arvalid[6]),
    .i_core6_m1_axi_s_awaddr(ds_cores_m1_axi_awaddr[6]),
    .i_core6_m1_axi_s_awburst(ds_cores_m1_axi_awburst[6]),
    .i_core6_m1_axi_s_awcache(ds_cores_m1_axi_awcache[6]),
    .i_core6_m1_axi_s_awid(ds_cores_m1_axi_awid[6]),
    .i_core6_m1_axi_s_awlen(ds_cores_m1_axi_awlen[6]),
    .i_core6_m1_axi_s_awlock(ds_cores_m1_axi_awlock[6]),
    .i_core6_m1_axi_s_awprot(ds_cores_m1_axi_awprot[6]),
    .i_core6_m1_axi_s_awsize(ds_cores_m1_axi_awsize[6]),
    .o_core6_m1_axi_s_awready(ds_cores_m1_axi_awready[6]),
    .i_core6_m1_axi_s_awvalid(ds_cores_m1_axi_awvalid[6]),
    .o_core6_m1_axi_s_bid(ds_cores_m1_axi_bid[6]),
    .o_core6_m1_axi_s_bresp(ds_cores_m1_axi_bresp[6]),
    .i_core6_m1_axi_s_bready(ds_cores_m1_axi_bready[6]),
    .o_core6_m1_axi_s_bvalid(ds_cores_m1_axi_bvalid[6]),
    .o_core6_m1_axi_s_rdata(ds_cores_m1_axi_rdata[6]),
    .o_core6_m1_axi_s_rid(ds_cores_m1_axi_rid[6]),
    .o_core6_m1_axi_s_rlast(ds_cores_m1_axi_rlast[6]),
    .o_core6_m1_axi_s_rresp(ds_cores_m1_axi_rresp[6]),
    .i_core6_m1_axi_s_rready(ds_cores_m1_axi_rready[6]),
    .o_core6_m1_axi_s_rvalid(ds_cores_m1_axi_rvalid[6]),
    .i_core6_m1_axi_s_wdata(ds_cores_m1_axi_wdata[6]),
    .i_core6_m1_axi_s_wlast(ds_cores_m1_axi_wlast[6]),
    .i_core6_m1_axi_s_wstrb(ds_cores_m1_axi_wstrb[6]),
    .o_core6_m1_axi_s_wready(ds_cores_m1_axi_wready[6]),
    .i_core6_m1_axi_s_wvalid(ds_cores_m1_axi_wvalid[6]),
    .i_core6_m2_a_address(ds_cores_m2_a_address[6]),
    .i_core6_m2_a_corrupt(ds_cores_m2_a_corrupt[6]),
    .i_core6_m2_a_data(ds_cores_m2_a_data[6]),
    .i_core6_m2_a_mask(ds_cores_m2_a_mask[6]),
    .i_core6_m2_a_opcode(ds_cores_m2_a_opcode[6]),
    .i_core6_m2_a_param(ds_cores_m2_a_param[6]),
    .i_core6_m2_a_size(ds_cores_m2_a_size[6]),
    .i_core6_m2_a_source(ds_cores_m2_a_source[6]),
    .i_core6_m2_a_user(ds_cores_m2_a_user[6]),
    .o_core6_m2_a_ready(ds_cores_m2_a_ready[6]),
    .i_core6_m2_a_valid(ds_cores_m2_a_valid[6]),
    .o_core6_m2_d_corrupt(ds_cores_m2_d_corrupt[6]),
    .o_core6_m2_d_data(ds_cores_m2_d_data[6]),
    .o_core6_m2_d_denied(ds_cores_m2_d_denied[6]),
    .o_core6_m2_d_opcode(ds_cores_m2_d_opcode[6]),
    .o_core6_m2_d_param(ds_cores_m2_d_param[6]),
    .o_core6_m2_d_size(ds_cores_m2_d_size[6]),
    .o_core6_m2_d_sink(ds_cores_m2_d_sink[6]),
    .o_core6_m2_d_source(ds_cores_m2_d_source[6]),
    .o_core6_m2_d_user(ds_cores_m2_d_user[6]),
    .i_core6_m2_d_ready(ds_cores_m2_d_ready[6]),
    .o_core6_m2_d_valid(ds_cores_m2_d_valid[6]),

    .i_core7_coherent_enable(ds_cores_coherent_enable[7]),
    .o_core7_coherent_state(ds_cores_coherent_state[7]),
    .i_core7_m0_a_address(ds_cores_m0_a_address[7]),
    .i_core7_m0_a_corrupt(ds_cores_m0_a_corrupt[7]),
    .i_core7_m0_a_data(ds_cores_m0_a_data[7]),
    .i_core7_m0_a_mask(ds_cores_m0_a_mask[7]),
    .i_core7_m0_a_opcode(ds_cores_m0_a_opcode[7]),
    .i_core7_m0_a_param(ds_cores_m0_a_param[7]),
    .i_core7_m0_a_size(ds_cores_m0_a_size[7]),
    .i_core7_m0_a_source(ds_cores_m0_a_source[7]),
    .i_core7_m0_a_user(ds_cores_m0_a_user[7]),
    .o_core7_m0_a_ready(ds_cores_m0_a_ready[7]),
    .i_core7_m0_a_valid(ds_cores_m0_a_valid[7]),
    .o_core7_m0_b_address(ds_cores_m0_b_address[7]),
    .o_core7_m0_b_corrupt(ds_cores_m0_b_corrupt[7]),
    .o_core7_m0_b_data(ds_cores_m0_b_data[7]),
    .o_core7_m0_b_mask(ds_cores_m0_b_mask[7]),
    .o_core7_m0_b_opcode(ds_cores_m0_b_opcode[7]),
    .o_core7_m0_b_param(ds_cores_m0_b_param[7]),
    .o_core7_m0_b_size(ds_cores_m0_b_size[7]),
    .o_core7_m0_b_source(ds_cores_m0_b_source[7]),
    .i_core7_m0_b_ready(ds_cores_m0_b_ready[7]),
    .o_core7_m0_b_valid(ds_cores_m0_b_valid[7]),
    .i_core7_m0_c_address(ds_cores_m0_c_address[7]),
    .i_core7_m0_c_corrupt(ds_cores_m0_c_corrupt[7]),
    .i_core7_m0_c_data(ds_cores_m0_c_data[7]),
    .i_core7_m0_c_opcode(ds_cores_m0_c_opcode[7]),
    .i_core7_m0_c_param(ds_cores_m0_c_param[7]),
    .i_core7_m0_c_size(ds_cores_m0_c_size[7]),
    .i_core7_m0_c_source(ds_cores_m0_c_source[7]),
    .i_core7_m0_c_user(ds_cores_m0_c_user[7]),
    .o_core7_m0_c_ready(ds_cores_m0_c_ready[7]),
    .i_core7_m0_c_valid(ds_cores_m0_c_valid[7]),
    .o_core7_m0_d_corrupt(ds_cores_m0_d_corrupt[7]),
    .o_core7_m0_d_data(ds_cores_m0_d_data[7]),
    .o_core7_m0_d_denied(ds_cores_m0_d_denied[7]),
    .o_core7_m0_d_opcode(ds_cores_m0_d_opcode[7]),
    .o_core7_m0_d_param(ds_cores_m0_d_param[7]),
    .o_core7_m0_d_size(ds_cores_m0_d_size[7]),
    .o_core7_m0_d_sink(ds_cores_m0_d_sink[7]),
    .o_core7_m0_d_source(ds_cores_m0_d_source[7]),
    .o_core7_m0_d_user(ds_cores_m0_d_user[7]),
    .i_core7_m0_d_ready(ds_cores_m0_d_ready[7]),
    .o_core7_m0_d_valid(ds_cores_m0_d_valid[7]),
    .i_core7_m0_e_sink(ds_cores_m0_e_sink[7]),
    .o_core7_m0_e_ready(ds_cores_m0_e_ready[7]),
    .i_core7_m0_e_valid(ds_cores_m0_e_valid[7]),
    .i_core7_m1_axi_s_araddr(ds_cores_m1_axi_araddr[7]),
    .i_core7_m1_axi_s_arburst(ds_cores_m1_axi_arburst[7]),
    .i_core7_m1_axi_s_arcache(ds_cores_m1_axi_arcache[7]),
    .i_core7_m1_axi_s_arid(ds_cores_m1_axi_arid[7]),
    .i_core7_m1_axi_s_arlen(ds_cores_m1_axi_arlen[7]),
    .i_core7_m1_axi_s_arlock(ds_cores_m1_axi_arlock[7]),
    .i_core7_m1_axi_s_arprot(ds_cores_m1_axi_arprot[7]),
    .i_core7_m1_axi_s_arsize(ds_cores_m1_axi_arsize[7]),
    .o_core7_m1_axi_s_arready(ds_cores_m1_axi_arready[7]),
    .i_core7_m1_axi_s_arvalid(ds_cores_m1_axi_arvalid[7]),
    .i_core7_m1_axi_s_awaddr(ds_cores_m1_axi_awaddr[7]),
    .i_core7_m1_axi_s_awburst(ds_cores_m1_axi_awburst[7]),
    .i_core7_m1_axi_s_awcache(ds_cores_m1_axi_awcache[7]),
    .i_core7_m1_axi_s_awid(ds_cores_m1_axi_awid[7]),
    .i_core7_m1_axi_s_awlen(ds_cores_m1_axi_awlen[7]),
    .i_core7_m1_axi_s_awlock(ds_cores_m1_axi_awlock[7]),
    .i_core7_m1_axi_s_awprot(ds_cores_m1_axi_awprot[7]),
    .i_core7_m1_axi_s_awsize(ds_cores_m1_axi_awsize[7]),
    .o_core7_m1_axi_s_awready(ds_cores_m1_axi_awready[7]),
    .i_core7_m1_axi_s_awvalid(ds_cores_m1_axi_awvalid[7]),
    .o_core7_m1_axi_s_bid(ds_cores_m1_axi_bid[7]),
    .o_core7_m1_axi_s_bresp(ds_cores_m1_axi_bresp[7]),
    .i_core7_m1_axi_s_bready(ds_cores_m1_axi_bready[7]),
    .o_core7_m1_axi_s_bvalid(ds_cores_m1_axi_bvalid[7]),
    .o_core7_m1_axi_s_rdata(ds_cores_m1_axi_rdata[7]),
    .o_core7_m1_axi_s_rid(ds_cores_m1_axi_rid[7]),
    .o_core7_m1_axi_s_rlast(ds_cores_m1_axi_rlast[7]),
    .o_core7_m1_axi_s_rresp(ds_cores_m1_axi_rresp[7]),
    .i_core7_m1_axi_s_rready(ds_cores_m1_axi_rready[7]),
    .o_core7_m1_axi_s_rvalid(ds_cores_m1_axi_rvalid[7]),
    .i_core7_m1_axi_s_wdata(ds_cores_m1_axi_wdata[7]),
    .i_core7_m1_axi_s_wlast(ds_cores_m1_axi_wlast[7]),
    .i_core7_m1_axi_s_wstrb(ds_cores_m1_axi_wstrb[7]),
    .o_core7_m1_axi_s_wready(ds_cores_m1_axi_wready[7]),
    .i_core7_m1_axi_s_wvalid(ds_cores_m1_axi_wvalid[7]),
    .i_core7_m2_a_address(ds_cores_m2_a_address[7]),
    .i_core7_m2_a_corrupt(ds_cores_m2_a_corrupt[7]),
    .i_core7_m2_a_data(ds_cores_m2_a_data[7]),
    .i_core7_m2_a_mask(ds_cores_m2_a_mask[7]),
    .i_core7_m2_a_opcode(ds_cores_m2_a_opcode[7]),
    .i_core7_m2_a_param(ds_cores_m2_a_param[7]),
    .i_core7_m2_a_size(ds_cores_m2_a_size[7]),
    .i_core7_m2_a_source(ds_cores_m2_a_source[7]),
    .i_core7_m2_a_user(ds_cores_m2_a_user[7]),
    .o_core7_m2_a_ready(ds_cores_m2_a_ready[7]),
    .i_core7_m2_a_valid(ds_cores_m2_a_valid[7]),
    .o_core7_m2_d_corrupt(ds_cores_m2_d_corrupt[7]),
    .o_core7_m2_d_data(ds_cores_m2_d_data[7]),
    .o_core7_m2_d_denied(ds_cores_m2_d_denied[7]),
    .o_core7_m2_d_opcode(ds_cores_m2_d_opcode[7]),
    .o_core7_m2_d_param(ds_cores_m2_d_param[7]),
    .o_core7_m2_d_size(ds_cores_m2_d_size[7]),
    .o_core7_m2_d_sink(ds_cores_m2_d_sink[7]),
    .o_core7_m2_d_source(ds_cores_m2_d_source[7]),
    .o_core7_m2_d_user(ds_cores_m2_d_user[7]),
    .i_core7_m2_d_ready(ds_cores_m2_d_ready[7]),
    .o_core7_m2_d_valid(ds_cores_m2_d_valid[7]),

    //////////////////////////////////////////////
    /// AXI sigs
    //////////////////////////////////////////////
    .i_iocp_axi_s_araddr(i_iocp_axi_s_ar.addr),
    .i_iocp_axi_s_arburst(i_iocp_axi_s_ar.burst),
    .i_iocp_axi_s_arcache(i_iocp_axi_s_ar.cache),
    .i_iocp_axi_s_arid(i_iocp_axi_s_ar.id),
    .i_iocp_axi_s_arlen(i_iocp_axi_s_ar.len),
    .i_iocp_axi_s_arlock(i_iocp_axi_s_ar.lock),
    .i_iocp_axi_s_arprot(i_iocp_axi_s_ar.prot),
    .i_iocp_axi_s_arsize(i_iocp_axi_s_ar.size),
    .o_iocp_axi_s_arready,
    .i_iocp_axi_s_arvalid,
    .i_iocp_axi_s_awaddr(i_iocp_axi_s_aw.addr),
    .i_iocp_axi_s_awburst(i_iocp_axi_s_aw.burst),
    .i_iocp_axi_s_awcache(i_iocp_axi_s_aw.cache),
    .i_iocp_axi_s_awid(i_iocp_axi_s_aw.id),
    .i_iocp_axi_s_awlen(i_iocp_axi_s_aw.len),
    .i_iocp_axi_s_awlock(i_iocp_axi_s_aw.lock),
    .i_iocp_axi_s_awprot(i_iocp_axi_s_aw.prot),
    .i_iocp_axi_s_awsize(i_iocp_axi_s_aw.size),
    .o_iocp_axi_s_awready,
    .i_iocp_axi_s_awvalid,
    .o_iocp_axi_s_bid(o_iocp_axi_s_b.id),
    .o_iocp_axi_s_bresp(o_iocp_axi_s_b.resp[axi_pkg::AXI_RESP_WIDTH-1:0]),
    .i_iocp_axi_s_bready,
    .o_iocp_axi_s_bvalid,
    .o_iocp_axi_s_rdata(o_iocp_axi_s_r.data),
    .o_iocp_axi_s_rid(o_iocp_axi_s_r.id),
    .o_iocp_axi_s_rlast(o_iocp_axi_s_r.last),
    .o_iocp_axi_s_rresp(o_iocp_axi_s_r.resp[axi_pkg::AXI_RESP_WIDTH-1:0]),
    .i_iocp_axi_s_rready,
    .o_iocp_axi_s_rvalid,
    .i_iocp_axi_s_wdata(i_iocp_axi_s_w.data),
    .i_iocp_axi_s_wlast(i_iocp_axi_s_w.last),
    .i_iocp_axi_s_wstrb(i_iocp_axi_s_w.strb),
    .o_iocp_axi_s_wready,
    .i_iocp_axi_s_wvalid,
    .o_mem_axi_m_araddr(o_mem_axi_m_ar.addr),
    .o_mem_axi_m_arburst(o_mem_axi_m_ar.burst[axi_pkg::AXI_BURST_WIDTH-1:0]),
    .o_mem_axi_m_arcache(o_mem_axi_m_ar.cache),
    .o_mem_axi_m_arid(o_mem_axi_m_ar.id),
    .o_mem_axi_m_arlen(o_mem_axi_m_ar.len),
    .o_mem_axi_m_arlock(o_mem_axi_m_ar.lock),
    .o_mem_axi_m_arprot(o_mem_axi_m_ar.prot),
    .o_mem_axi_m_arsize(o_mem_axi_m_ar.size[axi_pkg::AXI_SIZE_WIDTH-1:0]),
    .i_mem_axi_m_arready,
    .o_mem_axi_m_arvalid,
    .o_mem_axi_m_awaddr(o_mem_axi_m_aw.addr),
    .o_mem_axi_m_awburst(o_mem_axi_m_aw.burst[axi_pkg::AXI_BURST_WIDTH-1:0]),
    .o_mem_axi_m_awcache(o_mem_axi_m_aw.cache),
    .o_mem_axi_m_awid(o_mem_axi_m_aw.id),
    .o_mem_axi_m_awlen(o_mem_axi_m_aw.len),
    .o_mem_axi_m_awlock(o_mem_axi_m_aw.lock),
    .o_mem_axi_m_awprot(o_mem_axi_m_aw.prot),
    .o_mem_axi_m_awsize(o_mem_axi_m_aw.size[axi_pkg::AXI_SIZE_WIDTH-1:0]),
    .i_mem_axi_m_awready,
    .o_mem_axi_m_awvalid,
    .i_mem_axi_m_bid(i_mem_axi_m_b.id),
    .i_mem_axi_m_bresp(i_mem_axi_m_b.resp),
    .o_mem_axi_m_bready,
    .i_mem_axi_m_bvalid,
    .i_mem_axi_m_rdata(i_mem_axi_m_r.data),
    .i_mem_axi_m_rid(i_mem_axi_m_r.id),
    .i_mem_axi_m_rlast(i_mem_axi_m_r.last),
    .i_mem_axi_m_rresp(i_mem_axi_m_r.resp),
    .o_mem_axi_m_rready,
    .i_mem_axi_m_rvalid,
    .o_mem_axi_m_wdata(o_mem_axi_m_w.data),
    .o_mem_axi_m_wlast(o_mem_axi_m_w.last),
    .o_mem_axi_m_wstrb(o_mem_axi_m_w.strb),
    .i_mem_axi_m_wready,
    .o_mem_axi_m_wvalid,
    .o_mmio_axi_m_araddr(o_mmio_axi_m_ar.addr),
    .o_mmio_axi_m_arburst(o_mmio_axi_m_ar.burst[axi_pkg::AXI_BURST_WIDTH-1:0]),
    .o_mmio_axi_m_arcache(o_mmio_axi_m_ar.cache),
    .o_mmio_axi_m_arid(o_mmio_axi_m_ar.id),
    .o_mmio_axi_m_arlen(o_mmio_axi_m_ar.len),
    .o_mmio_axi_m_arlock(o_mmio_axi_m_ar.lock),
    .o_mmio_axi_m_arprot(o_mmio_axi_m_ar.prot),
    .o_mmio_axi_m_arsize(o_mmio_axi_m_ar.size[axi_pkg::AXI_SIZE_WIDTH-1:0]),
    .i_mmio_axi_m_arready,
    .o_mmio_axi_m_arvalid,
    .o_mmio_axi_m_awaddr(o_mmio_axi_m_aw.addr),
    .o_mmio_axi_m_awburst(o_mmio_axi_m_aw.burst[axi_pkg::AXI_BURST_WIDTH-1:0]),
    .o_mmio_axi_m_awcache(o_mmio_axi_m_aw.cache),
    .o_mmio_axi_m_awid(o_mmio_axi_m_aw.id),
    .o_mmio_axi_m_awlen(o_mmio_axi_m_aw.len),
    .o_mmio_axi_m_awlock(o_mmio_axi_m_aw.lock),
    .o_mmio_axi_m_awprot(o_mmio_axi_m_aw.prot),
    .o_mmio_axi_m_awsize(o_mmio_axi_m_aw.size[axi_pkg::AXI_SIZE_WIDTH-1:0]),
    .i_mmio_axi_m_awready,
    .o_mmio_axi_m_awvalid,
    .i_mmio_axi_m_bid(i_mmio_axi_m_b.id),
    .i_mmio_axi_m_bresp(i_mmio_axi_m_b.resp),
    .o_mmio_axi_m_bready,
    .i_mmio_axi_m_bvalid,
    .i_mmio_axi_m_rdata(i_mmio_axi_m_r.data),
    .i_mmio_axi_m_rid(i_mmio_axi_m_r.id),
    .i_mmio_axi_m_rlast(i_mmio_axi_m_r.last),
    .i_mmio_axi_m_rresp(i_mmio_axi_m_r.resp),
    .o_mmio_axi_m_rready,
    .i_mmio_axi_m_rvalid,
    .o_mmio_axi_m_wdata(o_mmio_axi_m_w.data),
    .o_mmio_axi_m_wlast(o_mmio_axi_m_w.last),
    .o_mmio_axi_m_wstrb(o_mmio_axi_m_w.strb),
    .i_mmio_axi_m_wready,
    .o_mmio_axi_m_wvalid,
    .o_plmt_axi_m_araddr(plmt_axi_ar.addr),
    .o_plmt_axi_m_arburst(plmt_axi_ar.burst[axi_pkg::AXI_BURST_WIDTH-1:0]),
    .o_plmt_axi_m_arcache(plmt_axi_ar.cache),
    .o_plmt_axi_m_arid(plmt_axi_ar.id),
    .o_plmt_axi_m_arlen(plmt_axi_ar.len),
    .o_plmt_axi_m_arlock(plmt_axi_ar.lock),
    .o_plmt_axi_m_arprot(plmt_axi_ar.prot),
    .o_plmt_axi_m_arsize(plmt_axi_ar.size[axi_pkg::AXI_SIZE_WIDTH-1:0]),
    .i_plmt_axi_m_arready(plmt_axi_arready),
    .o_plmt_axi_m_arvalid(plmt_axi_arvalid),
    .o_plmt_axi_m_awaddr(plmt_axi_aw.addr),
    .o_plmt_axi_m_awburst(plmt_axi_aw.burst[axi_pkg::AXI_BURST_WIDTH-1:0]),
    .o_plmt_axi_m_awcache(plmt_axi_aw.cache),
    .o_plmt_axi_m_awid(plmt_axi_aw.id),
    .o_plmt_axi_m_awlen(plmt_axi_aw.len),
    .o_plmt_axi_m_awlock(plmt_axi_aw.lock),
    .o_plmt_axi_m_awprot(plmt_axi_aw.prot),
    .o_plmt_axi_m_awsize(plmt_axi_aw.size[axi_pkg::AXI_SIZE_WIDTH-1:0]),
    .i_plmt_axi_m_awready(plmt_axi_awready),
    .o_plmt_axi_m_awvalid(plmt_axi_awvalid),
    .i_plmt_axi_m_bid(plmt_axi_b.id),
    .i_plmt_axi_m_bresp(plmt_axi_b.resp),
    .o_plmt_axi_m_bready(plmt_axi_bready),
    .i_plmt_axi_m_bvalid(plmt_axi_bvalid),
    .i_plmt_axi_m_rdata(plmt_axi_r.data),
    .i_plmt_axi_m_rid(plmt_axi_r.id),
    .i_plmt_axi_m_rlast(plmt_axi_r.last),
    .i_plmt_axi_m_rresp(plmt_axi_r.resp),
    .o_plmt_axi_m_rready(plmt_axi_rready),
    .i_plmt_axi_m_rvalid(plmt_axi_rvalid),
    .o_plmt_axi_m_wdata(plmt_axi_w.data),
    .o_plmt_axi_m_wlast(plmt_axi_w.last),
    .o_plmt_axi_m_wstrb(plmt_axi_w.strb),
    .i_plmt_axi_m_wready(plmt_axi_wready),
    .o_plmt_axi_m_wvalid(plmt_axi_wvalid),
    //////////////////////////////////////////////
    /// L2C bank sigs
    //////////////////////////////////////////////
    .i_l2c_ctrl,
    .o_l2c_ctrl,
    .i_l2c_disable_init,
    .o_l2c_err_int
  );

  // Drive AXI optional to 0
  always_comb o_mem_axi_m_ar.qos    = 'b0;
  always_comb o_mem_axi_m_ar.region = 'b0;
  always_comb o_mem_axi_m_ar.user   = 'b0;
  always_comb o_mem_axi_m_aw.atop   = 'b0;
  always_comb o_mem_axi_m_aw.qos    = 'b0;
  always_comb o_mem_axi_m_aw.region = 'b0;
  always_comb o_mem_axi_m_aw.user   = 'b0;
  always_comb o_mem_axi_m_w.user    = 'b0;

  always_comb o_mmio_axi_m_ar.qos    = 'b0;
  always_comb o_mmio_axi_m_ar.region = 'b0;
  always_comb o_mmio_axi_m_ar.user   = 'b0;
  always_comb o_mmio_axi_m_aw.atop   = 'b0;
  always_comb o_mmio_axi_m_aw.qos    = 'b0;
  always_comb o_mmio_axi_m_aw.region = 'b0;
  always_comb o_mmio_axi_m_aw.user   = 'b0;
  always_comb o_mmio_axi_m_w.user    = 'b0;

  ax65_peripheral_wrapper #(
    .CORE_WIDTH(CORE_WIDTH + APU_AIC_WIDTH),
    .ADDR_WIDTH(chip_pkg::CHIP_AXI_ADDR_W),
    .DATA_WIDTH(chip_pkg::CHIP_AXI_LT_DATA_W),
    .ID_WIDTH(APU_AXI_LT_M_ID_W)
  ) u_peripheral_wrapper (
    .i_aclk,
    .i_arst_n,
    .i_mtime_clk,
    .i_por_rst_n,
    .o_cores_mtip(all_cores_mtip),
    .i_cores_stoptime(all_cores_stoptime),
    .i_test_mode,
    .i_plmt_axi_s_araddr(plmt_axi_ar.addr),
    .i_plmt_axi_s_arburst(plmt_axi_ar.burst),
    .i_plmt_axi_s_arcache(plmt_axi_ar.cache),
    .i_plmt_axi_s_arid(plmt_axi_ar.id),
    .i_plmt_axi_s_arlen(plmt_axi_ar.len),
    .i_plmt_axi_s_arlock(plmt_axi_ar.lock),
    .i_plmt_axi_s_arprot(plmt_axi_ar.prot),
    .i_plmt_axi_s_arsize(plmt_axi_ar.size),
    .o_plmt_axi_s_arready(plmt_axi_arready),
    .i_plmt_axi_s_arvalid(plmt_axi_arvalid),
    .i_plmt_axi_s_awaddr(plmt_axi_aw.addr),
    .i_plmt_axi_s_awburst(plmt_axi_aw.burst),
    .i_plmt_axi_s_awcache(plmt_axi_aw.cache),
    .i_plmt_axi_s_awid(plmt_axi_aw.id),
    .i_plmt_axi_s_awlen(plmt_axi_aw.len),
    .i_plmt_axi_s_awlock(plmt_axi_aw.lock),
    .i_plmt_axi_s_awprot(plmt_axi_aw.prot),
    .i_plmt_axi_s_awsize(plmt_axi_aw.size),
    .o_plmt_axi_s_awready(plmt_axi_awready),
    .i_plmt_axi_s_awvalid(plmt_axi_awvalid),
    .o_plmt_axi_s_bid(plmt_axi_b.id),
    .o_plmt_axi_s_bresp(plmt_axi_b.resp[axi_pkg::AXI_RESP_WIDTH-1:0]),
    .i_plmt_axi_s_bready(plmt_axi_bready),
    .o_plmt_axi_s_bvalid(plmt_axi_bvalid),
    .o_plmt_axi_s_rdata(plmt_axi_r.data),
    .o_plmt_axi_s_rid(plmt_axi_r.id),
    .o_plmt_axi_s_rlast(plmt_axi_r.last),
    .o_plmt_axi_s_rresp(plmt_axi_r.resp[axi_pkg::AXI_RESP_WIDTH-1:0]),
    .i_plmt_axi_s_rready(plmt_axi_rready),
    .o_plmt_axi_s_rvalid(plmt_axi_rvalid),
    .i_plmt_axi_s_wdata(plmt_axi_w.data),
    .i_plmt_axi_s_wlast(plmt_axi_w.last),
    .i_plmt_axi_s_wstrb(plmt_axi_w.strb),
    .o_plmt_axi_s_wready(plmt_axi_wready),
    .i_plmt_axi_s_wvalid(plmt_axi_wvalid)
  );

endmodule
