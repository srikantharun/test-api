
// (C) Copyright 2025 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_noc_tok_v_center
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_tok_v_center (
  output logic [41:0] o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld,
  input wire  i_noc_clk,
  input wire  i_noc_rst_n,
  input logic  scan_en,
  input wire  i_sdma_0_clk,
  input wire  i_sdma_0_clken,
  input logic [7:0] i_sdma_0_init_tok_ocpl_s_maddr,
  input logic [2:0] i_sdma_0_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_sdma_0_init_tok_ocpl_s_mdata,
  output logic  o_sdma_0_init_tok_ocpl_s_scmdaccept,
  output logic  o_sdma_0_pwr_tok_idle_val,
  output logic  o_sdma_0_pwr_tok_idle_ack,
  input logic  i_sdma_0_pwr_tok_idle_req,
  input wire  i_sdma_0_rst_n,
  output logic [7:0] o_sdma_0_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_sdma_0_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_sdma_0_targ_tok_ocpl_m_mdata,
  input logic  i_sdma_0_targ_tok_ocpl_m_scmdaccept,
  input wire  i_sdma_1_clk,
  input wire  i_sdma_1_clken,
  input logic [7:0] i_sdma_1_init_tok_ocpl_s_maddr,
  input logic [2:0] i_sdma_1_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_sdma_1_init_tok_ocpl_s_mdata,
  output logic  o_sdma_1_init_tok_ocpl_s_scmdaccept,
  output logic  o_sdma_1_pwr_tok_idle_val,
  output logic  o_sdma_1_pwr_tok_idle_ack,
  input logic  i_sdma_1_pwr_tok_idle_req,
  input wire  i_sdma_1_rst_n,
  output logic [7:0] o_sdma_1_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_sdma_1_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_sdma_1_targ_tok_ocpl_m_mdata,
  input logic  i_sdma_1_targ_tok_ocpl_m_scmdaccept
);

noc_tok_art_v_center u_noc_tok_art_v_center (
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Data(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data),
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Head(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head),
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Rdy(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy),
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Tail(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail),
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Vld(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Data(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Head(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Rdy(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Tail(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Vld(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Data(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Head(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Rdy(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Tail(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Vld(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Data(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Head(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Rdy(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Tail(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Vld(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Data(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Head(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Rdy(i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Tail(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail),
  .dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_Vld(o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Data(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Head(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Rdy(i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Tail(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail),
  .dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_Vld(o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Data(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Head(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Rdy(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Tail(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Vld(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Data(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Head(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Rdy(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Tail(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Vld(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Data(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Head(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Rdy(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Tail(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Vld(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Data(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Head(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Rdy(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Tail(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Vld(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Data(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Head(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Rdy(o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Tail(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail),
  .dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_Vld(i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Data(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Head(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Rdy(o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Tail(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail),
  .dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_Vld(i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld),
  .noc_clk(i_noc_clk),
  .noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en),
  .sdma_0_clk(i_sdma_0_clk),
  .sdma_0_clken(i_sdma_0_clken),
  .sdma_0_init_tok_MAddr(i_sdma_0_init_tok_ocpl_s_maddr),
  .sdma_0_init_tok_MCmd(i_sdma_0_init_tok_ocpl_s_mcmd),
  .sdma_0_init_tok_MData(i_sdma_0_init_tok_ocpl_s_mdata),
  .sdma_0_init_tok_SCmdAccept(o_sdma_0_init_tok_ocpl_s_scmdaccept),
  .sdma_0_pwr_tok_Idle(o_sdma_0_pwr_tok_idle_val),
  .sdma_0_pwr_tok_IdleAck(o_sdma_0_pwr_tok_idle_ack),
  .sdma_0_pwr_tok_IdleReq(i_sdma_0_pwr_tok_idle_req),
  .sdma_0_rst_n(i_sdma_0_rst_n),
  .sdma_0_targ_tok_MAddr(o_sdma_0_targ_tok_ocpl_m_maddr),
  .sdma_0_targ_tok_MCmd(o_sdma_0_targ_tok_ocpl_m_mcmd),
  .sdma_0_targ_tok_MData(o_sdma_0_targ_tok_ocpl_m_mdata),
  .sdma_0_targ_tok_SCmdAccept(i_sdma_0_targ_tok_ocpl_m_scmdaccept),
  .sdma_1_clk(i_sdma_1_clk),
  .sdma_1_clken(i_sdma_1_clken),
  .sdma_1_init_tok_MAddr(i_sdma_1_init_tok_ocpl_s_maddr),
  .sdma_1_init_tok_MCmd(i_sdma_1_init_tok_ocpl_s_mcmd),
  .sdma_1_init_tok_MData(i_sdma_1_init_tok_ocpl_s_mdata),
  .sdma_1_init_tok_SCmdAccept(o_sdma_1_init_tok_ocpl_s_scmdaccept),
  .sdma_1_pwr_tok_Idle(o_sdma_1_pwr_tok_idle_val),
  .sdma_1_pwr_tok_IdleAck(o_sdma_1_pwr_tok_idle_ack),
  .sdma_1_pwr_tok_IdleReq(i_sdma_1_pwr_tok_idle_req),
  .sdma_1_rst_n(i_sdma_1_rst_n),
  .sdma_1_targ_tok_MAddr(o_sdma_1_targ_tok_ocpl_m_maddr),
  .sdma_1_targ_tok_MCmd(o_sdma_1_targ_tok_ocpl_m_mcmd),
  .sdma_1_targ_tok_MData(o_sdma_1_targ_tok_ocpl_m_mdata),
  .sdma_1_targ_tok_SCmdAccept(i_sdma_1_targ_tok_ocpl_m_scmdaccept)
);
endmodule
