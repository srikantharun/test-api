 import lpddr_axi_pkg::*;

 bind lpddr_p Axi4PC # (
				.DATA_WIDTH(512),
        .ADDR_WIDTH(36),
				.RID_WIDTH  (8),
				.WID_WIDTH  (8),
        .MAXWBURSTS(20),
        .MAXRBURSTS(20),
        .RecommendOn(0),
				.RecMaxWaitOn( 0 ),
        .AWREADY_MAXWAITS ( 50 ),
        .ARREADY_MAXWAITS ( 50 ),
        .WREADY_MAXWAITS ( 50 ),
        .BREADY_MAXWAITS ( 16 ),
        .RREADY_MAXWAITS ( 16 )
				)
	AXI_AIP_DDR_axi_hp_s
				(
				.ACLK(lpddr_ctrl_axi_s_aclk),
				.ARESETn(lpddr_ctrl_axi_s_aclk),
				.ARVALID(lpddr_ctrl_axi_s_arvalid),
				.ARADDR(lpddr_ctrl_axi_s_araddr ),
				.ARLEN(lpddr_ctrl_axi_s_arlen),
				.ARSIZE( lpddr_ctrl_axi_s_arsize),
				.ARBURST( lpddr_ctrl_axi_s_arburst ),
				.ARLOCK( lpddr_ctrl_axi_s_arlock),
				.ARCACHE( lpddr_ctrl_axi_s_arcache ),
				.ARPROT( lpddr_ctrl_axi_s_arprot ),
				.ARID( lpddr_ctrl_axi_s_arid ),
				.ARREADY( lpddr_ctrl_axi_s_arready ),
				.RREADY( lpddr_ctrl_axi_s_rready ),
				.RVALID( lpddr_ctrl_axi_s_rvalid ),
				.RLAST( lpddr_ctrl_axi_s_rlast ),
				.RDATA( lpddr_ctrl_axi_s_rdata ),
				.RRESP( lpddr_ctrl_axi_s_rresp ),
				.RID( lpddr_ctrl_axi_s_rid ),
				.AWVALID( lpddr_ctrl_axi_s_awvalid ),
				.AWADDR( lpddr_ctrl_axi_s_awaddr ),
				.AWLEN( lpddr_ctrl_axi_s_awlen),
				.AWSIZE( lpddr_ctrl_axi_s_awsize ),
				.AWBURST( lpddr_ctrl_axi_s_awburst ),
				.AWLOCK( lpddr_ctrl_axi_s_awlock ),
				.AWCACHE( lpddr_ctrl_axi_s_awcache ),
				.AWPROT( lpddr_ctrl_axi_s_awprot ),
				.AWID( lpddr_ctrl_axi_s_awid ),
				.AWREADY( lpddr_ctrl_axi_s_awready ),
				.WVALID( lpddr_ctrl_axi_s_wvalid ),
				.WLAST( lpddr_ctrl_axi_s_wlast ),
				.WDATA( lpddr_ctrl_axi_s_wdata ),
				.WSTRB( lpddr_ctrl_axi_s_wstrb ),
				.WREADY( lpddr_ctrl_axi_s_wready),
				.BREADY( lpddr_ctrl_axi_s_bready ),
				.BVALID( lpddr_ctrl_axi_s_bvalid ),
				.BRESP( lpddr_ctrl_axi_s_bresp ),
				.BID( lpddr_ctrl_axi_s_bid  ),
				.AWUSER( 32'h0 ),
				.WUSER( 32'h0 ),
				.ARUSER( 32'h0 ),
				.RUSER( 32'h0 ),
				.BUSER( 32'h0 )
				);



