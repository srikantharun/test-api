// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description:
// Owner: abond

`ifndef AXE_DMA_CHANNEL_SEQUENCER_SVH
`define AXE_DMA_CHANNEL_SEQUENCER_SVH

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(uvm_sequence_item) axe_dma_channel_sequencer;


`endif // AXE_DMA_CHANNEL_SEQUENCER_SVH
