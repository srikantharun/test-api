bind ai_core_dwpu_p Axi4PC # (
  .DATA_WIDTH      (ai_core_axi_pkg::AI_CORE_LP_AXI_DATA_WIDTH),
  .ADDR_WIDTH      (ai_core_axi_pkg::AI_CORE_LP_AXI_LOCAL_ADDR_WIDTH),
  .RID_WIDTH       (ai_core_axi_pkg::AI_CORE_LP_AXI_S_ID_WIDTH),
  .WID_WIDTH       (ai_core_axi_pkg::AI_CORE_LP_AXI_S_ID_WIDTH),
  .MAXWBURSTS      (20),
  .MAXRBURSTS      (20),
  .RecommendOn     (0),
  .RecMaxWaitOn    (0),
  .AWREADY_MAXWAITS(256),
  .ARREADY_MAXWAITS(256),
  .WREADY_MAXWAITS (256),
  .BREADY_MAXWAITS (16),
  .RREADY_MAXWAITS (16)
) AXI_AIP_ai_core_dwpu_PROTOCOL_CHECKER (
  .ACLK    (clk),
  .ARESETn (rst_n),
  .ARVALID (ai_core_dwpu_axi_s_arvalid),
  .ARADDR  (ai_core_dwpu_axi_s_araddr),
  .ARLEN   (ai_core_dwpu_axi_s_arlen),
  .ARSIZE  (ai_core_dwpu_axi_s_arsize),
  .ARBURST (ai_core_dwpu_axi_s_arburst),
  .ARLOCK  (ai_core_dwpu_axi_s_arlock),
  .ARCACHE (ai_core_dwpu_axi_s_arcache),
  .ARPROT  (ai_core_dwpu_axi_s_arprot),
  .ARID    (ai_core_dwpu_axi_s_arid),
  .ARREADY (ai_core_dwpu_axi_s_arready),
  .RREADY  (ai_core_dwpu_axi_s_rready),
  .RVALID  (ai_core_dwpu_axi_s_rvalid),
  .RLAST   (ai_core_dwpu_axi_s_rlast),
  .RDATA   (ai_core_dwpu_axi_s_rdata),
  .RRESP   (ai_core_dwpu_axi_s_rresp),
  .RID     (ai_core_dwpu_axi_s_rid),
  .AWVALID (ai_core_dwpu_axi_s_awvalid),
  .AWADDR  (ai_core_dwpu_axi_s_awaddr),
  .AWLEN   (ai_core_dwpu_axi_s_awlen),
  .AWSIZE  (ai_core_dwpu_axi_s_awsize),
  .AWBURST (ai_core_dwpu_axi_s_awburst),
  .AWLOCK  (ai_core_dwpu_axi_s_awlock),
  .AWCACHE (ai_core_dwpu_axi_s_awcache),
  .AWPROT  (ai_core_dwpu_axi_s_awprot),
  .AWID    (ai_core_dwpu_axi_s_awid),
  .AWREADY (ai_core_dwpu_axi_s_awready),
  .WVALID  (ai_core_dwpu_axi_s_wvalid),
  .WLAST   (ai_core_dwpu_axi_s_wlast),
  .WDATA   (ai_core_dwpu_axi_s_wdata),
  .WSTRB   (ai_core_dwpu_axi_s_wstrb),
  .WREADY  (ai_core_dwpu_axi_s_wready),
  .BREADY  (ai_core_dwpu_axi_s_bready),
  .BVALID  (ai_core_dwpu_axi_s_bvalid),
  .BRESP   (ai_core_dwpu_axi_s_bresp),
  .BID     (ai_core_dwpu_axi_s_bid),
  .AWUSER  (32'h0),
  .WUSER   (32'h0),
  .ARUSER  (32'h0),
  .RUSER   (32'h0),
  .BUSER   (32'h0),
  .AWREGION(4'b0),
  .AWQOS   (4'b0),
  .ARQOS   (4'b0),
  .ARREGION(4'b0),
  .CACTIVE (1'b0),
  .CSYSREQ (1'b0),
  .CSYSACK (1'b0)
);
