module ax65_peripheral_wrapper #(
  parameter int unsigned CORE_WIDTH = 6,
  parameter int unsigned ADDR_WIDTH = 40,
  parameter int unsigned DATA_WIDTH = 64,
  parameter int unsigned ID_WIDTH = 8
) (
  input wire i_aclk,
  input wire i_arst_n,
  input wire i_mtime_clk,
  input wire i_por_rst_n,
  output logic [CORE_WIDTH - 1:0] o_cores_mtip,
  input logic [CORE_WIDTH - 1:0] i_cores_stoptime,
  input logic i_test_mode,
  input logic [ADDR_WIDTH-1:0] i_plmt_axi_s_araddr,
  input logic [1:0] i_plmt_axi_s_arburst,
  input logic [3:0] i_plmt_axi_s_arcache,
  input logic [ID_WIDTH-1:0] i_plmt_axi_s_arid,
  input logic [7:0] i_plmt_axi_s_arlen,
  input logic i_plmt_axi_s_arlock,
  input logic [2:0] i_plmt_axi_s_arprot,
  input logic [2:0] i_plmt_axi_s_arsize,
  output logic o_plmt_axi_s_arready,
  input logic i_plmt_axi_s_arvalid,
  input logic [ADDR_WIDTH-1:0] i_plmt_axi_s_awaddr,
  input logic [1:0] i_plmt_axi_s_awburst,
  input logic [3:0] i_plmt_axi_s_awcache,
  input logic [ID_WIDTH-1:0] i_plmt_axi_s_awid,
  input logic [7:0] i_plmt_axi_s_awlen,
  input logic i_plmt_axi_s_awlock,
  input logic [2:0] i_plmt_axi_s_awprot,
  input logic [2:0] i_plmt_axi_s_awsize,
  output logic o_plmt_axi_s_awready,
  input logic i_plmt_axi_s_awvalid,
  output logic [ID_WIDTH-1:0] o_plmt_axi_s_bid,
  output logic [1:0] o_plmt_axi_s_bresp,
  input logic i_plmt_axi_s_bready,
  output logic o_plmt_axi_s_bvalid,
  output logic [DATA_WIDTH-1:0] o_plmt_axi_s_rdata,
  output logic [ID_WIDTH-1:0] o_plmt_axi_s_rid,
  output logic o_plmt_axi_s_rlast,
  output logic [1:0] o_plmt_axi_s_rresp,
  input logic i_plmt_axi_s_rready,
  output logic o_plmt_axi_s_rvalid,
  input logic [DATA_WIDTH-1:0] i_plmt_axi_s_wdata,
  input logic i_plmt_axi_s_wlast,
  input logic [(DATA_WIDTH / 8) - 1:0] i_plmt_axi_s_wstrb,
  output logic o_plmt_axi_s_wready,
  input logic i_plmt_axi_s_wvalid
);

  logic [DATA_WIDTH-1:0] unused_plmt_hrdata;
  logic unused_plmt_hreadyout;
  logic [1:0] unused_plmt_hresp;

  logic stoptime;
  always_comb stoptime = &i_cores_stoptime;

  nceplmt100 #(
    .ADDR_WIDTH(ADDR_WIDTH),
    .BUS_TYPE("axi"),
    .DATA_WIDTH(DATA_WIDTH),
    .GRAY_WIDTH(2),
    .ID_WIDTH(ID_WIDTH),
    .NHART(CORE_WIDTH),
    .SYNC_STAGE(3)
  ) u_plmt (
    .clk(i_aclk),
    .resetn(i_arst_n),
    .mtime_clk(i_mtime_clk),
    .por_rstn(i_por_rst_n),
    .araddr(i_plmt_axi_s_araddr),
    .arburst(i_plmt_axi_s_arburst),
    .arcache(i_plmt_axi_s_arcache),
    .arid(i_plmt_axi_s_arid),
    .arlen(i_plmt_axi_s_arlen),
    .arlock(i_plmt_axi_s_arlock),
    .arprot(i_plmt_axi_s_arprot),
    .arready(o_plmt_axi_s_arready),
    .arsize(i_plmt_axi_s_arsize),
    .arvalid(i_plmt_axi_s_arvalid),
    .awaddr(i_plmt_axi_s_awaddr),
    .awburst(i_plmt_axi_s_awburst),
    .awcache(i_plmt_axi_s_awcache),
    .awid(i_plmt_axi_s_awid),
    .awlen(i_plmt_axi_s_awlen),
    .awlock(i_plmt_axi_s_awlock),
    .awprot(i_plmt_axi_s_awprot),
    .awready(o_plmt_axi_s_awready),
    .awsize(i_plmt_axi_s_awsize),
    .awvalid(i_plmt_axi_s_awvalid),
    .bid(o_plmt_axi_s_bid),
    .bready(i_plmt_axi_s_bready),
    .bresp(o_plmt_axi_s_bresp),
    .bvalid(o_plmt_axi_s_bvalid),
    .haddr({ADDR_WIDTH{1'b0}}),
    .hburst(3'd0),
    .hrdata(unused_plmt_hrdata),
    .hready(1'd0),
    .hreadyout(unused_plmt_hreadyout),
    .hresp(unused_plmt_hresp),
    .hsel(1'd0),
    .hsize(3'd0),
    .htrans(2'd0),
    .hwdata({DATA_WIDTH{1'b0}}),
    .hwrite(1'd0),
    .rdata(o_plmt_axi_s_rdata),
    .rid(o_plmt_axi_s_rid),
    .rlast(o_plmt_axi_s_rlast),
    .rready(i_plmt_axi_s_rready),
    .rresp(o_plmt_axi_s_rresp),
    .rvalid(o_plmt_axi_s_rvalid),
    .wdata(i_plmt_axi_s_wdata),
    .wlast(i_plmt_axi_s_wlast),
    .wready(o_plmt_axi_s_wready),
    .wstrb(i_plmt_axi_s_wstrb),
    .wvalid(i_plmt_axi_s_wvalid),
    .test_mode(i_test_mode),
    .mtip(o_cores_mtip),
    .stoptime(stoptime)
  );

endmodule
