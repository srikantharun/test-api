
// (C) Copyright 2025 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_noc_tok_h_north
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_tok_h_north (
  input wire  i_aic_4_clk,
  input wire  i_aic_4_clken,
  input logic [7:0] i_aic_4_init_tok_ocpl_s_maddr,
  input logic [2:0] i_aic_4_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_4_init_tok_ocpl_s_mdata,
  output logic  o_aic_4_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_4_pwr_tok_idle_val,
  output logic  o_aic_4_pwr_tok_idle_ack,
  input logic  i_aic_4_pwr_tok_idle_req,
  input wire  i_aic_4_rst_n,
  output logic [7:0] o_aic_4_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_aic_4_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_4_targ_tok_ocpl_m_mdata,
  input logic  i_aic_4_targ_tok_ocpl_m_scmdaccept,
  input wire  i_aic_5_clk,
  input wire  i_aic_5_clken,
  input logic [7:0] i_aic_5_init_tok_ocpl_s_maddr,
  input logic [2:0] i_aic_5_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_5_init_tok_ocpl_s_mdata,
  output logic  o_aic_5_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_5_pwr_tok_idle_val,
  output logic  o_aic_5_pwr_tok_idle_ack,
  input logic  i_aic_5_pwr_tok_idle_req,
  input wire  i_aic_5_rst_n,
  output logic [7:0] o_aic_5_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_aic_5_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_5_targ_tok_ocpl_m_mdata,
  input logic  i_aic_5_targ_tok_ocpl_m_scmdaccept,
  input wire  i_aic_6_clk,
  input wire  i_aic_6_clken,
  input logic [7:0] i_aic_6_init_tok_ocpl_s_maddr,
  input logic [2:0] i_aic_6_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_6_init_tok_ocpl_s_mdata,
  output logic  o_aic_6_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_6_pwr_tok_idle_val,
  output logic  o_aic_6_pwr_tok_idle_ack,
  input logic  i_aic_6_pwr_tok_idle_req,
  input wire  i_aic_6_rst_n,
  output logic [7:0] o_aic_6_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_aic_6_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_6_targ_tok_ocpl_m_mdata,
  input logic  i_aic_6_targ_tok_ocpl_m_scmdaccept,
  input wire  i_aic_7_clk,
  input wire  i_aic_7_clken,
  input logic [7:0] i_aic_7_init_tok_ocpl_s_maddr,
  input logic [2:0] i_aic_7_init_tok_ocpl_s_mcmd,
  input logic [7:0] i_aic_7_init_tok_ocpl_s_mdata,
  output logic  o_aic_7_init_tok_ocpl_s_scmdaccept,
  output logic  o_aic_7_pwr_tok_idle_val,
  output logic  o_aic_7_pwr_tok_idle_ack,
  input logic  i_aic_7_pwr_tok_idle_req,
  input wire  i_aic_7_rst_n,
  output logic [7:0] o_aic_7_targ_tok_ocpl_m_maddr,
  output logic [2:0] o_aic_7_targ_tok_ocpl_m_mcmd,
  output logic [7:0] o_aic_7_targ_tok_ocpl_m_mdata,
  input logic  i_aic_7_targ_tok_ocpl_m_scmdaccept,
  input logic [41:0] i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld,
  input wire  i_noc_clk,
  input wire  i_noc_rst_n,
  input logic  scan_en
);

noc_tok_art_h_north u_noc_tok_art_h_north (
  .aic_4_clk(i_aic_4_clk),
  .aic_4_clken(i_aic_4_clken),
  .aic_4_init_tok_MAddr(i_aic_4_init_tok_ocpl_s_maddr),
  .aic_4_init_tok_MCmd(i_aic_4_init_tok_ocpl_s_mcmd),
  .aic_4_init_tok_MData(i_aic_4_init_tok_ocpl_s_mdata),
  .aic_4_init_tok_SCmdAccept(o_aic_4_init_tok_ocpl_s_scmdaccept),
  .aic_4_pwr_tok_Idle(o_aic_4_pwr_tok_idle_val),
  .aic_4_pwr_tok_IdleAck(o_aic_4_pwr_tok_idle_ack),
  .aic_4_pwr_tok_IdleReq(i_aic_4_pwr_tok_idle_req),
  .aic_4_rst_n(i_aic_4_rst_n),
  .aic_4_targ_tok_MAddr(o_aic_4_targ_tok_ocpl_m_maddr),
  .aic_4_targ_tok_MCmd(o_aic_4_targ_tok_ocpl_m_mcmd),
  .aic_4_targ_tok_MData(o_aic_4_targ_tok_ocpl_m_mdata),
  .aic_4_targ_tok_SCmdAccept(i_aic_4_targ_tok_ocpl_m_scmdaccept),
  .aic_5_clk(i_aic_5_clk),
  .aic_5_clken(i_aic_5_clken),
  .aic_5_init_tok_MAddr(i_aic_5_init_tok_ocpl_s_maddr),
  .aic_5_init_tok_MCmd(i_aic_5_init_tok_ocpl_s_mcmd),
  .aic_5_init_tok_MData(i_aic_5_init_tok_ocpl_s_mdata),
  .aic_5_init_tok_SCmdAccept(o_aic_5_init_tok_ocpl_s_scmdaccept),
  .aic_5_pwr_tok_Idle(o_aic_5_pwr_tok_idle_val),
  .aic_5_pwr_tok_IdleAck(o_aic_5_pwr_tok_idle_ack),
  .aic_5_pwr_tok_IdleReq(i_aic_5_pwr_tok_idle_req),
  .aic_5_rst_n(i_aic_5_rst_n),
  .aic_5_targ_tok_MAddr(o_aic_5_targ_tok_ocpl_m_maddr),
  .aic_5_targ_tok_MCmd(o_aic_5_targ_tok_ocpl_m_mcmd),
  .aic_5_targ_tok_MData(o_aic_5_targ_tok_ocpl_m_mdata),
  .aic_5_targ_tok_SCmdAccept(i_aic_5_targ_tok_ocpl_m_scmdaccept),
  .aic_6_clk(i_aic_6_clk),
  .aic_6_clken(i_aic_6_clken),
  .aic_6_init_tok_MAddr(i_aic_6_init_tok_ocpl_s_maddr),
  .aic_6_init_tok_MCmd(i_aic_6_init_tok_ocpl_s_mcmd),
  .aic_6_init_tok_MData(i_aic_6_init_tok_ocpl_s_mdata),
  .aic_6_init_tok_SCmdAccept(o_aic_6_init_tok_ocpl_s_scmdaccept),
  .aic_6_pwr_tok_Idle(o_aic_6_pwr_tok_idle_val),
  .aic_6_pwr_tok_IdleAck(o_aic_6_pwr_tok_idle_ack),
  .aic_6_pwr_tok_IdleReq(i_aic_6_pwr_tok_idle_req),
  .aic_6_rst_n(i_aic_6_rst_n),
  .aic_6_targ_tok_MAddr(o_aic_6_targ_tok_ocpl_m_maddr),
  .aic_6_targ_tok_MCmd(o_aic_6_targ_tok_ocpl_m_mcmd),
  .aic_6_targ_tok_MData(o_aic_6_targ_tok_ocpl_m_mdata),
  .aic_6_targ_tok_SCmdAccept(i_aic_6_targ_tok_ocpl_m_scmdaccept),
  .aic_7_clk(i_aic_7_clk),
  .aic_7_clken(i_aic_7_clken),
  .aic_7_init_tok_MAddr(i_aic_7_init_tok_ocpl_s_maddr),
  .aic_7_init_tok_MCmd(i_aic_7_init_tok_ocpl_s_mcmd),
  .aic_7_init_tok_MData(i_aic_7_init_tok_ocpl_s_mdata),
  .aic_7_init_tok_SCmdAccept(o_aic_7_init_tok_ocpl_s_scmdaccept),
  .aic_7_pwr_tok_Idle(o_aic_7_pwr_tok_idle_val),
  .aic_7_pwr_tok_IdleAck(o_aic_7_pwr_tok_idle_ack),
  .aic_7_pwr_tok_IdleReq(i_aic_7_pwr_tok_idle_req),
  .aic_7_rst_n(i_aic_7_rst_n),
  .aic_7_targ_tok_MAddr(o_aic_7_targ_tok_ocpl_m_maddr),
  .aic_7_targ_tok_MCmd(o_aic_7_targ_tok_ocpl_m_mcmd),
  .aic_7_targ_tok_MData(o_aic_7_targ_tok_ocpl_m_mdata),
  .aic_7_targ_tok_SCmdAccept(i_aic_7_targ_tok_ocpl_m_scmdaccept),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Data(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Head(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Rdy(o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Tail(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail),
  .dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_Vld(i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Data(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Head(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Rdy(o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Tail(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail),
  .dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_Vld(i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Data(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Head(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Rdy(i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Tail(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail),
  .dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_Vld(o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Data(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Head(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Rdy(i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Tail(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail),
  .dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_Vld(o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld),
  .noc_clk(i_noc_clk),
  .noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en)
);
endmodule
