
// (C) Copyright 2025 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_noc_tok_h_east
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_tok_h_east (
  input logic [41:0] i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld,
  input wire  i_noc_clk,
  input wire  i_noc_rst_n,
  input logic  scan_en
);

noc_tok_art_h_east u_noc_tok_art_h_east (
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Data(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data),
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Head(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head),
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Rdy(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy),
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Tail(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail),
  .dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_Vld(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Data(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Head(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Rdy(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Tail(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail),
  .dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_Vld(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Data(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Head(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Rdy(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Tail(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail),
  .dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_Vld(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Data(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Head(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Rdy(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Tail(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail),
  .dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_Vld(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Data(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Head(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Rdy(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Tail(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail),
  .dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_Vld(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Data(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Head(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Rdy(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Tail(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail),
  .dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_Vld(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Data(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Head(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Rdy(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Tail(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail),
  .dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_Vld(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Data(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Head(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Rdy(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Tail(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail),
  .dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_Vld(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld),
  .noc_clk(i_noc_clk),
  .noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en)
);
endmodule
