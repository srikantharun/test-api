// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024


`ifndef __TREK_DELAY_REQ_SV__
`define __TREK_DELAY_REQ_SV__

// User-defined TLM datatype for data in/out of TrekSoC.
//
class trek_delay_req extends uvm_pkg::uvm_transaction;

       bit[63:0]  m_delay = 64'h0000000000000000;

  `uvm_object_utils_begin(trek_delay_req)
    `uvm_field_int(m_delay, UVM_DEFAULT | UVM_HEX)
  `uvm_object_utils_end

  function new(input string name = "trek_delay_req");
    super.new(name);
  endfunction

endclass: trek_delay_req

`endif  // __TREK_DELAY_REQ_SV__
