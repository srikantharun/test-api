// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_ddr_west
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_ddr_west_p (
    input  wire                                        i_ddr_wpll_aon_clk,
    input  wire                                        i_ddr_wpll_aon_rst_n,
    output chip_pkg::chip_syscfg_addr_t                o_ddr_wpll_targ_syscfg_apb_m_paddr,
    output logic                                       o_ddr_wpll_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_ddr_wpll_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_ddr_wpll_targ_syscfg_apb_m_prdata,
    input  logic                                       i_ddr_wpll_targ_syscfg_apb_m_pready,
    output logic                                       o_ddr_wpll_targ_syscfg_apb_m_psel,
    input  logic                                       i_ddr_wpll_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_ddr_wpll_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_ddr_wpll_targ_syscfg_apb_m_pwdata,
    output logic                                       o_ddr_wpll_targ_syscfg_apb_m_pwrite,
    input  logic [398:0]                               i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld,
    output logic [398:0]                               o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld,
    input  logic [398:0]                               i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld,
    output logic [398:0]                               o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld,
    input  logic [398:0]                               i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld,
    output logic [398:0]                               o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld,
    input  logic [398:0]                               i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld,
    output logic [398:0]                               o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld,
    input  logic [146:0]                               i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld,
    output logic [146:0]                               o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head,
    input  logic                                       i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail,
    output logic                                       o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld,
    input  wire                                        i_lpddr_graph_0_aon_clk,
    input  wire                                        i_lpddr_graph_0_aon_rst_n,
    output logic                                       o_lpddr_graph_0_cfg_pwr_idle_val,
    output logic                                       o_lpddr_graph_0_cfg_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_0_cfg_pwr_idle_req,
    input  wire                                        i_lpddr_graph_0_clk,
    input  wire                                        i_lpddr_graph_0_clken,
    output logic                                       o_lpddr_graph_0_pwr_idle_val,
    output logic                                       o_lpddr_graph_0_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_0_pwr_idle_req,
    input  wire                                        i_lpddr_graph_0_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t   o_lpddr_graph_0_targ_cfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_0_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_0_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   i_lpddr_graph_0_targ_cfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_0_targ_cfg_apb_m_pready,
    output logic                                       o_lpddr_graph_0_targ_cfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_0_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                 o_lpddr_graph_0_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   o_lpddr_graph_0_targ_cfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_0_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_0_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_0_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_0_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_0_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_0_targ_ht_axi_m_arlen,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_0_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_0_targ_ht_axi_m_arqos,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_0_targ_ht_axi_m_arsize,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_0_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_0_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_0_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_0_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_0_targ_ht_axi_m_awlen,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_0_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_0_targ_ht_axi_m_awqos,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_0_targ_ht_axi_m_awsize,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_0_targ_ht_axi_m_bid,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_0_targ_ht_axi_m_bresp,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   i_lpddr_graph_0_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_0_targ_ht_axi_m_rid,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_rlast,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_0_targ_ht_axi_m_rresp,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   o_lpddr_graph_0_targ_ht_axi_m_wdata,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_wlast,
    input  logic                                       i_lpddr_graph_0_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t   o_lpddr_graph_0_targ_ht_axi_m_wstrb,
    output logic                                       o_lpddr_graph_0_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                o_lpddr_graph_0_targ_syscfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_lpddr_graph_0_targ_syscfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_0_targ_syscfg_apb_m_pready,
    output logic                                       o_lpddr_graph_0_targ_syscfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_lpddr_graph_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_lpddr_graph_0_targ_syscfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_0_targ_syscfg_apb_m_pwrite,
    input  wire                                        i_lpddr_graph_1_aon_clk,
    input  wire                                        i_lpddr_graph_1_aon_rst_n,
    output logic                                       o_lpddr_graph_1_cfg_pwr_idle_val,
    output logic                                       o_lpddr_graph_1_cfg_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_1_cfg_pwr_idle_req,
    input  wire                                        i_lpddr_graph_1_clk,
    input  wire                                        i_lpddr_graph_1_clken,
    output logic                                       o_lpddr_graph_1_pwr_idle_val,
    output logic                                       o_lpddr_graph_1_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_1_pwr_idle_req,
    input  wire                                        i_lpddr_graph_1_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t   o_lpddr_graph_1_targ_cfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_1_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_1_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   i_lpddr_graph_1_targ_cfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_1_targ_cfg_apb_m_pready,
    output logic                                       o_lpddr_graph_1_targ_cfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_1_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                 o_lpddr_graph_1_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   o_lpddr_graph_1_targ_cfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_1_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_1_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_1_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_1_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_1_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_1_targ_ht_axi_m_arlen,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_1_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_1_targ_ht_axi_m_arqos,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_1_targ_ht_axi_m_arsize,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_1_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_1_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_1_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_1_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_1_targ_ht_axi_m_awlen,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_1_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_1_targ_ht_axi_m_awqos,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_1_targ_ht_axi_m_awsize,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_1_targ_ht_axi_m_bid,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_1_targ_ht_axi_m_bresp,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   i_lpddr_graph_1_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_1_targ_ht_axi_m_rid,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_rlast,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_1_targ_ht_axi_m_rresp,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   o_lpddr_graph_1_targ_ht_axi_m_wdata,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_wlast,
    input  logic                                       i_lpddr_graph_1_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t   o_lpddr_graph_1_targ_ht_axi_m_wstrb,
    output logic                                       o_lpddr_graph_1_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                o_lpddr_graph_1_targ_syscfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_lpddr_graph_1_targ_syscfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_1_targ_syscfg_apb_m_pready,
    output logic                                       o_lpddr_graph_1_targ_syscfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_lpddr_graph_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_lpddr_graph_1_targ_syscfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_1_targ_syscfg_apb_m_pwrite,
    input  wire                                        i_lpddr_graph_2_aon_clk,
    input  wire                                        i_lpddr_graph_2_aon_rst_n,
    output logic                                       o_lpddr_graph_2_cfg_pwr_idle_val,
    output logic                                       o_lpddr_graph_2_cfg_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_2_cfg_pwr_idle_req,
    input  wire                                        i_lpddr_graph_2_clk,
    input  wire                                        i_lpddr_graph_2_clken,
    output logic                                       o_lpddr_graph_2_pwr_idle_val,
    output logic                                       o_lpddr_graph_2_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_2_pwr_idle_req,
    input  wire                                        i_lpddr_graph_2_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t   o_lpddr_graph_2_targ_cfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_2_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_2_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   i_lpddr_graph_2_targ_cfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_2_targ_cfg_apb_m_pready,
    output logic                                       o_lpddr_graph_2_targ_cfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_2_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                 o_lpddr_graph_2_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   o_lpddr_graph_2_targ_cfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_2_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_2_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_2_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_2_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_2_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_2_targ_ht_axi_m_arlen,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_2_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_2_targ_ht_axi_m_arqos,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_2_targ_ht_axi_m_arsize,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_2_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_2_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_2_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_2_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_2_targ_ht_axi_m_awlen,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_2_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_2_targ_ht_axi_m_awqos,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_2_targ_ht_axi_m_awsize,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_2_targ_ht_axi_m_bid,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_2_targ_ht_axi_m_bresp,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   i_lpddr_graph_2_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_2_targ_ht_axi_m_rid,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_rlast,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_2_targ_ht_axi_m_rresp,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   o_lpddr_graph_2_targ_ht_axi_m_wdata,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_wlast,
    input  logic                                       i_lpddr_graph_2_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t   o_lpddr_graph_2_targ_ht_axi_m_wstrb,
    output logic                                       o_lpddr_graph_2_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                o_lpddr_graph_2_targ_syscfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_lpddr_graph_2_targ_syscfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_2_targ_syscfg_apb_m_pready,
    output logic                                       o_lpddr_graph_2_targ_syscfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_lpddr_graph_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_lpddr_graph_2_targ_syscfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_2_targ_syscfg_apb_m_pwrite,
    input  wire                                        i_lpddr_graph_3_aon_clk,
    input  wire                                        i_lpddr_graph_3_aon_rst_n,
    output logic                                       o_lpddr_graph_3_cfg_pwr_idle_val,
    output logic                                       o_lpddr_graph_3_cfg_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_3_cfg_pwr_idle_req,
    input  wire                                        i_lpddr_graph_3_clk,
    input  wire                                        i_lpddr_graph_3_clken,
    output logic                                       o_lpddr_graph_3_pwr_idle_val,
    output logic                                       o_lpddr_graph_3_pwr_idle_ack,
    input  logic                                       i_lpddr_graph_3_pwr_idle_req,
    input  wire                                        i_lpddr_graph_3_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t   o_lpddr_graph_3_targ_cfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_3_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_3_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   i_lpddr_graph_3_targ_cfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_3_targ_cfg_apb_m_pready,
    output logic                                       o_lpddr_graph_3_targ_cfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_3_targ_cfg_apb_m_pslverr,
    output logic [3:0]                                 o_lpddr_graph_3_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t   o_lpddr_graph_3_targ_cfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_3_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_3_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_3_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_3_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_3_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_3_targ_ht_axi_m_arlen,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_3_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_3_targ_ht_axi_m_arqos,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_3_targ_ht_axi_m_arsize,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                   o_lpddr_graph_3_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                        o_lpddr_graph_3_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                        o_lpddr_graph_3_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     o_lpddr_graph_3_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                          o_lpddr_graph_3_targ_ht_axi_m_awlen,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                         o_lpddr_graph_3_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                          o_lpddr_graph_3_targ_ht_axi_m_awqos,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                         o_lpddr_graph_3_targ_ht_axi_m_awsize,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_3_targ_ht_axi_m_bid,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_3_targ_ht_axi_m_bresp,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   i_lpddr_graph_3_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t     i_lpddr_graph_3_targ_ht_axi_m_rid,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_rlast,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                         i_lpddr_graph_3_targ_ht_axi_m_rresp,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t   o_lpddr_graph_3_targ_ht_axi_m_wdata,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_wlast,
    input  logic                                       i_lpddr_graph_3_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t   o_lpddr_graph_3_targ_ht_axi_m_wstrb,
    output logic                                       o_lpddr_graph_3_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                o_lpddr_graph_3_targ_syscfg_apb_m_paddr,
    output logic                                       o_lpddr_graph_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                     o_lpddr_graph_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t            i_lpddr_graph_3_targ_syscfg_apb_m_prdata,
    input  logic                                       i_lpddr_graph_3_targ_syscfg_apb_m_pready,
    output logic                                       o_lpddr_graph_3_targ_syscfg_apb_m_psel,
    input  logic                                       i_lpddr_graph_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t            o_lpddr_graph_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t            o_lpddr_graph_3_targ_syscfg_apb_m_pwdata,
    output logic                                       o_lpddr_graph_3_targ_syscfg_apb_m_pwrite,
    input  wire                                        i_noc_clk,
    input  wire                                        i_noc_rst_n,
    // DFT Interface
    input  wire           tck,
    input  wire           trst,
    input  logic          tms,
    input  logic          tdi,
    output logic          tdo_en,
    output logic          tdo,
    input  wire           test_clk,
    input  logic          test_mode,
    input  logic          edt_update,
    input  logic          scan_en,
    input  logic [12-1:0] scan_in,
    output logic [12-1:0] scan_out
);
    // -- Automatically-generated Reset Synchronizers -- //
    wire lpddr_graph_0_aon_rst_n_synced;
    wire lpddr_graph_1_aon_rst_n_synced;
    wire lpddr_graph_2_aon_rst_n_synced;
    wire lpddr_graph_3_aon_rst_n_synced;
    wire ddr_wpll_aon_rst_n_synced;

    // LPDDR GRAPH 0 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_lpddr_graph_0_aon_rst_n_sync (
        .i_clk          (i_lpddr_graph_0_aon_clk),
        .i_rst_n        (i_lpddr_graph_0_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (lpddr_graph_0_aon_rst_n_synced)
    );

    // LPDDR GRAPH 1 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_lpddr_graph_1_aon_rst_n_sync (
        .i_clk          (i_lpddr_graph_1_aon_clk),
        .i_rst_n        (i_lpddr_graph_1_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (lpddr_graph_1_aon_rst_n_synced)
    );

    // LPDDR GRAPH 2 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_lpddr_graph_2_aon_rst_n_sync (
        .i_clk          (i_lpddr_graph_2_aon_clk),
        .i_rst_n        (i_lpddr_graph_2_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (lpddr_graph_2_aon_rst_n_synced)
    );

    // LPDDR GRAPH 3 AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_lpddr_graph_3_aon_rst_n_sync (
        .i_clk          (i_lpddr_graph_3_aon_clk),
        .i_rst_n        (i_lpddr_graph_3_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (lpddr_graph_3_aon_rst_n_synced)
    );

    // DDR WPLL AON Reset Synchronizer
    axe_ccl_rst_n_sync #(
        .SyncStages (2)
    ) u_ddr_wpll_aon_rst_n_sync (
        .i_clk          (i_ddr_wpll_aon_clk),
        .i_rst_n        (i_ddr_wpll_aon_rst_n),
        .i_test_mode    (test_mode),
        .o_rst_n        (ddr_wpll_aon_rst_n_synced)
    );

    noc_ddr_west u_noc_ddr_west (
    .i_ddr_wpll_aon_clk(i_ddr_wpll_aon_clk),
    .i_ddr_wpll_aon_rst_n(ddr_wpll_aon_rst_n_synced),
    .o_ddr_wpll_targ_syscfg_apb_m_paddr(o_ddr_wpll_targ_syscfg_apb_m_paddr),
    .o_ddr_wpll_targ_syscfg_apb_m_penable(o_ddr_wpll_targ_syscfg_apb_m_penable),
    .o_ddr_wpll_targ_syscfg_apb_m_pprot(o_ddr_wpll_targ_syscfg_apb_m_pprot),
    .i_ddr_wpll_targ_syscfg_apb_m_prdata(i_ddr_wpll_targ_syscfg_apb_m_prdata),
    .i_ddr_wpll_targ_syscfg_apb_m_pready(i_ddr_wpll_targ_syscfg_apb_m_pready),
    .o_ddr_wpll_targ_syscfg_apb_m_psel(o_ddr_wpll_targ_syscfg_apb_m_psel),
    .i_ddr_wpll_targ_syscfg_apb_m_pslverr(i_ddr_wpll_targ_syscfg_apb_m_pslverr),
    .o_ddr_wpll_targ_syscfg_apb_m_pstrb(o_ddr_wpll_targ_syscfg_apb_m_pstrb),
    .o_ddr_wpll_targ_syscfg_apb_m_pwdata(o_ddr_wpll_targ_syscfg_apb_m_pwdata),
    .o_ddr_wpll_targ_syscfg_apb_m_pwrite(o_ddr_wpll_targ_syscfg_apb_m_pwrite),
    .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data),
    .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head),
    .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy(o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy),
    .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail),
    .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld(i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld),
    .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data),
    .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head),
    .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy(i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy),
    .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail),
    .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld(o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld),
    .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data),
    .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head),
    .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy(o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy),
    .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail),
    .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld(i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld),
    .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data),
    .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head),
    .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy(i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy),
    .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail),
    .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld(o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld),
    .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data),
    .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head),
    .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy(o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy),
    .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail),
    .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld(i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld),
    .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data),
    .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head),
    .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy(i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy),
    .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail),
    .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld(o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld),
    .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data),
    .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head),
    .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy(o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy),
    .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail),
    .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld(i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld),
    .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data),
    .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head),
    .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy(i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy),
    .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail),
    .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld(o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld),
    .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data),
    .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head),
    .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy(o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy),
    .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail),
    .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld(i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld),
    .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data),
    .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head),
    .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy(i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy),
    .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail),
    .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld(o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld),
    .i_lpddr_graph_0_aon_clk(i_lpddr_graph_0_aon_clk),
    .i_lpddr_graph_0_aon_rst_n(lpddr_graph_0_aon_rst_n_synced),
    .o_lpddr_graph_0_cfg_pwr_idle_val(o_lpddr_graph_0_cfg_pwr_idle_val),
    .o_lpddr_graph_0_cfg_pwr_idle_ack(o_lpddr_graph_0_cfg_pwr_idle_ack),
    .i_lpddr_graph_0_cfg_pwr_idle_req(i_lpddr_graph_0_cfg_pwr_idle_req),
    .i_lpddr_graph_0_clk(i_lpddr_graph_0_clk),
    .i_lpddr_graph_0_clken(i_lpddr_graph_0_clken),
    .o_lpddr_graph_0_pwr_idle_val(o_lpddr_graph_0_pwr_idle_val),
    .o_lpddr_graph_0_pwr_idle_ack(o_lpddr_graph_0_pwr_idle_ack),
    .i_lpddr_graph_0_pwr_idle_req(i_lpddr_graph_0_pwr_idle_req),
    .i_lpddr_graph_0_rst_n(i_lpddr_graph_0_rst_n),
    .o_lpddr_graph_0_targ_cfg_apb_m_paddr(o_lpddr_graph_0_targ_cfg_apb_m_paddr),
    .o_lpddr_graph_0_targ_cfg_apb_m_penable(o_lpddr_graph_0_targ_cfg_apb_m_penable),
    .o_lpddr_graph_0_targ_cfg_apb_m_pprot(o_lpddr_graph_0_targ_cfg_apb_m_pprot),
    .i_lpddr_graph_0_targ_cfg_apb_m_prdata(i_lpddr_graph_0_targ_cfg_apb_m_prdata),
    .i_lpddr_graph_0_targ_cfg_apb_m_pready(i_lpddr_graph_0_targ_cfg_apb_m_pready),
    .o_lpddr_graph_0_targ_cfg_apb_m_psel(o_lpddr_graph_0_targ_cfg_apb_m_psel),
    .i_lpddr_graph_0_targ_cfg_apb_m_pslverr(i_lpddr_graph_0_targ_cfg_apb_m_pslverr),
    .o_lpddr_graph_0_targ_cfg_apb_m_pstrb(o_lpddr_graph_0_targ_cfg_apb_m_pstrb),
    .o_lpddr_graph_0_targ_cfg_apb_m_pwdata(o_lpddr_graph_0_targ_cfg_apb_m_pwdata),
    .o_lpddr_graph_0_targ_cfg_apb_m_pwrite(o_lpddr_graph_0_targ_cfg_apb_m_pwrite),
    .o_lpddr_graph_0_targ_ht_axi_m_araddr(o_lpddr_graph_0_targ_ht_axi_m_araddr),
    .o_lpddr_graph_0_targ_ht_axi_m_arburst(o_lpddr_graph_0_targ_ht_axi_m_arburst),
    .o_lpddr_graph_0_targ_ht_axi_m_arcache(o_lpddr_graph_0_targ_ht_axi_m_arcache),
    .o_lpddr_graph_0_targ_ht_axi_m_arid(o_lpddr_graph_0_targ_ht_axi_m_arid),
    .o_lpddr_graph_0_targ_ht_axi_m_arlen(o_lpddr_graph_0_targ_ht_axi_m_arlen),
    .o_lpddr_graph_0_targ_ht_axi_m_arlock(o_lpddr_graph_0_targ_ht_axi_m_arlock),
    .o_lpddr_graph_0_targ_ht_axi_m_arprot(o_lpddr_graph_0_targ_ht_axi_m_arprot),
    .o_lpddr_graph_0_targ_ht_axi_m_arqos(o_lpddr_graph_0_targ_ht_axi_m_arqos),
    .i_lpddr_graph_0_targ_ht_axi_m_arready(i_lpddr_graph_0_targ_ht_axi_m_arready),
    .o_lpddr_graph_0_targ_ht_axi_m_arsize(o_lpddr_graph_0_targ_ht_axi_m_arsize),
    .o_lpddr_graph_0_targ_ht_axi_m_arvalid(o_lpddr_graph_0_targ_ht_axi_m_arvalid),
    .o_lpddr_graph_0_targ_ht_axi_m_awaddr(o_lpddr_graph_0_targ_ht_axi_m_awaddr),
    .o_lpddr_graph_0_targ_ht_axi_m_awburst(o_lpddr_graph_0_targ_ht_axi_m_awburst),
    .o_lpddr_graph_0_targ_ht_axi_m_awcache(o_lpddr_graph_0_targ_ht_axi_m_awcache),
    .o_lpddr_graph_0_targ_ht_axi_m_awid(o_lpddr_graph_0_targ_ht_axi_m_awid),
    .o_lpddr_graph_0_targ_ht_axi_m_awlen(o_lpddr_graph_0_targ_ht_axi_m_awlen),
    .o_lpddr_graph_0_targ_ht_axi_m_awlock(o_lpddr_graph_0_targ_ht_axi_m_awlock),
    .o_lpddr_graph_0_targ_ht_axi_m_awprot(o_lpddr_graph_0_targ_ht_axi_m_awprot),
    .o_lpddr_graph_0_targ_ht_axi_m_awqos(o_lpddr_graph_0_targ_ht_axi_m_awqos),
    .i_lpddr_graph_0_targ_ht_axi_m_awready(i_lpddr_graph_0_targ_ht_axi_m_awready),
    .o_lpddr_graph_0_targ_ht_axi_m_awsize(o_lpddr_graph_0_targ_ht_axi_m_awsize),
    .o_lpddr_graph_0_targ_ht_axi_m_awvalid(o_lpddr_graph_0_targ_ht_axi_m_awvalid),
    .i_lpddr_graph_0_targ_ht_axi_m_bid(i_lpddr_graph_0_targ_ht_axi_m_bid),
    .o_lpddr_graph_0_targ_ht_axi_m_bready(o_lpddr_graph_0_targ_ht_axi_m_bready),
    .i_lpddr_graph_0_targ_ht_axi_m_bresp(i_lpddr_graph_0_targ_ht_axi_m_bresp),
    .i_lpddr_graph_0_targ_ht_axi_m_bvalid(i_lpddr_graph_0_targ_ht_axi_m_bvalid),
    .i_lpddr_graph_0_targ_ht_axi_m_rdata(i_lpddr_graph_0_targ_ht_axi_m_rdata),
    .i_lpddr_graph_0_targ_ht_axi_m_rid(i_lpddr_graph_0_targ_ht_axi_m_rid),
    .i_lpddr_graph_0_targ_ht_axi_m_rlast(i_lpddr_graph_0_targ_ht_axi_m_rlast),
    .o_lpddr_graph_0_targ_ht_axi_m_rready(o_lpddr_graph_0_targ_ht_axi_m_rready),
    .i_lpddr_graph_0_targ_ht_axi_m_rresp(i_lpddr_graph_0_targ_ht_axi_m_rresp),
    .i_lpddr_graph_0_targ_ht_axi_m_rvalid(i_lpddr_graph_0_targ_ht_axi_m_rvalid),
    .o_lpddr_graph_0_targ_ht_axi_m_wdata(o_lpddr_graph_0_targ_ht_axi_m_wdata),
    .o_lpddr_graph_0_targ_ht_axi_m_wlast(o_lpddr_graph_0_targ_ht_axi_m_wlast),
    .i_lpddr_graph_0_targ_ht_axi_m_wready(i_lpddr_graph_0_targ_ht_axi_m_wready),
    .o_lpddr_graph_0_targ_ht_axi_m_wstrb(o_lpddr_graph_0_targ_ht_axi_m_wstrb),
    .o_lpddr_graph_0_targ_ht_axi_m_wvalid(o_lpddr_graph_0_targ_ht_axi_m_wvalid),
    .o_lpddr_graph_0_targ_syscfg_apb_m_paddr(o_lpddr_graph_0_targ_syscfg_apb_m_paddr),
    .o_lpddr_graph_0_targ_syscfg_apb_m_penable(o_lpddr_graph_0_targ_syscfg_apb_m_penable),
    .o_lpddr_graph_0_targ_syscfg_apb_m_pprot(o_lpddr_graph_0_targ_syscfg_apb_m_pprot),
    .i_lpddr_graph_0_targ_syscfg_apb_m_prdata(i_lpddr_graph_0_targ_syscfg_apb_m_prdata),
    .i_lpddr_graph_0_targ_syscfg_apb_m_pready(i_lpddr_graph_0_targ_syscfg_apb_m_pready),
    .o_lpddr_graph_0_targ_syscfg_apb_m_psel(o_lpddr_graph_0_targ_syscfg_apb_m_psel),
    .i_lpddr_graph_0_targ_syscfg_apb_m_pslverr(i_lpddr_graph_0_targ_syscfg_apb_m_pslverr),
    .o_lpddr_graph_0_targ_syscfg_apb_m_pstrb(o_lpddr_graph_0_targ_syscfg_apb_m_pstrb),
    .o_lpddr_graph_0_targ_syscfg_apb_m_pwdata(o_lpddr_graph_0_targ_syscfg_apb_m_pwdata),
    .o_lpddr_graph_0_targ_syscfg_apb_m_pwrite(o_lpddr_graph_0_targ_syscfg_apb_m_pwrite),
    .i_lpddr_graph_1_aon_clk(i_lpddr_graph_1_aon_clk),
    .i_lpddr_graph_1_aon_rst_n(lpddr_graph_1_aon_rst_n_synced),
    .o_lpddr_graph_1_cfg_pwr_idle_val(o_lpddr_graph_1_cfg_pwr_idle_val),
    .o_lpddr_graph_1_cfg_pwr_idle_ack(o_lpddr_graph_1_cfg_pwr_idle_ack),
    .i_lpddr_graph_1_cfg_pwr_idle_req(i_lpddr_graph_1_cfg_pwr_idle_req),
    .i_lpddr_graph_1_clk(i_lpddr_graph_1_clk),
    .i_lpddr_graph_1_clken(i_lpddr_graph_1_clken),
    .o_lpddr_graph_1_pwr_idle_val(o_lpddr_graph_1_pwr_idle_val),
    .o_lpddr_graph_1_pwr_idle_ack(o_lpddr_graph_1_pwr_idle_ack),
    .i_lpddr_graph_1_pwr_idle_req(i_lpddr_graph_1_pwr_idle_req),
    .i_lpddr_graph_1_rst_n(i_lpddr_graph_1_rst_n),
    .o_lpddr_graph_1_targ_cfg_apb_m_paddr(o_lpddr_graph_1_targ_cfg_apb_m_paddr),
    .o_lpddr_graph_1_targ_cfg_apb_m_penable(o_lpddr_graph_1_targ_cfg_apb_m_penable),
    .o_lpddr_graph_1_targ_cfg_apb_m_pprot(o_lpddr_graph_1_targ_cfg_apb_m_pprot),
    .i_lpddr_graph_1_targ_cfg_apb_m_prdata(i_lpddr_graph_1_targ_cfg_apb_m_prdata),
    .i_lpddr_graph_1_targ_cfg_apb_m_pready(i_lpddr_graph_1_targ_cfg_apb_m_pready),
    .o_lpddr_graph_1_targ_cfg_apb_m_psel(o_lpddr_graph_1_targ_cfg_apb_m_psel),
    .i_lpddr_graph_1_targ_cfg_apb_m_pslverr(i_lpddr_graph_1_targ_cfg_apb_m_pslverr),
    .o_lpddr_graph_1_targ_cfg_apb_m_pstrb(o_lpddr_graph_1_targ_cfg_apb_m_pstrb),
    .o_lpddr_graph_1_targ_cfg_apb_m_pwdata(o_lpddr_graph_1_targ_cfg_apb_m_pwdata),
    .o_lpddr_graph_1_targ_cfg_apb_m_pwrite(o_lpddr_graph_1_targ_cfg_apb_m_pwrite),
    .o_lpddr_graph_1_targ_ht_axi_m_araddr(o_lpddr_graph_1_targ_ht_axi_m_araddr),
    .o_lpddr_graph_1_targ_ht_axi_m_arburst(o_lpddr_graph_1_targ_ht_axi_m_arburst),
    .o_lpddr_graph_1_targ_ht_axi_m_arcache(o_lpddr_graph_1_targ_ht_axi_m_arcache),
    .o_lpddr_graph_1_targ_ht_axi_m_arid(o_lpddr_graph_1_targ_ht_axi_m_arid),
    .o_lpddr_graph_1_targ_ht_axi_m_arlen(o_lpddr_graph_1_targ_ht_axi_m_arlen),
    .o_lpddr_graph_1_targ_ht_axi_m_arlock(o_lpddr_graph_1_targ_ht_axi_m_arlock),
    .o_lpddr_graph_1_targ_ht_axi_m_arprot(o_lpddr_graph_1_targ_ht_axi_m_arprot),
    .o_lpddr_graph_1_targ_ht_axi_m_arqos(o_lpddr_graph_1_targ_ht_axi_m_arqos),
    .i_lpddr_graph_1_targ_ht_axi_m_arready(i_lpddr_graph_1_targ_ht_axi_m_arready),
    .o_lpddr_graph_1_targ_ht_axi_m_arsize(o_lpddr_graph_1_targ_ht_axi_m_arsize),
    .o_lpddr_graph_1_targ_ht_axi_m_arvalid(o_lpddr_graph_1_targ_ht_axi_m_arvalid),
    .o_lpddr_graph_1_targ_ht_axi_m_awaddr(o_lpddr_graph_1_targ_ht_axi_m_awaddr),
    .o_lpddr_graph_1_targ_ht_axi_m_awburst(o_lpddr_graph_1_targ_ht_axi_m_awburst),
    .o_lpddr_graph_1_targ_ht_axi_m_awcache(o_lpddr_graph_1_targ_ht_axi_m_awcache),
    .o_lpddr_graph_1_targ_ht_axi_m_awid(o_lpddr_graph_1_targ_ht_axi_m_awid),
    .o_lpddr_graph_1_targ_ht_axi_m_awlen(o_lpddr_graph_1_targ_ht_axi_m_awlen),
    .o_lpddr_graph_1_targ_ht_axi_m_awlock(o_lpddr_graph_1_targ_ht_axi_m_awlock),
    .o_lpddr_graph_1_targ_ht_axi_m_awprot(o_lpddr_graph_1_targ_ht_axi_m_awprot),
    .o_lpddr_graph_1_targ_ht_axi_m_awqos(o_lpddr_graph_1_targ_ht_axi_m_awqos),
    .i_lpddr_graph_1_targ_ht_axi_m_awready(i_lpddr_graph_1_targ_ht_axi_m_awready),
    .o_lpddr_graph_1_targ_ht_axi_m_awsize(o_lpddr_graph_1_targ_ht_axi_m_awsize),
    .o_lpddr_graph_1_targ_ht_axi_m_awvalid(o_lpddr_graph_1_targ_ht_axi_m_awvalid),
    .i_lpddr_graph_1_targ_ht_axi_m_bid(i_lpddr_graph_1_targ_ht_axi_m_bid),
    .o_lpddr_graph_1_targ_ht_axi_m_bready(o_lpddr_graph_1_targ_ht_axi_m_bready),
    .i_lpddr_graph_1_targ_ht_axi_m_bresp(i_lpddr_graph_1_targ_ht_axi_m_bresp),
    .i_lpddr_graph_1_targ_ht_axi_m_bvalid(i_lpddr_graph_1_targ_ht_axi_m_bvalid),
    .i_lpddr_graph_1_targ_ht_axi_m_rdata(i_lpddr_graph_1_targ_ht_axi_m_rdata),
    .i_lpddr_graph_1_targ_ht_axi_m_rid(i_lpddr_graph_1_targ_ht_axi_m_rid),
    .i_lpddr_graph_1_targ_ht_axi_m_rlast(i_lpddr_graph_1_targ_ht_axi_m_rlast),
    .o_lpddr_graph_1_targ_ht_axi_m_rready(o_lpddr_graph_1_targ_ht_axi_m_rready),
    .i_lpddr_graph_1_targ_ht_axi_m_rresp(i_lpddr_graph_1_targ_ht_axi_m_rresp),
    .i_lpddr_graph_1_targ_ht_axi_m_rvalid(i_lpddr_graph_1_targ_ht_axi_m_rvalid),
    .o_lpddr_graph_1_targ_ht_axi_m_wdata(o_lpddr_graph_1_targ_ht_axi_m_wdata),
    .o_lpddr_graph_1_targ_ht_axi_m_wlast(o_lpddr_graph_1_targ_ht_axi_m_wlast),
    .i_lpddr_graph_1_targ_ht_axi_m_wready(i_lpddr_graph_1_targ_ht_axi_m_wready),
    .o_lpddr_graph_1_targ_ht_axi_m_wstrb(o_lpddr_graph_1_targ_ht_axi_m_wstrb),
    .o_lpddr_graph_1_targ_ht_axi_m_wvalid(o_lpddr_graph_1_targ_ht_axi_m_wvalid),
    .o_lpddr_graph_1_targ_syscfg_apb_m_paddr(o_lpddr_graph_1_targ_syscfg_apb_m_paddr),
    .o_lpddr_graph_1_targ_syscfg_apb_m_penable(o_lpddr_graph_1_targ_syscfg_apb_m_penable),
    .o_lpddr_graph_1_targ_syscfg_apb_m_pprot(o_lpddr_graph_1_targ_syscfg_apb_m_pprot),
    .i_lpddr_graph_1_targ_syscfg_apb_m_prdata(i_lpddr_graph_1_targ_syscfg_apb_m_prdata),
    .i_lpddr_graph_1_targ_syscfg_apb_m_pready(i_lpddr_graph_1_targ_syscfg_apb_m_pready),
    .o_lpddr_graph_1_targ_syscfg_apb_m_psel(o_lpddr_graph_1_targ_syscfg_apb_m_psel),
    .i_lpddr_graph_1_targ_syscfg_apb_m_pslverr(i_lpddr_graph_1_targ_syscfg_apb_m_pslverr),
    .o_lpddr_graph_1_targ_syscfg_apb_m_pstrb(o_lpddr_graph_1_targ_syscfg_apb_m_pstrb),
    .o_lpddr_graph_1_targ_syscfg_apb_m_pwdata(o_lpddr_graph_1_targ_syscfg_apb_m_pwdata),
    .o_lpddr_graph_1_targ_syscfg_apb_m_pwrite(o_lpddr_graph_1_targ_syscfg_apb_m_pwrite),
    .i_lpddr_graph_2_aon_clk(i_lpddr_graph_2_aon_clk),
    .i_lpddr_graph_2_aon_rst_n(lpddr_graph_2_aon_rst_n_synced),
    .o_lpddr_graph_2_cfg_pwr_idle_val(o_lpddr_graph_2_cfg_pwr_idle_val),
    .o_lpddr_graph_2_cfg_pwr_idle_ack(o_lpddr_graph_2_cfg_pwr_idle_ack),
    .i_lpddr_graph_2_cfg_pwr_idle_req(i_lpddr_graph_2_cfg_pwr_idle_req),
    .i_lpddr_graph_2_clk(i_lpddr_graph_2_clk),
    .i_lpddr_graph_2_clken(i_lpddr_graph_2_clken),
    .o_lpddr_graph_2_pwr_idle_val(o_lpddr_graph_2_pwr_idle_val),
    .o_lpddr_graph_2_pwr_idle_ack(o_lpddr_graph_2_pwr_idle_ack),
    .i_lpddr_graph_2_pwr_idle_req(i_lpddr_graph_2_pwr_idle_req),
    .i_lpddr_graph_2_rst_n(i_lpddr_graph_2_rst_n),
    .o_lpddr_graph_2_targ_cfg_apb_m_paddr(o_lpddr_graph_2_targ_cfg_apb_m_paddr),
    .o_lpddr_graph_2_targ_cfg_apb_m_penable(o_lpddr_graph_2_targ_cfg_apb_m_penable),
    .o_lpddr_graph_2_targ_cfg_apb_m_pprot(o_lpddr_graph_2_targ_cfg_apb_m_pprot),
    .i_lpddr_graph_2_targ_cfg_apb_m_prdata(i_lpddr_graph_2_targ_cfg_apb_m_prdata),
    .i_lpddr_graph_2_targ_cfg_apb_m_pready(i_lpddr_graph_2_targ_cfg_apb_m_pready),
    .o_lpddr_graph_2_targ_cfg_apb_m_psel(o_lpddr_graph_2_targ_cfg_apb_m_psel),
    .i_lpddr_graph_2_targ_cfg_apb_m_pslverr(i_lpddr_graph_2_targ_cfg_apb_m_pslverr),
    .o_lpddr_graph_2_targ_cfg_apb_m_pstrb(o_lpddr_graph_2_targ_cfg_apb_m_pstrb),
    .o_lpddr_graph_2_targ_cfg_apb_m_pwdata(o_lpddr_graph_2_targ_cfg_apb_m_pwdata),
    .o_lpddr_graph_2_targ_cfg_apb_m_pwrite(o_lpddr_graph_2_targ_cfg_apb_m_pwrite),
    .o_lpddr_graph_2_targ_ht_axi_m_araddr(o_lpddr_graph_2_targ_ht_axi_m_araddr),
    .o_lpddr_graph_2_targ_ht_axi_m_arburst(o_lpddr_graph_2_targ_ht_axi_m_arburst),
    .o_lpddr_graph_2_targ_ht_axi_m_arcache(o_lpddr_graph_2_targ_ht_axi_m_arcache),
    .o_lpddr_graph_2_targ_ht_axi_m_arid(o_lpddr_graph_2_targ_ht_axi_m_arid),
    .o_lpddr_graph_2_targ_ht_axi_m_arlen(o_lpddr_graph_2_targ_ht_axi_m_arlen),
    .o_lpddr_graph_2_targ_ht_axi_m_arlock(o_lpddr_graph_2_targ_ht_axi_m_arlock),
    .o_lpddr_graph_2_targ_ht_axi_m_arprot(o_lpddr_graph_2_targ_ht_axi_m_arprot),
    .o_lpddr_graph_2_targ_ht_axi_m_arqos(o_lpddr_graph_2_targ_ht_axi_m_arqos),
    .i_lpddr_graph_2_targ_ht_axi_m_arready(i_lpddr_graph_2_targ_ht_axi_m_arready),
    .o_lpddr_graph_2_targ_ht_axi_m_arsize(o_lpddr_graph_2_targ_ht_axi_m_arsize),
    .o_lpddr_graph_2_targ_ht_axi_m_arvalid(o_lpddr_graph_2_targ_ht_axi_m_arvalid),
    .o_lpddr_graph_2_targ_ht_axi_m_awaddr(o_lpddr_graph_2_targ_ht_axi_m_awaddr),
    .o_lpddr_graph_2_targ_ht_axi_m_awburst(o_lpddr_graph_2_targ_ht_axi_m_awburst),
    .o_lpddr_graph_2_targ_ht_axi_m_awcache(o_lpddr_graph_2_targ_ht_axi_m_awcache),
    .o_lpddr_graph_2_targ_ht_axi_m_awid(o_lpddr_graph_2_targ_ht_axi_m_awid),
    .o_lpddr_graph_2_targ_ht_axi_m_awlen(o_lpddr_graph_2_targ_ht_axi_m_awlen),
    .o_lpddr_graph_2_targ_ht_axi_m_awlock(o_lpddr_graph_2_targ_ht_axi_m_awlock),
    .o_lpddr_graph_2_targ_ht_axi_m_awprot(o_lpddr_graph_2_targ_ht_axi_m_awprot),
    .o_lpddr_graph_2_targ_ht_axi_m_awqos(o_lpddr_graph_2_targ_ht_axi_m_awqos),
    .i_lpddr_graph_2_targ_ht_axi_m_awready(i_lpddr_graph_2_targ_ht_axi_m_awready),
    .o_lpddr_graph_2_targ_ht_axi_m_awsize(o_lpddr_graph_2_targ_ht_axi_m_awsize),
    .o_lpddr_graph_2_targ_ht_axi_m_awvalid(o_lpddr_graph_2_targ_ht_axi_m_awvalid),
    .i_lpddr_graph_2_targ_ht_axi_m_bid(i_lpddr_graph_2_targ_ht_axi_m_bid),
    .o_lpddr_graph_2_targ_ht_axi_m_bready(o_lpddr_graph_2_targ_ht_axi_m_bready),
    .i_lpddr_graph_2_targ_ht_axi_m_bresp(i_lpddr_graph_2_targ_ht_axi_m_bresp),
    .i_lpddr_graph_2_targ_ht_axi_m_bvalid(i_lpddr_graph_2_targ_ht_axi_m_bvalid),
    .i_lpddr_graph_2_targ_ht_axi_m_rdata(i_lpddr_graph_2_targ_ht_axi_m_rdata),
    .i_lpddr_graph_2_targ_ht_axi_m_rid(i_lpddr_graph_2_targ_ht_axi_m_rid),
    .i_lpddr_graph_2_targ_ht_axi_m_rlast(i_lpddr_graph_2_targ_ht_axi_m_rlast),
    .o_lpddr_graph_2_targ_ht_axi_m_rready(o_lpddr_graph_2_targ_ht_axi_m_rready),
    .i_lpddr_graph_2_targ_ht_axi_m_rresp(i_lpddr_graph_2_targ_ht_axi_m_rresp),
    .i_lpddr_graph_2_targ_ht_axi_m_rvalid(i_lpddr_graph_2_targ_ht_axi_m_rvalid),
    .o_lpddr_graph_2_targ_ht_axi_m_wdata(o_lpddr_graph_2_targ_ht_axi_m_wdata),
    .o_lpddr_graph_2_targ_ht_axi_m_wlast(o_lpddr_graph_2_targ_ht_axi_m_wlast),
    .i_lpddr_graph_2_targ_ht_axi_m_wready(i_lpddr_graph_2_targ_ht_axi_m_wready),
    .o_lpddr_graph_2_targ_ht_axi_m_wstrb(o_lpddr_graph_2_targ_ht_axi_m_wstrb),
    .o_lpddr_graph_2_targ_ht_axi_m_wvalid(o_lpddr_graph_2_targ_ht_axi_m_wvalid),
    .o_lpddr_graph_2_targ_syscfg_apb_m_paddr(o_lpddr_graph_2_targ_syscfg_apb_m_paddr),
    .o_lpddr_graph_2_targ_syscfg_apb_m_penable(o_lpddr_graph_2_targ_syscfg_apb_m_penable),
    .o_lpddr_graph_2_targ_syscfg_apb_m_pprot(o_lpddr_graph_2_targ_syscfg_apb_m_pprot),
    .i_lpddr_graph_2_targ_syscfg_apb_m_prdata(i_lpddr_graph_2_targ_syscfg_apb_m_prdata),
    .i_lpddr_graph_2_targ_syscfg_apb_m_pready(i_lpddr_graph_2_targ_syscfg_apb_m_pready),
    .o_lpddr_graph_2_targ_syscfg_apb_m_psel(o_lpddr_graph_2_targ_syscfg_apb_m_psel),
    .i_lpddr_graph_2_targ_syscfg_apb_m_pslverr(i_lpddr_graph_2_targ_syscfg_apb_m_pslverr),
    .o_lpddr_graph_2_targ_syscfg_apb_m_pstrb(o_lpddr_graph_2_targ_syscfg_apb_m_pstrb),
    .o_lpddr_graph_2_targ_syscfg_apb_m_pwdata(o_lpddr_graph_2_targ_syscfg_apb_m_pwdata),
    .o_lpddr_graph_2_targ_syscfg_apb_m_pwrite(o_lpddr_graph_2_targ_syscfg_apb_m_pwrite),
    .i_lpddr_graph_3_aon_clk(i_lpddr_graph_3_aon_clk),
    .i_lpddr_graph_3_aon_rst_n(lpddr_graph_3_aon_rst_n_synced),
    .o_lpddr_graph_3_cfg_pwr_idle_val(o_lpddr_graph_3_cfg_pwr_idle_val),
    .o_lpddr_graph_3_cfg_pwr_idle_ack(o_lpddr_graph_3_cfg_pwr_idle_ack),
    .i_lpddr_graph_3_cfg_pwr_idle_req(i_lpddr_graph_3_cfg_pwr_idle_req),
    .i_lpddr_graph_3_clk(i_lpddr_graph_3_clk),
    .i_lpddr_graph_3_clken(i_lpddr_graph_3_clken),
    .o_lpddr_graph_3_pwr_idle_val(o_lpddr_graph_3_pwr_idle_val),
    .o_lpddr_graph_3_pwr_idle_ack(o_lpddr_graph_3_pwr_idle_ack),
    .i_lpddr_graph_3_pwr_idle_req(i_lpddr_graph_3_pwr_idle_req),
    .i_lpddr_graph_3_rst_n(i_lpddr_graph_3_rst_n),
    .o_lpddr_graph_3_targ_cfg_apb_m_paddr(o_lpddr_graph_3_targ_cfg_apb_m_paddr),
    .o_lpddr_graph_3_targ_cfg_apb_m_penable(o_lpddr_graph_3_targ_cfg_apb_m_penable),
    .o_lpddr_graph_3_targ_cfg_apb_m_pprot(o_lpddr_graph_3_targ_cfg_apb_m_pprot),
    .i_lpddr_graph_3_targ_cfg_apb_m_prdata(i_lpddr_graph_3_targ_cfg_apb_m_prdata),
    .i_lpddr_graph_3_targ_cfg_apb_m_pready(i_lpddr_graph_3_targ_cfg_apb_m_pready),
    .o_lpddr_graph_3_targ_cfg_apb_m_psel(o_lpddr_graph_3_targ_cfg_apb_m_psel),
    .i_lpddr_graph_3_targ_cfg_apb_m_pslverr(i_lpddr_graph_3_targ_cfg_apb_m_pslverr),
    .o_lpddr_graph_3_targ_cfg_apb_m_pstrb(o_lpddr_graph_3_targ_cfg_apb_m_pstrb),
    .o_lpddr_graph_3_targ_cfg_apb_m_pwdata(o_lpddr_graph_3_targ_cfg_apb_m_pwdata),
    .o_lpddr_graph_3_targ_cfg_apb_m_pwrite(o_lpddr_graph_3_targ_cfg_apb_m_pwrite),
    .o_lpddr_graph_3_targ_ht_axi_m_araddr(o_lpddr_graph_3_targ_ht_axi_m_araddr),
    .o_lpddr_graph_3_targ_ht_axi_m_arburst(o_lpddr_graph_3_targ_ht_axi_m_arburst),
    .o_lpddr_graph_3_targ_ht_axi_m_arcache(o_lpddr_graph_3_targ_ht_axi_m_arcache),
    .o_lpddr_graph_3_targ_ht_axi_m_arid(o_lpddr_graph_3_targ_ht_axi_m_arid),
    .o_lpddr_graph_3_targ_ht_axi_m_arlen(o_lpddr_graph_3_targ_ht_axi_m_arlen),
    .o_lpddr_graph_3_targ_ht_axi_m_arlock(o_lpddr_graph_3_targ_ht_axi_m_arlock),
    .o_lpddr_graph_3_targ_ht_axi_m_arprot(o_lpddr_graph_3_targ_ht_axi_m_arprot),
    .o_lpddr_graph_3_targ_ht_axi_m_arqos(o_lpddr_graph_3_targ_ht_axi_m_arqos),
    .i_lpddr_graph_3_targ_ht_axi_m_arready(i_lpddr_graph_3_targ_ht_axi_m_arready),
    .o_lpddr_graph_3_targ_ht_axi_m_arsize(o_lpddr_graph_3_targ_ht_axi_m_arsize),
    .o_lpddr_graph_3_targ_ht_axi_m_arvalid(o_lpddr_graph_3_targ_ht_axi_m_arvalid),
    .o_lpddr_graph_3_targ_ht_axi_m_awaddr(o_lpddr_graph_3_targ_ht_axi_m_awaddr),
    .o_lpddr_graph_3_targ_ht_axi_m_awburst(o_lpddr_graph_3_targ_ht_axi_m_awburst),
    .o_lpddr_graph_3_targ_ht_axi_m_awcache(o_lpddr_graph_3_targ_ht_axi_m_awcache),
    .o_lpddr_graph_3_targ_ht_axi_m_awid(o_lpddr_graph_3_targ_ht_axi_m_awid),
    .o_lpddr_graph_3_targ_ht_axi_m_awlen(o_lpddr_graph_3_targ_ht_axi_m_awlen),
    .o_lpddr_graph_3_targ_ht_axi_m_awlock(o_lpddr_graph_3_targ_ht_axi_m_awlock),
    .o_lpddr_graph_3_targ_ht_axi_m_awprot(o_lpddr_graph_3_targ_ht_axi_m_awprot),
    .o_lpddr_graph_3_targ_ht_axi_m_awqos(o_lpddr_graph_3_targ_ht_axi_m_awqos),
    .i_lpddr_graph_3_targ_ht_axi_m_awready(i_lpddr_graph_3_targ_ht_axi_m_awready),
    .o_lpddr_graph_3_targ_ht_axi_m_awsize(o_lpddr_graph_3_targ_ht_axi_m_awsize),
    .o_lpddr_graph_3_targ_ht_axi_m_awvalid(o_lpddr_graph_3_targ_ht_axi_m_awvalid),
    .i_lpddr_graph_3_targ_ht_axi_m_bid(i_lpddr_graph_3_targ_ht_axi_m_bid),
    .o_lpddr_graph_3_targ_ht_axi_m_bready(o_lpddr_graph_3_targ_ht_axi_m_bready),
    .i_lpddr_graph_3_targ_ht_axi_m_bresp(i_lpddr_graph_3_targ_ht_axi_m_bresp),
    .i_lpddr_graph_3_targ_ht_axi_m_bvalid(i_lpddr_graph_3_targ_ht_axi_m_bvalid),
    .i_lpddr_graph_3_targ_ht_axi_m_rdata(i_lpddr_graph_3_targ_ht_axi_m_rdata),
    .i_lpddr_graph_3_targ_ht_axi_m_rid(i_lpddr_graph_3_targ_ht_axi_m_rid),
    .i_lpddr_graph_3_targ_ht_axi_m_rlast(i_lpddr_graph_3_targ_ht_axi_m_rlast),
    .o_lpddr_graph_3_targ_ht_axi_m_rready(o_lpddr_graph_3_targ_ht_axi_m_rready),
    .i_lpddr_graph_3_targ_ht_axi_m_rresp(i_lpddr_graph_3_targ_ht_axi_m_rresp),
    .i_lpddr_graph_3_targ_ht_axi_m_rvalid(i_lpddr_graph_3_targ_ht_axi_m_rvalid),
    .o_lpddr_graph_3_targ_ht_axi_m_wdata(o_lpddr_graph_3_targ_ht_axi_m_wdata),
    .o_lpddr_graph_3_targ_ht_axi_m_wlast(o_lpddr_graph_3_targ_ht_axi_m_wlast),
    .i_lpddr_graph_3_targ_ht_axi_m_wready(i_lpddr_graph_3_targ_ht_axi_m_wready),
    .o_lpddr_graph_3_targ_ht_axi_m_wstrb(o_lpddr_graph_3_targ_ht_axi_m_wstrb),
    .o_lpddr_graph_3_targ_ht_axi_m_wvalid(o_lpddr_graph_3_targ_ht_axi_m_wvalid),
    .o_lpddr_graph_3_targ_syscfg_apb_m_paddr(o_lpddr_graph_3_targ_syscfg_apb_m_paddr),
    .o_lpddr_graph_3_targ_syscfg_apb_m_penable(o_lpddr_graph_3_targ_syscfg_apb_m_penable),
    .o_lpddr_graph_3_targ_syscfg_apb_m_pprot(o_lpddr_graph_3_targ_syscfg_apb_m_pprot),
    .i_lpddr_graph_3_targ_syscfg_apb_m_prdata(i_lpddr_graph_3_targ_syscfg_apb_m_prdata),
    .i_lpddr_graph_3_targ_syscfg_apb_m_pready(i_lpddr_graph_3_targ_syscfg_apb_m_pready),
    .o_lpddr_graph_3_targ_syscfg_apb_m_psel(o_lpddr_graph_3_targ_syscfg_apb_m_psel),
    .i_lpddr_graph_3_targ_syscfg_apb_m_pslverr(i_lpddr_graph_3_targ_syscfg_apb_m_pslverr),
    .o_lpddr_graph_3_targ_syscfg_apb_m_pstrb(o_lpddr_graph_3_targ_syscfg_apb_m_pstrb),
    .o_lpddr_graph_3_targ_syscfg_apb_m_pwdata(o_lpddr_graph_3_targ_syscfg_apb_m_pwdata),
    .o_lpddr_graph_3_targ_syscfg_apb_m_pwrite(o_lpddr_graph_3_targ_syscfg_apb_m_pwrite),
    .i_noc_clk(i_noc_clk),
    .i_noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
);

endmodule
