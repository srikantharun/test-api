const phy_init_data_t ddrctl_init2_details[string][] = '{
"A" : '{
'{step_type : POLL,	value:32'd0,	reg_addr:32'd66836},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd66836},
'{step_type:REG_WRITE,	value:32'd0,	reg_addr:32'd68736},
'{step_type:REG_WRITE,	value:32'd65556,	reg_addr:32'd66832},
'{step_type:REG_WRITE,	value:32'd1,	reg_addr:32'd68736},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd68740},
'{step_type:REG_WRITE,	value:32'd0,	reg_addr:32'd68736},
'{step_type:REG_WRITE,	value:32'd65557,	reg_addr:32'd66832},
'{step_type:REG_WRITE,	value:32'd1,	reg_addr:32'd68736},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd68740},
'{step_type:REG_WRITE,	value:32'd0,	reg_addr:32'd65920},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65556},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65556},
'{step_type : POLL,	value:32'd10468,	reg_addr:32'd2688},
'{step_type:REG_WRITE,	value:32'd10468,	reg_addr:32'd2688},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd9566,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd10334,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd10496,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd11776,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd9566,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd10334,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd10496,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd11776,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd2097152000,	reg_addr:32'd66840},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd4096,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd4096,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd4638,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd4638,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd432,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd432,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd699,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd699,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd774,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd774,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd2648,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd2648,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd2869,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd2869,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd3119,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd3119,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd3328,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd3328,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd3603,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd3603,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd3918,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd3918,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd4410,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd4410,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd4864,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd4864,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd5122,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd5122,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd5632,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd5632,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd5888,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd5888,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd6290,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd6290,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd6400,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd6400,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd7168,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd7168,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd9566,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd9566,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd10334,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd10334,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd10496,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd10496,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd16,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd11776,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483664,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd32,	reg_addr:32'd65664},
'{step_type:REG_WRITE,	value:32'd11776,	reg_addr:32'd65668},
'{step_type:REG_WRITE,	value:32'd2147483680,	reg_addr:32'd65664},
'{step_type : POLL,	value:32'd1,	reg_addr:32'd65680},
'{step_type : POLL,	value:32'd0,	reg_addr:32'd65680},
'{step_type:REG_WRITE,	value:32'd2097152001,	reg_addr:32'd66840},
'{step_type:REG_WRITE,	value:32'd0,	reg_addr:32'd66056},
'{step_type:REG_WRITE,	value:32'd0,	reg_addr:32'd65920},
'{step_type:REG_WRITE,	value:32'd1,	reg_addr:32'd65920},
'{step_type:REG_WRITE,	value:32'd1,	reg_addr:32'd65920},
'{step_type:REG_WRITE,	value:32'd1,	reg_addr:32'd65792},
'{step_type:REG_WRITE,	value:32'd10468,	reg_addr:32'd2688},
'{step_type:REG_WRITE,	value:32'd0,	reg_addr:32'd65920},
'{step_type : POLL,	value:32'd50855944,	reg_addr:32'd65536},
'{step_type:REG_WRITE,	value:32'd0,	reg_addr:32'd65920},
'{step_type : POLL,	value:32'd50855944,	reg_addr:32'd65536}

}};

