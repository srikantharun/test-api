//
// File: test_packages.svh
//
// Generated from Questa VIP Configurator (20240520)
// Generated using Questa VIP Library ( 2024.2 : 05/29/2024:10:31 )
//

import lpddr_subsystem_test_pkg::*;

// Add other packages here as required
