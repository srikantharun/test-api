// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: Milos Stanisavljevic <milos.stanisavljevic@axelera.ai>


/// TODO:__one_line_summary_of_lpddr_subsys_pkg__
///
package lpddr_subsys_pkg;

endpackage
