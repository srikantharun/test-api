// COPYRIGHT (c) Breker Verification Systems
// This software has been provided pursuant to a License Agreement
// containing restrictions on its use.  This software contains
// valuable trade secrets and proprietary information of
// Breker Verification Systems and is protected by law.  It may
// not be copied or distributed in any form or medium, disclosed
// to third parties, reverse engineered or used in any manner not
// provided for in said License Agreement except with the prior
// written authorization from Breker Verification Systems.
//
// Auto-generated by Breker TrekSoC version 2.1.3 at Wed Aug 28 07:36:38 2024



`ifndef GUARD__TREK_MASTER_PORT_DELAY_REQ_DELAY_REQ__SV
`define GUARD__TREK_MASTER_PORT_DELAY_REQ_DELAY_REQ__SV

class trek_master_port_delay_req_delay_req
    extends trek_master_port#(.T1(trek_delay_req),
                              .T2(trek_delay_req));

  function new(input string name = "");
    super.new(name);  // get_name() should return the tb_path
    trek_uvm_pkg::audit_port_info(.name(name),
        .port_type("trek_master_port_delay_req_delay_req"),
        .primary_type(T1::type_name),
        .secondary_type(T2::type_name));
    trek_uvm_pkg::port_built(name);
  endfunction

  // User methods are in the base class.
  // This method is called by the user methods to get
  // data from Trek via a "put_port" or a "master_port".
  //
  virtual function trek_delay_req pull(
    input trek_delay_req t = null, bit call_item_done = 1'b1);
    bit[63:0] tid;

    if (! trek_uvm_pkg::trek_started) begin: not_started
      `uvm_error({get_name(), "::pull()"},
        "You must start Trek before calling this function.")
      return null;
    end

    if (trek_uvm_events::end_of_test()) begin: test_is_done
      `uvm_info({get_name(), "::pull()"},
        "The trek test has already finished.", UVM_DEBUG)
      return null;
    end

    if (! trek_dpi_pkg::trek_can_get(get_name())) begin: nothing_there
      `uvm_error({get_name(), "::pull()"},
        {"You must ensure the port 'trek_delay_port' has",
        " a transaction ready to retrieve before calling this function."})
      return null;
    end

    if (t == null) begin: no_object_provided
      t = T1::type_id::create("req");
    end

    tid = trek_get_transaction_id(get_name());
    if ((tid[63:31] == 33'h1_ffff_ffff) || (tid[63:32] == 32'h0000_0000))
    begin: _tid
      t.set_transaction_id(tid);
    end else begin: _no_tid
      `uvm_error(get_name(), $sformatf({"PSS uses a 64-bit transaction_id",
           " but UVM uses a 32-bit signed integer. Your transaction_id ",
           "(64'h%016h) does not fit in a 32-bit signed integer."}, tid))
    end

    t.m_delay = trek_get_longint_unsigned(get_name(), "m_delay");

    if (call_item_done) begin: pop_transaction_with_no_response
      item_done();
    end
    return t;
  endfunction: pull

  // User methods are in the base class.
  // This method is called by the user methods to send
  // data to Trek via a "check_port" or a "master_port".
  //
  virtual function void push(input trek_delay_req t);
    int errno = 0;
    // Trek5 uses a 64-bit unsigned id, but uvm uses a 32-bit signed id
    errno += trek_put_transaction_id(get_name(), t.get_transaction_id());
    errno += trek_put_longint_unsigned(get_name(), "m_delay", t.m_delay);
    errno += trek_put_done(get_name()); 
    if (errno != 0) begin: bad_return_status
      `uvm_fatal(get_name(), {"trek_master_port_delay_req_delay_req::push(",
          get_name(), ") encountered non-zero return status"})
    end
  endfunction: push

endclass: trek_master_port_delay_req_delay_req

`endif  // GUARD__TREK_MASTER_PORT_DELAY_REQ_DELAY_REQ__SV
