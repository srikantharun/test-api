// (C) Copyright Axelera AI 2024
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description:
// UVM Scoreboards
// Pre-configured scoreboards for testbench construction
// Owner: abond

// Package: axe_uvm_scoreboard_pkg 
package axe_uvm_scoreboard_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  `include "axe_uvm_scoreboard.svh"
  `include "axe_uvm_indexed_scoreboard.svh"

endpackage : axe_uvm_scoreboard_pkg
