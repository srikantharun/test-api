// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Owner: andrew dickson <andrew.dickson@axelera.ai>

// Assertions to check connectivity for the deubgger
// I/Os to debugger IP in soc_mgmt

always_comb begin

  a_dbg_con000 : assert #0 ( o_debugint         === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_debugint         ) else con_fail_rpt("o_debugint         ", o_debugint        , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_debugint        );
  a_dbg_con001 : assert #0 ( o_resethaltreq     === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_resethaltreq     ) else con_fail_rpt("o_resethaltreq     ", o_resethaltreq    , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_resethaltreq    );
  a_dbg_con004 : assert #0 ( i_hart_unavail     === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_hart_unavail     ) else con_fail_rpt("i_hart_unavail     ", i_hart_unavail    , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_hart_unavail    );
  a_dbg_con005 : assert #0 ( i_hart_under_reset === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_hart_under_reset ) else con_fail_rpt("i_hart_under_reset ", i_hart_under_reset, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_hart_under_reset);
  a_dbg_con006 : assert #0 ( o_lt_axi_m_awid    === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awid         ) else con_fail_rpt("o_lt_axi_m_awid    ", o_lt_axi_m_awid   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awid        );
  a_dbg_con007 : assert #0 ( o_lt_axi_m_awaddr  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awaddr       ) else con_fail_rpt("o_lt_axi_m_awaddr  ", o_lt_axi_m_awaddr , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awaddr      );
  a_dbg_con008 : assert #0 ( o_lt_axi_m_awlen   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awlen        ) else con_fail_rpt("o_lt_axi_m_awlen   ", o_lt_axi_m_awlen  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awlen       );
  a_dbg_con009 : assert #0 ( o_lt_axi_m_awsize  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awsize       ) else con_fail_rpt("o_lt_axi_m_awsize  ", o_lt_axi_m_awsize , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awsize      );
  a_dbg_con010 : assert #0 ( o_lt_axi_m_awburst === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awburst      ) else con_fail_rpt("o_lt_axi_m_awburst ", o_lt_axi_m_awburst, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awburst     );
  a_dbg_con011 : assert #0 ( o_lt_axi_m_awlock  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awlock       ) else con_fail_rpt("o_lt_axi_m_awlock  ", o_lt_axi_m_awlock , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awlock      );
  a_dbg_con012 : assert #0 ( o_lt_axi_m_awcache === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awcache      ) else con_fail_rpt("o_lt_axi_m_awcache ", o_lt_axi_m_awcache, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awcache     );
  a_dbg_con013 : assert #0 ( o_lt_axi_m_awprot  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awprot       ) else con_fail_rpt("o_lt_axi_m_awprot  ", o_lt_axi_m_awprot , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awprot      );
  a_dbg_con014 : assert #0 ( o_lt_axi_m_awvalid === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awvalid      ) else con_fail_rpt("o_lt_axi_m_awvalid ", o_lt_axi_m_awvalid, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_awvalid     );
  a_dbg_con015 : assert #0 ( i_lt_axi_m_awready === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_awready      ) else con_fail_rpt("i_lt_axi_m_awready ", i_lt_axi_m_awready, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_awready     );
  a_dbg_con016 : assert #0 ( o_lt_axi_m_wdata   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_wdata        ) else con_fail_rpt("o_lt_axi_m_wdata   ", o_lt_axi_m_wdata  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_wdata       );
  a_dbg_con017 : assert #0 ( o_lt_axi_m_wstrb   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_wstrb        ) else con_fail_rpt("o_lt_axi_m_wstrb   ", o_lt_axi_m_wstrb  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_wstrb       );
  a_dbg_con018 : assert #0 ( o_lt_axi_m_wlast   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_wlast        ) else con_fail_rpt("o_lt_axi_m_wlast   ", o_lt_axi_m_wlast  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_wlast       );
  a_dbg_con019 : assert #0 ( o_lt_axi_m_wvalid  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_wvalid       ) else con_fail_rpt("o_lt_axi_m_wvalid  ", o_lt_axi_m_wvalid , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_wvalid      );
  a_dbg_con020 : assert #0 ( i_lt_axi_m_wready  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_wready       ) else con_fail_rpt("i_lt_axi_m_wready  ", i_lt_axi_m_wready , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_wready      );
  a_dbg_con021 : assert #0 ( i_lt_axi_m_bid     === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_bid          ) else con_fail_rpt("i_lt_axi_m_bid     ", i_lt_axi_m_bid    , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_bid         );
  a_dbg_con022 : assert #0 ( i_lt_axi_m_bresp   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_bresp        ) else con_fail_rpt("i_lt_axi_m_bresp   ", i_lt_axi_m_bresp  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_bresp       );
  a_dbg_con023 : assert #0 ( i_lt_axi_m_bvalid  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_bvalid       ) else con_fail_rpt("i_lt_axi_m_bvalid  ", i_lt_axi_m_bvalid , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_bvalid      );
  a_dbg_con024 : assert #0 ( o_lt_axi_m_bready  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_bready       ) else con_fail_rpt("o_lt_axi_m_bready  ", o_lt_axi_m_bready , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_bready      );
  a_dbg_con025 : assert #0 ( o_lt_axi_m_arid    === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arid         ) else con_fail_rpt("o_lt_axi_m_arid    ", o_lt_axi_m_arid   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arid        );
  a_dbg_con026 : assert #0 ( o_lt_axi_m_araddr  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_araddr       ) else con_fail_rpt("o_lt_axi_m_araddr  ", o_lt_axi_m_araddr , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_araddr      );
  a_dbg_con027 : assert #0 ( o_lt_axi_m_arlen   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arlen        ) else con_fail_rpt("o_lt_axi_m_arlen   ", o_lt_axi_m_arlen  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arlen       );
  a_dbg_con028 : assert #0 ( o_lt_axi_m_arsize  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arsize       ) else con_fail_rpt("o_lt_axi_m_arsize  ", o_lt_axi_m_arsize , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arsize      );
  a_dbg_con029 : assert #0 ( o_lt_axi_m_arburst === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arburst      ) else con_fail_rpt("o_lt_axi_m_arburst ", o_lt_axi_m_arburst, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arburst     );
  a_dbg_con030 : assert #0 ( o_lt_axi_m_arlock  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arlock       ) else con_fail_rpt("o_lt_axi_m_arlock  ", o_lt_axi_m_arlock , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arlock      );
  a_dbg_con031 : assert #0 ( o_lt_axi_m_arcache === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arcache      ) else con_fail_rpt("o_lt_axi_m_arcache ", o_lt_axi_m_arcache, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arcache     );
  a_dbg_con032 : assert #0 ( o_lt_axi_m_arprot  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arprot       ) else con_fail_rpt("o_lt_axi_m_arprot  ", o_lt_axi_m_arprot , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arprot      );
  a_dbg_con033 : assert #0 ( o_lt_axi_m_arvalid === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arvalid      ) else con_fail_rpt("o_lt_axi_m_arvalid ", o_lt_axi_m_arvalid, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_arvalid     );
  a_dbg_con034 : assert #0 ( i_lt_axi_m_arready === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_arready      ) else con_fail_rpt("i_lt_axi_m_arready ", i_lt_axi_m_arready, i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_arready     );
  a_dbg_con035 : assert #0 ( i_lt_axi_m_rid     === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rid          ) else con_fail_rpt("i_lt_axi_m_rid     ", i_lt_axi_m_rid    , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rid         );
  a_dbg_con036 : assert #0 ( i_lt_axi_m_rdata   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rdata        ) else con_fail_rpt("i_lt_axi_m_rdata   ", i_lt_axi_m_rdata  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rdata       );
  a_dbg_con037 : assert #0 ( i_lt_axi_m_rresp   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rresp        ) else con_fail_rpt("i_lt_axi_m_rresp   ", i_lt_axi_m_rresp  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rresp       );
  a_dbg_con038 : assert #0 ( i_lt_axi_m_rlast   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rlast        ) else con_fail_rpt("i_lt_axi_m_rlast   ", i_lt_axi_m_rlast  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rlast       );
  a_dbg_con039 : assert #0 ( i_lt_axi_m_rvalid  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rvalid       ) else con_fail_rpt("i_lt_axi_m_rvalid  ", i_lt_axi_m_rvalid , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_sys_rvalid      );
  a_dbg_con040 : assert #0 ( o_lt_axi_m_rready  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_rready       ) else con_fail_rpt("o_lt_axi_m_rready  ", o_lt_axi_m_rready , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_sys_rready      );

  a_dbg_con100 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arready === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_arready   ) else con_fail_rpt("o_rv_arready ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arready , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_arready   );
  a_dbg_con101 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awready === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_awready   ) else con_fail_rpt("o_rv_awready ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awready , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_awready   );
  a_dbg_con102 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_bid     === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_bid       ) else con_fail_rpt("o_rv_bid     ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_bid     , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_bid       );
  a_dbg_con103 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_bresp   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_bresp     ) else con_fail_rpt("o_rv_bresp   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_bresp   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_bresp     );
  a_dbg_con104 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_bvalid  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_bvalid    ) else con_fail_rpt("o_rv_bvalid  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_bvalid  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_bvalid    );
  a_dbg_con105 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rdata   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rdata     ) else con_fail_rpt("o_rv_rdata   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rdata   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rdata     );
  a_dbg_con106 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rid     === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rid       ) else con_fail_rpt("o_rv_rid     ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rid     , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rid       );
  a_dbg_con107 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rlast   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rlast     ) else con_fail_rpt("o_rv_rlast   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rlast   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rlast     );
  a_dbg_con108 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rresp   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rresp     ) else con_fail_rpt("o_rv_rresp   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rresp   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rresp     );
  a_dbg_con109 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rvalid  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rvalid    ) else con_fail_rpt("o_rv_rvalid  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rvalid  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_rvalid    );
  a_dbg_con110 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wready  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_wready    ) else con_fail_rpt("o_rv_wready  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wready  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.o_rv_wready    );
  a_dbg_con111 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_araddr  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_araddr    ) else con_fail_rpt("i_rv_araddr  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_araddr  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_araddr    );
  a_dbg_con112 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arburst === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arburst   ) else con_fail_rpt("i_rv_arburst ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arburst , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arburst   );
  a_dbg_con113 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arcache === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arcache   ) else con_fail_rpt("i_rv_arcache ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arcache , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arcache   );
  a_dbg_con114 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arid    === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arid      ) else con_fail_rpt("i_rv_arid    ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arid    , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arid      );
  a_dbg_con115 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arlen   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arlen     ) else con_fail_rpt("i_rv_arlen   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arlen   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arlen     );
  a_dbg_con116 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arlock  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arlock    ) else con_fail_rpt("i_rv_arlock  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arlock  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arlock    );
  a_dbg_con117 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arprot  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arprot    ) else con_fail_rpt("i_rv_arprot  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arprot  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arprot    );
  a_dbg_con118 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arsize  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arsize    ) else con_fail_rpt("i_rv_arsize  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arsize  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arsize    );
  a_dbg_con119 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arvalid === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arvalid   ) else con_fail_rpt("i_rv_arvalid ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_arvalid , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_arvalid   );
  a_dbg_con120 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awaddr  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awaddr    ) else con_fail_rpt("i_rv_awaddr  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awaddr  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awaddr    );
  a_dbg_con121 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awburst === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awburst   ) else con_fail_rpt("i_rv_awburst ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awburst , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awburst   );
  a_dbg_con122 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awcache === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awcache   ) else con_fail_rpt("i_rv_awcache ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awcache , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awcache   );
  a_dbg_con123 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awid    === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awid      ) else con_fail_rpt("i_rv_awid    ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awid    , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awid      );
  a_dbg_con124 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awlen   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awlen     ) else con_fail_rpt("i_rv_awlen   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awlen   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awlen     );
  a_dbg_con125 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awlock  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awlock    ) else con_fail_rpt("i_rv_awlock  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awlock  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awlock    );
  a_dbg_con126 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awprot  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awprot    ) else con_fail_rpt("i_rv_awprot  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awprot  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awprot    );
  a_dbg_con127 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awsize  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awsize    ) else con_fail_rpt("i_rv_awsize  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awsize  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awsize    );
  a_dbg_con128 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awvalid === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awvalid   ) else con_fail_rpt("i_rv_awvalid ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_awvalid , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_awvalid   );
  a_dbg_con129 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_bready  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_bready    ) else con_fail_rpt("i_rv_bready  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_bready  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_bready    );
  a_dbg_con130 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rready  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_rready    ) else con_fail_rpt("i_rv_rready  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_rready  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_rready    );
  a_dbg_con131 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wdata   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_wdata     ) else con_fail_rpt("i_rv_wdata   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wdata   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_wdata     );
  a_dbg_con132 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wlast   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_wlast     ) else con_fail_rpt("i_rv_wlast   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wlast   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_wlast     );
  a_dbg_con133 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wstrb   === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_wstrb     ) else con_fail_rpt("i_rv_wstrb   ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wstrb   , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_wstrb     );
  a_dbg_con134 : assert #0 ( i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wvalid  === i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_wvalid    ) else con_fail_rpt("i_rv_wvalid  ", i_soc_mgmt_p_dut.u_soc_mgmt.u_soc_mgmt_bus_fabric_wrapper.u_smu_fabric_subsys.ex_smu_axi_fabric_lt_axi_dbgr_m_wvalid  , i_soc_mgmt_p_dut.u_soc_mgmt.u_nds_pldm_wrapper.i_rv_wvalid    );

end

function void con_fail_rpt(string sig_name, logic [63:0] lhs, rhs);
  `uvm_error("DEBUG_ASSERT", $sformatf("ERROR Assertion failed for signal %0s LHS: %0x RHS: %0x", sig_name, lhs, rhs))
  fail_cnt++;
endfunction



