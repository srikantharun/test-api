`ifndef RAL_DWC_DDRPHYA_DBYTE3_P1_PKG
`define RAL_DWC_DDRPHYA_DBYTE3_P1_PKG

package ral_DWC_DDRPHYA_DBYTE3_p1_pkg;
import uvm_pkg::*;

class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DFIMRL_p1 extends uvm_reg;
	rand uvm_reg_field DFIMRL_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DFIMRL_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DFIMRL_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DFIMRL_p1 = uvm_reg_field::type_id::create("DFIMRL_p1",,get_full_name());
      this.DFIMRL_p1.configure(this, 6, 0, "RW", 0, 6'h6, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DFIMRL_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DFIMRL_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_EnableWriteLinkEcc_p1 extends uvm_reg;
	rand uvm_reg_field EnableWriteLinkEcc_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   EnableWriteLinkEcc_p1: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_EnableWriteLinkEcc_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.EnableWriteLinkEcc_p1 = uvm_reg_field::type_id::create("EnableWriteLinkEcc_p1",,get_full_name());
      this.EnableWriteLinkEcc_p1.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_EnableWriteLinkEcc_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_EnableWriteLinkEcc_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxDfiClkDis_p1 extends uvm_reg;
	rand uvm_reg_field DfiClkDqDis;
	rand uvm_reg_field DfiClkDqsDis;
	rand uvm_reg_field DfiClkWckDis;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DfiClkDqDis: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	   DfiClkDqsDis: coverpoint {m_data[9:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   DfiClkWckDis: coverpoint {m_data[10:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DxDfiClkDis_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DfiClkDqDis = uvm_reg_field::type_id::create("DfiClkDqDis",,get_full_name());
      this.DfiClkDqDis.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 0);
      this.DfiClkDqsDis = uvm_reg_field::type_id::create("DfiClkDqsDis",,get_full_name());
      this.DfiClkDqsDis.configure(this, 1, 9, "RW", 0, 1'h0, 1, 0, 0);
      this.DfiClkWckDis = uvm_reg_field::type_id::create("DfiClkWckDis",,get_full_name());
      this.DfiClkWckDis.configure(this, 1, 10, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxDfiClkDis_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxDfiClkDis_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPClkDis_p1 extends uvm_reg;
	rand uvm_reg_field PClkDqDis;
	rand uvm_reg_field PClkDqsDis;
	rand uvm_reg_field PClkWckDis;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PClkDqDis: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	   PClkDqsDis: coverpoint {m_data[9:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PClkWckDis: coverpoint {m_data[10:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DxPClkDis_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PClkDqDis = uvm_reg_field::type_id::create("PClkDqDis",,get_full_name());
      this.PClkDqDis.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 0);
      this.PClkDqsDis = uvm_reg_field::type_id::create("PClkDqsDis",,get_full_name());
      this.PClkDqsDis.configure(this, 1, 9, "RW", 0, 1'h0, 1, 0, 0);
      this.PClkWckDis = uvm_reg_field::type_id::create("PClkWckDis",,get_full_name());
      this.PClkWckDis.configure(this, 1, 10, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPClkDis_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPClkDis_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_LP5DfiDataEnLatency_p1 extends uvm_reg;
	rand uvm_reg_field LP5RLm13;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   LP5RLm13: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_LP5DfiDataEnLatency_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.LP5RLm13 = uvm_reg_field::type_id::create("LP5RLm13",,get_full_name());
      this.LP5RLm13.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_LP5DfiDataEnLatency_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_LP5DfiDataEnLatency_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg0_p1 extends uvm_reg;
	rand uvm_reg_field PptDqsCntInvTrnTg0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PptDqsCntInvTrnTg0_p1: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PptDqsCntInvTrnTg0_p1 = uvm_reg_field::type_id::create("PptDqsCntInvTrnTg0_p1",,get_full_name());
      this.PptDqsCntInvTrnTg0_p1.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg1_p1 extends uvm_reg;
	rand uvm_reg_field PptDqsCntInvTrnTg1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PptDqsCntInvTrnTg1_p1: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PptDqsCntInvTrnTg1_p1 = uvm_reg_field::type_id::create("PptDqsCntInvTrnTg1_p1",,get_full_name());
      this.PptDqsCntInvTrnTg1_p1.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TrackingModeCntrl_p1 extends uvm_reg;
	rand uvm_reg_field EnWck2DqoSnoopTracking;
	rand uvm_reg_field Twck2dqoTrackingLimit;
	rand uvm_reg_field ReservedTrackingModeCntrl;
	rand uvm_reg_field Tdqs2dqTrackingLimit;
	rand uvm_reg_field DqsOscRunTimeSel;
	rand uvm_reg_field RxDqsTrackingThreshold;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   EnWck2DqoSnoopTracking: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   Twck2dqoTrackingLimit: coverpoint {m_data[3:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	   ReservedTrackingModeCntrl: coverpoint {m_data[4:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   Tdqs2dqTrackingLimit: coverpoint {m_data[7:5], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	   DqsOscRunTimeSel: coverpoint {m_data[11:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   RxDqsTrackingThreshold: coverpoint {m_data[14:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TrackingModeCntrl_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.EnWck2DqoSnoopTracking = uvm_reg_field::type_id::create("EnWck2DqoSnoopTracking",,get_full_name());
      this.EnWck2DqoSnoopTracking.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.Twck2dqoTrackingLimit = uvm_reg_field::type_id::create("Twck2dqoTrackingLimit",,get_full_name());
      this.Twck2dqoTrackingLimit.configure(this, 3, 1, "RW", 0, 3'h0, 1, 0, 0);
      this.ReservedTrackingModeCntrl = uvm_reg_field::type_id::create("ReservedTrackingModeCntrl",,get_full_name());
      this.ReservedTrackingModeCntrl.configure(this, 1, 4, "RW", 0, 1'h0, 1, 0, 0);
      this.Tdqs2dqTrackingLimit = uvm_reg_field::type_id::create("Tdqs2dqTrackingLimit",,get_full_name());
      this.Tdqs2dqTrackingLimit.configure(this, 3, 5, "RW", 0, 3'h0, 1, 0, 0);
      this.DqsOscRunTimeSel = uvm_reg_field::type_id::create("DqsOscRunTimeSel",,get_full_name());
      this.DqsOscRunTimeSel.configure(this, 4, 8, "RW", 0, 4'h3, 1, 0, 0);
      this.RxDqsTrackingThreshold = uvm_reg_field::type_id::create("RxDqsTrackingThreshold",,get_full_name());
      this.RxDqsTrackingThreshold.configure(this, 3, 12, "RW", 0, 3'h1, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TrackingModeCntrl_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TrackingModeCntrl_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r0_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r0_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r0_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r0_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r0_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r0_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r0_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r0_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r0_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r0_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r0_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r0_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r0_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r0_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r0_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r0_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg0_p1 extends uvm_reg;
	rand uvm_reg_field PptWck2DqoCntInvTrnTg0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PptWck2DqoCntInvTrnTg0_p1: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PptWck2DqoCntInvTrnTg0_p1 = uvm_reg_field::type_id::create("PptWck2DqoCntInvTrnTg0_p1",,get_full_name());
      this.PptWck2DqoCntInvTrnTg0_p1.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg1_p1 extends uvm_reg;
	rand uvm_reg_field PptWck2DqoCntInvTrnTg1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PptWck2DqoCntInvTrnTg1_p1: coverpoint {m_data[15:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {17'b???????????????00};
	      wildcard bins bit_0_wr_as_1 = {17'b???????????????10};
	      wildcard bins bit_0_rd_as_0 = {17'b???????????????01};
	      wildcard bins bit_0_rd_as_1 = {17'b???????????????11};
	      wildcard bins bit_1_wr_as_0 = {17'b??????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {17'b??????????????1?0};
	      wildcard bins bit_1_rd_as_0 = {17'b??????????????0?1};
	      wildcard bins bit_1_rd_as_1 = {17'b??????????????1?1};
	      wildcard bins bit_2_wr_as_0 = {17'b?????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {17'b?????????????1??0};
	      wildcard bins bit_2_rd_as_0 = {17'b?????????????0??1};
	      wildcard bins bit_2_rd_as_1 = {17'b?????????????1??1};
	      wildcard bins bit_3_wr_as_0 = {17'b????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {17'b????????????1???0};
	      wildcard bins bit_3_rd_as_0 = {17'b????????????0???1};
	      wildcard bins bit_3_rd_as_1 = {17'b????????????1???1};
	      wildcard bins bit_4_wr_as_0 = {17'b???????????0????0};
	      wildcard bins bit_4_wr_as_1 = {17'b???????????1????0};
	      wildcard bins bit_4_rd_as_0 = {17'b???????????0????1};
	      wildcard bins bit_4_rd_as_1 = {17'b???????????1????1};
	      wildcard bins bit_5_wr_as_0 = {17'b??????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {17'b??????????1?????0};
	      wildcard bins bit_5_rd_as_0 = {17'b??????????0?????1};
	      wildcard bins bit_5_rd_as_1 = {17'b??????????1?????1};
	      wildcard bins bit_6_wr_as_0 = {17'b?????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {17'b?????????1??????0};
	      wildcard bins bit_6_rd_as_0 = {17'b?????????0??????1};
	      wildcard bins bit_6_rd_as_1 = {17'b?????????1??????1};
	      wildcard bins bit_7_wr_as_0 = {17'b????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {17'b????????1???????0};
	      wildcard bins bit_7_rd_as_0 = {17'b????????0???????1};
	      wildcard bins bit_7_rd_as_1 = {17'b????????1???????1};
	      wildcard bins bit_8_wr_as_0 = {17'b???????0????????0};
	      wildcard bins bit_8_wr_as_1 = {17'b???????1????????0};
	      wildcard bins bit_8_rd_as_0 = {17'b???????0????????1};
	      wildcard bins bit_8_rd_as_1 = {17'b???????1????????1};
	      wildcard bins bit_9_wr_as_0 = {17'b??????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {17'b??????1?????????0};
	      wildcard bins bit_9_rd_as_0 = {17'b??????0?????????1};
	      wildcard bins bit_9_rd_as_1 = {17'b??????1?????????1};
	      wildcard bins bit_10_wr_as_0 = {17'b?????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {17'b?????1??????????0};
	      wildcard bins bit_10_rd_as_0 = {17'b?????0??????????1};
	      wildcard bins bit_10_rd_as_1 = {17'b?????1??????????1};
	      wildcard bins bit_11_wr_as_0 = {17'b????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {17'b????1???????????0};
	      wildcard bins bit_11_rd_as_0 = {17'b????0???????????1};
	      wildcard bins bit_11_rd_as_1 = {17'b????1???????????1};
	      wildcard bins bit_12_wr_as_0 = {17'b???0????????????0};
	      wildcard bins bit_12_wr_as_1 = {17'b???1????????????0};
	      wildcard bins bit_12_rd_as_0 = {17'b???0????????????1};
	      wildcard bins bit_12_rd_as_1 = {17'b???1????????????1};
	      wildcard bins bit_13_wr_as_0 = {17'b??0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {17'b??1?????????????0};
	      wildcard bins bit_13_rd_as_0 = {17'b??0?????????????1};
	      wildcard bins bit_13_rd_as_1 = {17'b??1?????????????1};
	      wildcard bins bit_14_wr_as_0 = {17'b?0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {17'b?1??????????????0};
	      wildcard bins bit_14_rd_as_0 = {17'b?0??????????????1};
	      wildcard bins bit_14_rd_as_1 = {17'b?1??????????????1};
	      wildcard bins bit_15_wr_as_0 = {17'b0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {17'b1???????????????0};
	      wildcard bins bit_15_rd_as_0 = {17'b0???????????????1};
	      wildcard bins bit_15_rd_as_1 = {17'b1???????????????1};
	      option.weight = 64;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PptWck2DqoCntInvTrnTg1_p1 = uvm_reg_field::type_id::create("PptWck2DqoCntInvTrnTg1_p1",,get_full_name());
      this.PptWck2DqoCntInvTrnTg1_p1.configure(this, 16, 0, "RW", 0, 16'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqsLeftEyeOffsetTg0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqsLeftEyeOffsetTg0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqsLeftEyeOffsetTg0_p1 = uvm_reg_field::type_id::create("TxDqsLeftEyeOffsetTg0_p1",,get_full_name());
      this.TxDqsLeftEyeOffsetTg0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqsLeftEyeOffsetTg1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqsLeftEyeOffsetTg1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqsLeftEyeOffsetTg1_p1 = uvm_reg_field::type_id::create("TxDqsLeftEyeOffsetTg1_p1",,get_full_name());
      this.TxDqsLeftEyeOffsetTg1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg0_p1 extends uvm_reg;
	rand uvm_reg_field RxEnDlyTg0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxEnDlyTg0_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxEnDlyTg0_p1 = uvm_reg_field::type_id::create("RxEnDlyTg0_p1",,get_full_name());
      this.RxEnDlyTg0_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg1_p1 extends uvm_reg;
	rand uvm_reg_field RxEnDlyTg1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxEnDlyTg1_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxEnDlyTg1_p1 = uvm_reg_field::type_id::create("RxEnDlyTg1_p1",,get_full_name());
      this.RxEnDlyTg1_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqsRightEyeOffsetTg0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqsRightEyeOffsetTg0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqsRightEyeOffsetTg0_p1 = uvm_reg_field::type_id::create("TxDqsRightEyeOffsetTg0_p1",,get_full_name());
      this.TxDqsRightEyeOffsetTg0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqsRightEyeOffsetTg1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqsRightEyeOffsetTg1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqsRightEyeOffsetTg1_p1 = uvm_reg_field::type_id::create("TxDqsRightEyeOffsetTg1_p1",,get_full_name());
      this.TxDqsRightEyeOffsetTg1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqsPreambleControl_p1 extends uvm_reg;
	uvm_reg_field Reserved;
	rand uvm_reg_field LP4PostambleExt;
	rand uvm_reg_field WDQSEXTENSION;
	rand uvm_reg_field WCKEXTENSION;
	rand uvm_reg_field DqPreOeExt;
	rand uvm_reg_field DqPstOeExt;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   Reserved: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd = {7'b??????1};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd = {7'b??????1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd = {7'b??????1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd = {7'b??????1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd = {7'b??????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd = {7'b??????1};
	      option.weight = 18;
	   }
	   LP4PostambleExt: coverpoint {m_data[6:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   WDQSEXTENSION: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   WCKEXTENSION: coverpoint {m_data[8:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   DqPreOeExt: coverpoint {m_data[9:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   DqPstOeExt: coverpoint {m_data[10:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqsPreambleControl_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.Reserved = uvm_reg_field::type_id::create("Reserved",,get_full_name());
      this.Reserved.configure(this, 6, 0, "RO", 1, 6'h0, 1, 0, 0);
      this.LP4PostambleExt = uvm_reg_field::type_id::create("LP4PostambleExt",,get_full_name());
      this.LP4PostambleExt.configure(this, 1, 6, "RW", 0, 1'h0, 1, 0, 0);
      this.WDQSEXTENSION = uvm_reg_field::type_id::create("WDQSEXTENSION",,get_full_name());
      this.WDQSEXTENSION.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.WCKEXTENSION = uvm_reg_field::type_id::create("WCKEXTENSION",,get_full_name());
      this.WCKEXTENSION.configure(this, 1, 8, "RW", 0, 1'h0, 1, 0, 0);
      this.DqPreOeExt = uvm_reg_field::type_id::create("DqPreOeExt",,get_full_name());
      this.DqPreOeExt.configure(this, 1, 9, "RW", 0, 1'h0, 1, 0, 0);
      this.DqPstOeExt = uvm_reg_field::type_id::create("DqPstOeExt",,get_full_name());
      this.DqPstOeExt.configure(this, 1, 10, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqsPreambleControl_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqsPreambleControl_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DbyteRxDqsModeCntrl_p1 extends uvm_reg;
	rand uvm_reg_field RxPostambleMode;
	rand uvm_reg_field RxPreambleMode;
	rand uvm_reg_field LPDDR5RdqsEn;
	rand uvm_reg_field LPDDR5RdqsPre;
	rand uvm_reg_field LPDDR5RdqsPst;
	rand uvm_reg_field PositionDfeInit;
	rand uvm_reg_field PositionRxPhaseUpdate;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxPostambleMode: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxPreambleMode: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   LPDDR5RdqsEn: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   LPDDR5RdqsPre: coverpoint {m_data[4:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	   LPDDR5RdqsPst: coverpoint {m_data[6:5], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	   PositionDfeInit: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PositionRxPhaseUpdate: coverpoint {m_data[8:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DbyteRxDqsModeCntrl_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxPostambleMode = uvm_reg_field::type_id::create("RxPostambleMode",,get_full_name());
      this.RxPostambleMode.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.RxPreambleMode = uvm_reg_field::type_id::create("RxPreambleMode",,get_full_name());
      this.RxPreambleMode.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.LPDDR5RdqsEn = uvm_reg_field::type_id::create("LPDDR5RdqsEn",,get_full_name());
      this.LPDDR5RdqsEn.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
      this.LPDDR5RdqsPre = uvm_reg_field::type_id::create("LPDDR5RdqsPre",,get_full_name());
      this.LPDDR5RdqsPre.configure(this, 2, 3, "RW", 0, 2'h0, 1, 0, 0);
      this.LPDDR5RdqsPst = uvm_reg_field::type_id::create("LPDDR5RdqsPst",,get_full_name());
      this.LPDDR5RdqsPst.configure(this, 2, 5, "RW", 0, 2'h0, 1, 0, 0);
      this.PositionDfeInit = uvm_reg_field::type_id::create("PositionDfeInit",,get_full_name());
      this.PositionDfeInit.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.PositionRxPhaseUpdate = uvm_reg_field::type_id::create("PositionRxPhaseUpdate",,get_full_name());
      this.PositionRxPhaseUpdate.configure(this, 1, 8, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DbyteRxDqsModeCntrl_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DbyteRxDqsModeCntrl_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCntl1_p1 extends uvm_reg;
	rand uvm_reg_field EnRxClkCor;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   EnRxClkCor: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCntl1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.EnRxClkCor = uvm_reg_field::type_id::create("EnRxClkCor",,get_full_name());
      this.EnRxClkCor.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCntl1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCntl1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqsDlyTg0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqsDlyTg0_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqsDlyTg0_p1 = uvm_reg_field::type_id::create("TxDqsDlyTg0_p1",,get_full_name());
      this.TxDqsDlyTg0_p1.configure(this, 10, 0, "RW", 0, 10'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqsDlyTg1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqsDlyTg1_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqsDlyTg1_p1 = uvm_reg_field::type_id::create("TxDqsDlyTg1_p1",,get_full_name());
      this.TxDqsDlyTg1_p1.configure(this, 10, 0, "RW", 0, 10'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg0_p1 extends uvm_reg;
	rand uvm_reg_field TxWckDlyTg0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxWckDlyTg0_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxWckDlyTg0_p1 = uvm_reg_field::type_id::create("TxWckDlyTg0_p1",,get_full_name());
      this.TxWckDlyTg0_p1.configure(this, 12, 0, "RW", 0, 12'h200, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg1_p1 extends uvm_reg;
	rand uvm_reg_field TxWckDlyTg1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxWckDlyTg1_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxWckDlyTg1_p1 = uvm_reg_field::type_id::create("TxWckDlyTg1_p1",,get_full_name());
      this.TxWckDlyTg1_p1.configure(this, 12, 0, "RW", 0, 12'h200, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxModeCtlRxReplica_p1 extends uvm_reg;
	rand uvm_reg_field RxModeCtlRxReplica_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxModeCtlRxReplica_p1: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxModeCtlRxReplica_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxModeCtlRxReplica_p1 = uvm_reg_field::type_id::create("RxModeCtlRxReplica_p1",,get_full_name());
      this.RxModeCtlRxReplica_p1.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxModeCtlRxReplica_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxModeCtlRxReplica_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxGainCurrAdjRxReplica_p1 extends uvm_reg;
	rand uvm_reg_field RxGainCurrAdjRxReplica_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxGainCurrAdjRxReplica_p1: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxGainCurrAdjRxReplica_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxGainCurrAdjRxReplica_p1 = uvm_reg_field::type_id::create("RxGainCurrAdjRxReplica_p1",,get_full_name());
      this.RxGainCurrAdjRxReplica_p1.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxGainCurrAdjRxReplica_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxGainCurrAdjRxReplica_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxRxStandbyEn_p1 extends uvm_reg;
	rand uvm_reg_field DxRxStandbyEn_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DxRxStandbyEn_p1: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DxRxStandbyEn_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DxRxStandbyEn_p1 = uvm_reg_field::type_id::create("DxRxStandbyEn_p1",,get_full_name());
      this.DxRxStandbyEn_p1.configure(this, 1, 0, "RW", 0, 1'h1, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxRxStandbyEn_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxRxStandbyEn_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r0_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r0_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r0_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r0_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r0_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r0_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r0_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r0_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r0_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r0_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r0_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r0_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r0_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r0_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r0_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r0_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r0_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r0_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r0_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r0_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r0_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r0_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r0_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r0_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r0_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r0_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r0_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r0_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r0_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r0_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r0_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r0_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r0_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r0_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r0_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r0_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r0_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r0_p1",,get_full_name());
      this.TxDqDlyTg0_r0_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r0_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r0_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r0_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r0_p1",,get_full_name());
      this.TxDqDlyTg1_r0_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_SingleEndedMode_p1 extends uvm_reg;
	rand uvm_reg_field SingleEndedModeReserved;
	rand uvm_reg_field SingleEndedDQS;
	rand uvm_reg_field SingleEndedWCK;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   SingleEndedModeReserved: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   SingleEndedDQS: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   SingleEndedWCK: coverpoint {m_data[3:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_SingleEndedMode_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.SingleEndedModeReserved = uvm_reg_field::type_id::create("SingleEndedModeReserved",,get_full_name());
      this.SingleEndedModeReserved.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.SingleEndedDQS = uvm_reg_field::type_id::create("SingleEndedDQS",,get_full_name());
      this.SingleEndedDQS.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.SingleEndedWCK = uvm_reg_field::type_id::create("SingleEndedWCK",,get_full_name());
      this.SingleEndedWCK.configure(this, 2, 2, "RW", 0, 2'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_SingleEndedMode_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_SingleEndedMode_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxTrainPattern8BitMode_p1 extends uvm_reg;
	rand uvm_reg_field RxTrainPattern8BitMode_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxTrainPattern8BitMode_p1: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxTrainPattern8BitMode_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxTrainPattern8BitMode_p1 = uvm_reg_field::type_id::create("RxTrainPattern8BitMode_p1",,get_full_name());
      this.RxTrainPattern8BitMode_p1.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxTrainPattern8BitMode_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxTrainPattern8BitMode_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r0_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r0_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r0_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r0_p1",,get_full_name());
      this.DqRxVrefDac_r0_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbEn_p1 extends uvm_reg;
	rand uvm_reg_field EnStrblssRdMode;
	rand uvm_reg_field RxReplicaPowerDownNoRDQS;
	rand uvm_reg_field OdtDisDqs;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   EnStrblssRdMode: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxReplicaPowerDownNoRDQS: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   OdtDisDqs: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbEn_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.EnStrblssRdMode = uvm_reg_field::type_id::create("EnStrblssRdMode",,get_full_name());
      this.EnStrblssRdMode.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.RxReplicaPowerDownNoRDQS = uvm_reg_field::type_id::create("RxReplicaPowerDownNoRDQS",,get_full_name());
      this.RxReplicaPowerDownNoRDQS.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.OdtDisDqs = uvm_reg_field::type_id::create("OdtDisDqs",,get_full_name());
      this.OdtDisDqs.configure(this, 1, 2, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbEn_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbEn_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPipeEn_p1 extends uvm_reg;
	rand uvm_reg_field DxWrPipeEn;
	rand uvm_reg_field DxRdPipeEn;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DxWrPipeEn: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   DxRdPipeEn: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DxPipeEn_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DxWrPipeEn = uvm_reg_field::type_id::create("DxWrPipeEn",,get_full_name());
      this.DxWrPipeEn.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.DxRdPipeEn = uvm_reg_field::type_id::create("DxRdPipeEn",,get_full_name());
      this.DxRdPipeEn.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPipeEn_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPipeEn_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCDCtrl_p1 extends uvm_reg;
	rand uvm_reg_field PclkDCDEn;
	rand uvm_reg_field PclkDCDOffsetMode;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PclkDCDEn: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PclkDCDOffsetMode: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PclkDCDCtrl_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PclkDCDEn = uvm_reg_field::type_id::create("PclkDCDEn",,get_full_name());
      this.PclkDCDEn.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.PclkDCDOffsetMode = uvm_reg_field::type_id::create("PclkDCDOffsetMode",,get_full_name());
      this.PclkDCDOffsetMode.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCDCtrl_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCDCtrl_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PPTTrainSetup2_p1 extends uvm_reg;
	rand uvm_reg_field PPTTrainSetup2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PPTTrainSetup2_p1: coverpoint {m_data[10:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {12'b??????????00};
	      wildcard bins bit_0_wr_as_1 = {12'b??????????10};
	      wildcard bins bit_0_rd_as_0 = {12'b??????????01};
	      wildcard bins bit_0_rd_as_1 = {12'b??????????11};
	      wildcard bins bit_1_wr_as_0 = {12'b?????????0?0};
	      wildcard bins bit_1_wr_as_1 = {12'b?????????1?0};
	      wildcard bins bit_1_rd_as_0 = {12'b?????????0?1};
	      wildcard bins bit_1_rd_as_1 = {12'b?????????1?1};
	      wildcard bins bit_2_wr_as_0 = {12'b????????0??0};
	      wildcard bins bit_2_wr_as_1 = {12'b????????1??0};
	      wildcard bins bit_2_rd_as_0 = {12'b????????0??1};
	      wildcard bins bit_2_rd_as_1 = {12'b????????1??1};
	      wildcard bins bit_3_wr_as_0 = {12'b???????0???0};
	      wildcard bins bit_3_wr_as_1 = {12'b???????1???0};
	      wildcard bins bit_3_rd_as_0 = {12'b???????0???1};
	      wildcard bins bit_3_rd_as_1 = {12'b???????1???1};
	      wildcard bins bit_4_wr_as_0 = {12'b??????0????0};
	      wildcard bins bit_4_wr_as_1 = {12'b??????1????0};
	      wildcard bins bit_4_rd_as_0 = {12'b??????0????1};
	      wildcard bins bit_4_rd_as_1 = {12'b??????1????1};
	      wildcard bins bit_5_wr_as_0 = {12'b?????0?????0};
	      wildcard bins bit_5_wr_as_1 = {12'b?????1?????0};
	      wildcard bins bit_5_rd_as_0 = {12'b?????0?????1};
	      wildcard bins bit_5_rd_as_1 = {12'b?????1?????1};
	      wildcard bins bit_6_wr_as_0 = {12'b????0??????0};
	      wildcard bins bit_6_wr_as_1 = {12'b????1??????0};
	      wildcard bins bit_6_rd_as_0 = {12'b????0??????1};
	      wildcard bins bit_6_rd_as_1 = {12'b????1??????1};
	      wildcard bins bit_7_wr_as_0 = {12'b???0???????0};
	      wildcard bins bit_7_wr_as_1 = {12'b???1???????0};
	      wildcard bins bit_7_rd_as_0 = {12'b???0???????1};
	      wildcard bins bit_7_rd_as_1 = {12'b???1???????1};
	      wildcard bins bit_8_wr_as_0 = {12'b??0????????0};
	      wildcard bins bit_8_wr_as_1 = {12'b??1????????0};
	      wildcard bins bit_8_rd_as_0 = {12'b??0????????1};
	      wildcard bins bit_8_rd_as_1 = {12'b??1????????1};
	      wildcard bins bit_9_wr_as_0 = {12'b?0?????????0};
	      wildcard bins bit_9_wr_as_1 = {12'b?1?????????0};
	      wildcard bins bit_9_rd_as_0 = {12'b?0?????????1};
	      wildcard bins bit_9_rd_as_1 = {12'b?1?????????1};
	      wildcard bins bit_10_wr_as_0 = {12'b0??????????0};
	      wildcard bins bit_10_wr_as_1 = {12'b1??????????0};
	      wildcard bins bit_10_rd_as_0 = {12'b0??????????1};
	      wildcard bins bit_10_rd_as_1 = {12'b1??????????1};
	      option.weight = 44;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PPTTrainSetup2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PPTTrainSetup2_p1 = uvm_reg_field::type_id::create("PPTTrainSetup2_p1",,get_full_name());
      this.PPTTrainSetup2_p1.configure(this, 11, 0, "RW", 0, 11'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PPTTrainSetup2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PPTTrainSetup2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DMIPinPresent_p1 extends uvm_reg;
	rand uvm_reg_field RdDbiEnabled;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RdDbiEnabled: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DMIPinPresent_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RdDbiEnabled = uvm_reg_field::type_id::create("RdDbiEnabled",,get_full_name());
      this.RdDbiEnabled.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DMIPinPresent_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DMIPinPresent_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_InhibitTxRdPtrInit_p1 extends uvm_reg;
	rand uvm_reg_field InhibitTxRdPtrInit_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   InhibitTxRdPtrInit_p1: coverpoint {m_data[1:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_InhibitTxRdPtrInit_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.InhibitTxRdPtrInit_p1 = uvm_reg_field::type_id::create("InhibitTxRdPtrInit_p1",,get_full_name());
      this.InhibitTxRdPtrInit_p1.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_InhibitTxRdPtrInit_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_InhibitTxRdPtrInit_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r1_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r1_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r1_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r1_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r1_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r1_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r1_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r1_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r1_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r1_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r1_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r1_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r1_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r1_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r1_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r1_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RDqRDqsCntrl_p1 extends uvm_reg;
	rand uvm_reg_field RxPubLcdlSeed;
	rand uvm_reg_field RDqRDqsCntrl9;
	rand uvm_reg_field RxPubCalModeIs1UI;
	rand uvm_reg_field RxPubCntlByPState;
	rand uvm_reg_field RxPubRxReplicaCalModeIs1UI;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxPubLcdlSeed: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	   RDqRDqsCntrl9: coverpoint {m_data[9:9], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxPubCalModeIs1UI: coverpoint {m_data[10:10], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxPubCntlByPState: coverpoint {m_data[11:11], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxPubRxReplicaCalModeIs1UI: coverpoint {m_data[12:12], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RDqRDqsCntrl_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxPubLcdlSeed = uvm_reg_field::type_id::create("RxPubLcdlSeed",,get_full_name());
      this.RxPubLcdlSeed.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 0);
      this.RDqRDqsCntrl9 = uvm_reg_field::type_id::create("RDqRDqsCntrl9",,get_full_name());
      this.RDqRDqsCntrl9.configure(this, 1, 9, "RW", 0, 1'h0, 1, 0, 0);
      this.RxPubCalModeIs1UI = uvm_reg_field::type_id::create("RxPubCalModeIs1UI",,get_full_name());
      this.RxPubCalModeIs1UI.configure(this, 1, 10, "RW", 0, 1'h0, 1, 0, 0);
      this.RxPubCntlByPState = uvm_reg_field::type_id::create("RxPubCntlByPState",,get_full_name());
      this.RxPubCntlByPState.configure(this, 1, 11, "RW", 0, 1'h0, 1, 0, 0);
      this.RxPubRxReplicaCalModeIs1UI = uvm_reg_field::type_id::create("RxPubRxReplicaCalModeIs1UI",,get_full_name());
      this.RxPubRxReplicaCalModeIs1UI.configure(this, 1, 12, "RW", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RDqRDqsCntrl_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RDqRDqsCntrl_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r1_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r1_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r1_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r1_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r1_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r1_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r1_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r1_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r1_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r1_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r1_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r1_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r1_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r1_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r1_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r1_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r1_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r1_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r1_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r1_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r1_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r1_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r1_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r1_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r1_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r1_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r1_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r1_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r1_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r1_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r1_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r1_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r1_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r1_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r1_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r1_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r1_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r1_p1",,get_full_name());
      this.TxDqDlyTg0_r1_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r1_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r1_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r1_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r1_p1",,get_full_name());
      this.TxDqDlyTg1_r1_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r1_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r1_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r1_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r1_p1",,get_full_name());
      this.DqRxVrefDac_r1_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaRangeVal_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaShortCalRangeA;
	rand uvm_reg_field RxReplicaShortCalRangeB;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaShortCalRangeA: coverpoint {m_data[7:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd_as_0 = {9'b???????01};
	      wildcard bins bit_0_rd_as_1 = {9'b???????11};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd_as_0 = {9'b??????0?1};
	      wildcard bins bit_1_rd_as_1 = {9'b??????1?1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd_as_0 = {9'b?????0??1};
	      wildcard bins bit_2_rd_as_1 = {9'b?????1??1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd_as_0 = {9'b????0???1};
	      wildcard bins bit_3_rd_as_1 = {9'b????1???1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd_as_0 = {9'b???0????1};
	      wildcard bins bit_4_rd_as_1 = {9'b???1????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd_as_0 = {9'b??0?????1};
	      wildcard bins bit_5_rd_as_1 = {9'b??1?????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd_as_0 = {9'b?0??????1};
	      wildcard bins bit_6_rd_as_1 = {9'b?1??????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd_as_0 = {9'b0???????1};
	      wildcard bins bit_7_rd_as_1 = {9'b1???????1};
	      option.weight = 32;
	   }
	   RxReplicaShortCalRangeB: coverpoint {m_data[15:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd_as_0 = {9'b???????01};
	      wildcard bins bit_0_rd_as_1 = {9'b???????11};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd_as_0 = {9'b??????0?1};
	      wildcard bins bit_1_rd_as_1 = {9'b??????1?1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd_as_0 = {9'b?????0??1};
	      wildcard bins bit_2_rd_as_1 = {9'b?????1??1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd_as_0 = {9'b????0???1};
	      wildcard bins bit_3_rd_as_1 = {9'b????1???1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd_as_0 = {9'b???0????1};
	      wildcard bins bit_4_rd_as_1 = {9'b???1????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd_as_0 = {9'b??0?????1};
	      wildcard bins bit_5_rd_as_1 = {9'b??1?????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd_as_0 = {9'b?0??????1};
	      wildcard bins bit_6_rd_as_1 = {9'b?1??????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd_as_0 = {9'b0???????1};
	      wildcard bins bit_7_rd_as_1 = {9'b1???????1};
	      option.weight = 32;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaRangeVal_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaShortCalRangeA = uvm_reg_field::type_id::create("RxReplicaShortCalRangeA",,get_full_name());
      this.RxReplicaShortCalRangeA.configure(this, 8, 0, "RW", 0, 8'h4, 1, 0, 1);
      this.RxReplicaShortCalRangeB = uvm_reg_field::type_id::create("RxReplicaShortCalRangeB",,get_full_name());
      this.RxReplicaShortCalRangeB.configure(this, 8, 8, "RW", 0, 8'h4, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaRangeVal_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaRangeVal_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl04_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaTrackEn;
	rand uvm_reg_field RxReplicaLongCal;
	rand uvm_reg_field RxReplicaStride;
	rand uvm_reg_field RxReplicaStandby;
	rand uvm_reg_field RxReplicaPDenFSM;
	rand uvm_reg_field RxReplicaPDRecoverytime;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaTrackEn: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxReplicaLongCal: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxReplicaStride: coverpoint {m_data[5:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	   RxReplicaStandby: coverpoint {m_data[6:6], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxReplicaPDenFSM: coverpoint {m_data[7:7], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   RxReplicaPDRecoverytime: coverpoint {m_data[15:8], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {9'b???????00};
	      wildcard bins bit_0_wr_as_1 = {9'b???????10};
	      wildcard bins bit_0_rd_as_0 = {9'b???????01};
	      wildcard bins bit_0_rd_as_1 = {9'b???????11};
	      wildcard bins bit_1_wr_as_0 = {9'b??????0?0};
	      wildcard bins bit_1_wr_as_1 = {9'b??????1?0};
	      wildcard bins bit_1_rd_as_0 = {9'b??????0?1};
	      wildcard bins bit_1_rd_as_1 = {9'b??????1?1};
	      wildcard bins bit_2_wr_as_0 = {9'b?????0??0};
	      wildcard bins bit_2_wr_as_1 = {9'b?????1??0};
	      wildcard bins bit_2_rd_as_0 = {9'b?????0??1};
	      wildcard bins bit_2_rd_as_1 = {9'b?????1??1};
	      wildcard bins bit_3_wr_as_0 = {9'b????0???0};
	      wildcard bins bit_3_wr_as_1 = {9'b????1???0};
	      wildcard bins bit_3_rd_as_0 = {9'b????0???1};
	      wildcard bins bit_3_rd_as_1 = {9'b????1???1};
	      wildcard bins bit_4_wr_as_0 = {9'b???0????0};
	      wildcard bins bit_4_wr_as_1 = {9'b???1????0};
	      wildcard bins bit_4_rd_as_0 = {9'b???0????1};
	      wildcard bins bit_4_rd_as_1 = {9'b???1????1};
	      wildcard bins bit_5_wr_as_0 = {9'b??0?????0};
	      wildcard bins bit_5_wr_as_1 = {9'b??1?????0};
	      wildcard bins bit_5_rd_as_0 = {9'b??0?????1};
	      wildcard bins bit_5_rd_as_1 = {9'b??1?????1};
	      wildcard bins bit_6_wr_as_0 = {9'b?0??????0};
	      wildcard bins bit_6_wr_as_1 = {9'b?1??????0};
	      wildcard bins bit_6_rd_as_0 = {9'b?0??????1};
	      wildcard bins bit_6_rd_as_1 = {9'b?1??????1};
	      wildcard bins bit_7_wr_as_0 = {9'b0???????0};
	      wildcard bins bit_7_wr_as_1 = {9'b1???????0};
	      wildcard bins bit_7_rd_as_0 = {9'b0???????1};
	      wildcard bins bit_7_rd_as_1 = {9'b1???????1};
	      option.weight = 32;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl04_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaTrackEn = uvm_reg_field::type_id::create("RxReplicaTrackEn",,get_full_name());
      this.RxReplicaTrackEn.configure(this, 1, 0, "RW", 0, 1'h1, 1, 0, 0);
      this.RxReplicaLongCal = uvm_reg_field::type_id::create("RxReplicaLongCal",,get_full_name());
      this.RxReplicaLongCal.configure(this, 1, 1, "RW", 0, 1'h1, 1, 0, 0);
      this.RxReplicaStride = uvm_reg_field::type_id::create("RxReplicaStride",,get_full_name());
      this.RxReplicaStride.configure(this, 4, 2, "RW", 0, 4'h1, 1, 0, 0);
      this.RxReplicaStandby = uvm_reg_field::type_id::create("RxReplicaStandby",,get_full_name());
      this.RxReplicaStandby.configure(this, 1, 6, "RW", 0, 1'h0, 1, 0, 0);
      this.RxReplicaPDenFSM = uvm_reg_field::type_id::create("RxReplicaPDenFSM",,get_full_name());
      this.RxReplicaPDenFSM.configure(this, 1, 7, "RW", 0, 1'h0, 1, 0, 0);
      this.RxReplicaPDRecoverytime = uvm_reg_field::type_id::create("RxReplicaPDRecoverytime",,get_full_name());
      this.RxReplicaPDRecoverytime.configure(this, 8, 8, "RW", 0, 8'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl04_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl04_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r2_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r2_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r2_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r2_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r2_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r2_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r2_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r2_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r2_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r2_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r2_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r2_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r2_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r2_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r2_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r2_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r2_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r2_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r2_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r2_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r2_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r2_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r2_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r2_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r2_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r2_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r2_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r2_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r2_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r2_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r2_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r2_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r2_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r2_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r2_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r2_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r2_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r2_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r2_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r2_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r2_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r2_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r2_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r2_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r2_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r2_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r2_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r2_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r2_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r2_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r2_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r2_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r2_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r2_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r2_p1",,get_full_name());
      this.TxDqDlyTg0_r2_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r2_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r2_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r2_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r2_p1",,get_full_name());
      this.TxDqDlyTg1_r2_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase0_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaPathPhase0_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaPathPhase0_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase0_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaPathPhase0_p1 = uvm_reg_field::type_id::create("RxReplicaPathPhase0_p1",,get_full_name());
      this.RxReplicaPathPhase0_p1.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase0_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase0_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase1_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaPathPhase1_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaPathPhase1_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase1_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaPathPhase1_p1 = uvm_reg_field::type_id::create("RxReplicaPathPhase1_p1",,get_full_name());
      this.RxReplicaPathPhase1_p1.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase1_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase1_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase2_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaPathPhase2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaPathPhase2_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaPathPhase2_p1 = uvm_reg_field::type_id::create("RxReplicaPathPhase2_p1",,get_full_name());
      this.RxReplicaPathPhase2_p1.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase3_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaPathPhase3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaPathPhase3_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaPathPhase3_p1 = uvm_reg_field::type_id::create("RxReplicaPathPhase3_p1",,get_full_name());
      this.RxReplicaPathPhase3_p1.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase4_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaPathPhase4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaPathPhase4_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaPathPhase4_p1 = uvm_reg_field::type_id::create("RxReplicaPathPhase4_p1",,get_full_name());
      this.RxReplicaPathPhase4_p1.configure(this, 9, 0, "RW", 0, 9'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl01_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaSelPathPhase;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaSelPathPhase: coverpoint {m_data[2:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {4'b??00};
	      wildcard bins bit_0_wr_as_1 = {4'b??10};
	      wildcard bins bit_0_rd_as_0 = {4'b??01};
	      wildcard bins bit_0_rd_as_1 = {4'b??11};
	      wildcard bins bit_1_wr_as_0 = {4'b?0?0};
	      wildcard bins bit_1_wr_as_1 = {4'b?1?0};
	      wildcard bins bit_1_rd_as_0 = {4'b?0?1};
	      wildcard bins bit_1_rd_as_1 = {4'b?1?1};
	      wildcard bins bit_2_wr_as_0 = {4'b0??0};
	      wildcard bins bit_2_wr_as_1 = {4'b1??0};
	      wildcard bins bit_2_rd_as_0 = {4'b0??1};
	      wildcard bins bit_2_rd_as_1 = {4'b1??1};
	      option.weight = 12;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl01_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaSelPathPhase = uvm_reg_field::type_id::create("RxReplicaSelPathPhase",,get_full_name());
      this.RxReplicaSelPathPhase.configure(this, 3, 0, "RW", 0, 3'h2, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl01_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl01_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl02_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaDiffLimit;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaDiffLimit: coverpoint {m_data[6:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl02_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaDiffLimit = uvm_reg_field::type_id::create("RxReplicaDiffLimit",,get_full_name());
      this.RxReplicaDiffLimit.configure(this, 7, 0, "RW", 0, 7'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl02_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl02_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl03_p1 extends uvm_reg;
	rand uvm_reg_field RxReplicaRatioTrn;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxReplicaRatioTrn: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl03_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxReplicaRatioTrn = uvm_reg_field::type_id::create("RxReplicaRatioTrn",,get_full_name());
      this.RxReplicaRatioTrn.configure(this, 10, 0, "RW", 0, 10'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl03_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl03_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r2_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r2_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r2_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r2_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r2_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r2_p1",,get_full_name());
      this.DqRxVrefDac_r2_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r2_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r2_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r3_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r3_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r3_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r3_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r3_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r3_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r3_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r3_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r3_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r3_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r3_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r3_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r3_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r3_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r3_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r3_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r3_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r3_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r3_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r3_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r3_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r3_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r3_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r3_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r3_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r3_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r3_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r3_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r3_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r3_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r3_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r3_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r3_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r3_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r3_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r3_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r3_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r3_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r3_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r3_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r3_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r3_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r3_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r3_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r3_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r3_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r3_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r3_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r3_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r3_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r3_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r3_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r3_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r3_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r3_p1",,get_full_name());
      this.TxDqDlyTg0_r3_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r3_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r3_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r3_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r3_p1",,get_full_name());
      this.TxDqDlyTg1_r3_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r3_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r3_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r3_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r3_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r3_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r3_p1",,get_full_name());
      this.DqRxVrefDac_r3_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r3_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r3_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r4_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r4_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r4_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r4_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r4_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r4_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r4_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r4_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r4_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r4_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r4_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r4_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r4_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r4_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r4_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r4_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r4_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r4_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r4_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r4_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r4_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r4_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r4_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r4_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r4_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r4_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r4_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r4_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r4_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r4_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r4_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r4_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r4_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r4_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r4_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r4_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r4_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r4_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r4_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r4_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r4_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r4_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r4_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r4_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r4_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r4_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r4_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r4_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r4_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r4_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r4_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r4_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r4_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r4_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r4_p1",,get_full_name());
      this.TxDqDlyTg0_r4_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r4_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r4_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r4_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r4_p1",,get_full_name());
      this.TxDqDlyTg1_r4_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r4_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r4_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r4_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r4_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r4_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r4_p1",,get_full_name());
      this.DqRxVrefDac_r4_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r4_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r4_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r5_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r5_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r5_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r5_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r5_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r5_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r5_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r5_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r5_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r5_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r5_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r5_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r5_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r5_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r5_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r5_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r5_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r5_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r5_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r5_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r5_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r5_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r5_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r5_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r5_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r5_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r5_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r5_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r5_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r5_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r5_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r5_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r5_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r5_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r5_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r5_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r5_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r5_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r5_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r5_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r5_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r5_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r5_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r5_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r5_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r5_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r5_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r5_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r5_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r5_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r5_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r5_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r5_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r5_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r5_p1",,get_full_name());
      this.TxDqDlyTg0_r5_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r5_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r5_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r5_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r5_p1",,get_full_name());
      this.TxDqDlyTg1_r5_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r5_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r5_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r5_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r5_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r5_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r5_p1",,get_full_name());
      this.DqRxVrefDac_r5_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r5_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r5_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r6_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r6_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r6_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r6_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r6_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r6_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r6_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r6_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r6_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r6_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r6_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r6_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r6_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r6_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r6_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r6_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r6_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r6_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r6_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r6_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r6_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r6_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r6_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r6_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r6_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r6_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r6_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r6_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r6_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r6_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r6_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r6_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r6_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r6_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r6_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r6_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r6_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r6_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r6_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r6_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r6_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r6_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r6_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r6_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r6_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r6_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r6_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r6_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r6_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r6_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r6_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r6_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r6_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r6_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r6_p1",,get_full_name());
      this.TxDqDlyTg0_r6_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r6_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r6_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r6_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r6_p1",,get_full_name());
      this.TxDqDlyTg1_r6_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r6_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r6_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r6_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r6_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r6_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r6_p1",,get_full_name());
      this.DqRxVrefDac_r6_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r6_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r6_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r7_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r7_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r7_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r7_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r7_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r7_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r7_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r7_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r7_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r7_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r7_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r7_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r7_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r7_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r7_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r7_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r7_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r7_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r7_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r7_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r7_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r7_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r7_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r7_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r7_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r7_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r7_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r7_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r7_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r7_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r7_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r7_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r7_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r7_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r7_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r7_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r7_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r7_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r7_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r7_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r7_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r7_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r7_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r7_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r7_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r7_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r7_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r7_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r7_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r7_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r7_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r7_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r7_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r7_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r7_p1",,get_full_name());
      this.TxDqDlyTg0_r7_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r7_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r7_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r7_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r7_p1",,get_full_name());
      this.TxDqDlyTg1_r7_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r7_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r7_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r7_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r7_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r7_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r7_p1",,get_full_name());
      this.DqRxVrefDac_r7_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r7_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r7_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl0DB_p1 extends uvm_reg;
	rand uvm_reg_field PclkDCACalModeDB;
	rand uvm_reg_field PclkDCAEnDB;
	rand uvm_reg_field PclkDCATxLcdlPhSelDB;
	rand uvm_reg_field PclkDCDSettleDB;
	rand uvm_reg_field PclkDCDSampTimeDB;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PclkDCACalModeDB: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PclkDCAEnDB: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PclkDCATxLcdlPhSelDB: coverpoint {m_data[3:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {3'b?00};
	      wildcard bins bit_0_wr_as_1 = {3'b?10};
	      wildcard bins bit_0_rd_as_0 = {3'b?01};
	      wildcard bins bit_0_rd_as_1 = {3'b?11};
	      wildcard bins bit_1_wr_as_0 = {3'b0?0};
	      wildcard bins bit_1_wr_as_1 = {3'b1?0};
	      wildcard bins bit_1_rd_as_0 = {3'b0?1};
	      wildcard bins bit_1_rd_as_1 = {3'b1?1};
	      option.weight = 8;
	   }
	   PclkDCDSettleDB: coverpoint {m_data[10:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	   PclkDCDSampTimeDB: coverpoint {m_data[14:11], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl0DB_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PclkDCACalModeDB = uvm_reg_field::type_id::create("PclkDCACalModeDB",,get_full_name());
      this.PclkDCACalModeDB.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.PclkDCAEnDB = uvm_reg_field::type_id::create("PclkDCAEnDB",,get_full_name());
      this.PclkDCAEnDB.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.PclkDCATxLcdlPhSelDB = uvm_reg_field::type_id::create("PclkDCATxLcdlPhSelDB",,get_full_name());
      this.PclkDCATxLcdlPhSelDB.configure(this, 2, 2, "RW", 0, 2'h0, 1, 0, 0);
      this.PclkDCDSettleDB = uvm_reg_field::type_id::create("PclkDCDSettleDB",,get_full_name());
      this.PclkDCDSettleDB.configure(this, 7, 4, "RW", 0, 7'h4, 1, 0, 0);
      this.PclkDCDSampTimeDB = uvm_reg_field::type_id::create("PclkDCDSampTimeDB",,get_full_name());
      this.PclkDCDSampTimeDB.configure(this, 4, 11, "RW", 0, 4'h2, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl0DB_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl0DB_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCASampDelayLCDLDB_p1 extends uvm_reg;
	rand uvm_reg_field PclkDCASampDelayLCDLDB_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PclkDCASampDelayLCDLDB_p1: coverpoint {m_data[3:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {5'b???00};
	      wildcard bins bit_0_wr_as_1 = {5'b???10};
	      wildcard bins bit_0_rd_as_0 = {5'b???01};
	      wildcard bins bit_0_rd_as_1 = {5'b???11};
	      wildcard bins bit_1_wr_as_0 = {5'b??0?0};
	      wildcard bins bit_1_wr_as_1 = {5'b??1?0};
	      wildcard bins bit_1_rd_as_0 = {5'b??0?1};
	      wildcard bins bit_1_rd_as_1 = {5'b??1?1};
	      wildcard bins bit_2_wr_as_0 = {5'b?0??0};
	      wildcard bins bit_2_wr_as_1 = {5'b?1??0};
	      wildcard bins bit_2_rd_as_0 = {5'b?0??1};
	      wildcard bins bit_2_rd_as_1 = {5'b?1??1};
	      wildcard bins bit_3_wr_as_0 = {5'b0???0};
	      wildcard bins bit_3_wr_as_1 = {5'b1???0};
	      wildcard bins bit_3_rd_as_0 = {5'b0???1};
	      wildcard bins bit_3_rd_as_1 = {5'b1???1};
	      option.weight = 16;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PclkDCASampDelayLCDLDB_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PclkDCASampDelayLCDLDB_p1 = uvm_reg_field::type_id::create("PclkDCASampDelayLCDLDB_p1",,get_full_name());
      this.PclkDCASampDelayLCDLDB_p1.configure(this, 4, 0, "RW", 0, 4'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCASampDelayLCDLDB_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCASampDelayLCDLDB_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg0_r8_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg0_r8_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg0_r8_p1",,get_full_name());
      this.RxClkT2UIDlyTg0_r8_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkT2UIDlyTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkT2UIDlyTg1_r8_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkT2UIDlyTg1_r8_p1 = uvm_reg_field::type_id::create("RxClkT2UIDlyTg1_r8_p1",,get_full_name());
      this.RxClkT2UIDlyTg1_r8_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg0_r8_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg0_r8_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg0_r8_p1",,get_full_name());
      this.RxClkC2UIDlyTg0_r8_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkC2UIDlyTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkC2UIDlyTg1_r8_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkC2UIDlyTg1_r8_p1 = uvm_reg_field::type_id::create("RxClkC2UIDlyTg1_r8_p1",,get_full_name());
      this.RxClkC2UIDlyTg1_r8_p1.configure(this, 10, 0, "RW", 0, 10'h110, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg0_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg0_r8_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg0_r8_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg0_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqLeftEyeOffsetTg1_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqLeftEyeOffsetTg1_r8_p1 = uvm_reg_field::type_id::create("TxDqLeftEyeOffsetTg1_r8_p1",,get_full_name());
      this.TxDqLeftEyeOffsetTg1_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg0_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg0_r8_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg0_r8_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg0_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqRightEyeOffsetTg1_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqRightEyeOffsetTg1_r8_p1 = uvm_reg_field::type_id::create("TxDqRightEyeOffsetTg1_r8_p1",,get_full_name());
      this.TxDqRightEyeOffsetTg1_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg0_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg0_r8_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg0_r8_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg0_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTLeftEyeOffsetTg1_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTLeftEyeOffsetTg1_r8_p1 = uvm_reg_field::type_id::create("RxClkTLeftEyeOffsetTg1_r8_p1",,get_full_name());
      this.RxClkTLeftEyeOffsetTg1_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg0_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg0_r8_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg0_r8_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg0_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkTRightEyeOffsetTg1_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkTRightEyeOffsetTg1_r8_p1 = uvm_reg_field::type_id::create("RxClkTRightEyeOffsetTg1_r8_p1",,get_full_name());
      this.RxClkTRightEyeOffsetTg1_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg0_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg0_r8_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg0_r8_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg0_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCLeftEyeOffsetTg1_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCLeftEyeOffsetTg1_r8_p1 = uvm_reg_field::type_id::create("RxClkCLeftEyeOffsetTg1_r8_p1",,get_full_name());
      this.RxClkCLeftEyeOffsetTg1_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg0_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg0_r8_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg0_r8_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg0_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxClkCRightEyeOffsetTg1_r8_p1: coverpoint {m_data[5:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {7'b?????00};
	      wildcard bins bit_0_wr_as_1 = {7'b?????10};
	      wildcard bins bit_0_rd_as_0 = {7'b?????01};
	      wildcard bins bit_0_rd_as_1 = {7'b?????11};
	      wildcard bins bit_1_wr_as_0 = {7'b????0?0};
	      wildcard bins bit_1_wr_as_1 = {7'b????1?0};
	      wildcard bins bit_1_rd_as_0 = {7'b????0?1};
	      wildcard bins bit_1_rd_as_1 = {7'b????1?1};
	      wildcard bins bit_2_wr_as_0 = {7'b???0??0};
	      wildcard bins bit_2_wr_as_1 = {7'b???1??0};
	      wildcard bins bit_2_rd_as_0 = {7'b???0??1};
	      wildcard bins bit_2_rd_as_1 = {7'b???1??1};
	      wildcard bins bit_3_wr_as_0 = {7'b??0???0};
	      wildcard bins bit_3_wr_as_1 = {7'b??1???0};
	      wildcard bins bit_3_rd_as_0 = {7'b??0???1};
	      wildcard bins bit_3_rd_as_1 = {7'b??1???1};
	      wildcard bins bit_4_wr_as_0 = {7'b?0????0};
	      wildcard bins bit_4_wr_as_1 = {7'b?1????0};
	      wildcard bins bit_4_rd_as_0 = {7'b?0????1};
	      wildcard bins bit_4_rd_as_1 = {7'b?1????1};
	      wildcard bins bit_5_wr_as_0 = {7'b0?????0};
	      wildcard bins bit_5_wr_as_1 = {7'b1?????0};
	      wildcard bins bit_5_rd_as_0 = {7'b0?????1};
	      wildcard bins bit_5_rd_as_1 = {7'b1?????1};
	      option.weight = 24;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r8_p1");
		super.new(name, 8,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxClkCRightEyeOffsetTg1_r8_p1 = uvm_reg_field::type_id::create("RxClkCRightEyeOffsetTg1_r8_p1",,get_full_name());
      this.RxClkCRightEyeOffsetTg1_r8_p1.configure(this, 6, 0, "RW", 0, 6'h1f, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg0_r8_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg0_r8_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg0_r8_p1",,get_full_name());
      this.RxDigStrbDlyTg0_r8_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field RxDigStrbDlyTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   RxDigStrbDlyTg1_r8_p1: coverpoint {m_data[11:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {13'b???????????00};
	      wildcard bins bit_0_wr_as_1 = {13'b???????????10};
	      wildcard bins bit_0_rd_as_0 = {13'b???????????01};
	      wildcard bins bit_0_rd_as_1 = {13'b???????????11};
	      wildcard bins bit_1_wr_as_0 = {13'b??????????0?0};
	      wildcard bins bit_1_wr_as_1 = {13'b??????????1?0};
	      wildcard bins bit_1_rd_as_0 = {13'b??????????0?1};
	      wildcard bins bit_1_rd_as_1 = {13'b??????????1?1};
	      wildcard bins bit_2_wr_as_0 = {13'b?????????0??0};
	      wildcard bins bit_2_wr_as_1 = {13'b?????????1??0};
	      wildcard bins bit_2_rd_as_0 = {13'b?????????0??1};
	      wildcard bins bit_2_rd_as_1 = {13'b?????????1??1};
	      wildcard bins bit_3_wr_as_0 = {13'b????????0???0};
	      wildcard bins bit_3_wr_as_1 = {13'b????????1???0};
	      wildcard bins bit_3_rd_as_0 = {13'b????????0???1};
	      wildcard bins bit_3_rd_as_1 = {13'b????????1???1};
	      wildcard bins bit_4_wr_as_0 = {13'b???????0????0};
	      wildcard bins bit_4_wr_as_1 = {13'b???????1????0};
	      wildcard bins bit_4_rd_as_0 = {13'b???????0????1};
	      wildcard bins bit_4_rd_as_1 = {13'b???????1????1};
	      wildcard bins bit_5_wr_as_0 = {13'b??????0?????0};
	      wildcard bins bit_5_wr_as_1 = {13'b??????1?????0};
	      wildcard bins bit_5_rd_as_0 = {13'b??????0?????1};
	      wildcard bins bit_5_rd_as_1 = {13'b??????1?????1};
	      wildcard bins bit_6_wr_as_0 = {13'b?????0??????0};
	      wildcard bins bit_6_wr_as_1 = {13'b?????1??????0};
	      wildcard bins bit_6_rd_as_0 = {13'b?????0??????1};
	      wildcard bins bit_6_rd_as_1 = {13'b?????1??????1};
	      wildcard bins bit_7_wr_as_0 = {13'b????0???????0};
	      wildcard bins bit_7_wr_as_1 = {13'b????1???????0};
	      wildcard bins bit_7_rd_as_0 = {13'b????0???????1};
	      wildcard bins bit_7_rd_as_1 = {13'b????1???????1};
	      wildcard bins bit_8_wr_as_0 = {13'b???0????????0};
	      wildcard bins bit_8_wr_as_1 = {13'b???1????????0};
	      wildcard bins bit_8_rd_as_0 = {13'b???0????????1};
	      wildcard bins bit_8_rd_as_1 = {13'b???1????????1};
	      wildcard bins bit_9_wr_as_0 = {13'b??0?????????0};
	      wildcard bins bit_9_wr_as_1 = {13'b??1?????????0};
	      wildcard bins bit_9_rd_as_0 = {13'b??0?????????1};
	      wildcard bins bit_9_rd_as_1 = {13'b??1?????????1};
	      wildcard bins bit_10_wr_as_0 = {13'b?0??????????0};
	      wildcard bins bit_10_wr_as_1 = {13'b?1??????????0};
	      wildcard bins bit_10_rd_as_0 = {13'b?0??????????1};
	      wildcard bins bit_10_rd_as_1 = {13'b?1??????????1};
	      wildcard bins bit_11_wr_as_0 = {13'b0???????????0};
	      wildcard bins bit_11_wr_as_1 = {13'b1???????????0};
	      wildcard bins bit_11_rd_as_0 = {13'b0???????????1};
	      wildcard bins bit_11_rd_as_1 = {13'b1???????????1};
	      option.weight = 48;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.RxDigStrbDlyTg1_r8_p1 = uvm_reg_field::type_id::create("RxDigStrbDlyTg1_r8_p1",,get_full_name());
      this.RxDigStrbDlyTg1_r8_p1.configure(this, 12, 0, "RW", 0, 12'h100, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r8_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg0_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg0_r8_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg0_r8_p1 = uvm_reg_field::type_id::create("TxDqDlyTg0_r8_p1",,get_full_name());
      this.TxDqDlyTg0_r8_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r8_p1 extends uvm_reg;
	rand uvm_reg_field TxDqDlyTg1_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   TxDqDlyTg1_r8_p1: coverpoint {m_data[9:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {11'b?????????00};
	      wildcard bins bit_0_wr_as_1 = {11'b?????????10};
	      wildcard bins bit_0_rd_as_0 = {11'b?????????01};
	      wildcard bins bit_0_rd_as_1 = {11'b?????????11};
	      wildcard bins bit_1_wr_as_0 = {11'b????????0?0};
	      wildcard bins bit_1_wr_as_1 = {11'b????????1?0};
	      wildcard bins bit_1_rd_as_0 = {11'b????????0?1};
	      wildcard bins bit_1_rd_as_1 = {11'b????????1?1};
	      wildcard bins bit_2_wr_as_0 = {11'b???????0??0};
	      wildcard bins bit_2_wr_as_1 = {11'b???????1??0};
	      wildcard bins bit_2_rd_as_0 = {11'b???????0??1};
	      wildcard bins bit_2_rd_as_1 = {11'b???????1??1};
	      wildcard bins bit_3_wr_as_0 = {11'b??????0???0};
	      wildcard bins bit_3_wr_as_1 = {11'b??????1???0};
	      wildcard bins bit_3_rd_as_0 = {11'b??????0???1};
	      wildcard bins bit_3_rd_as_1 = {11'b??????1???1};
	      wildcard bins bit_4_wr_as_0 = {11'b?????0????0};
	      wildcard bins bit_4_wr_as_1 = {11'b?????1????0};
	      wildcard bins bit_4_rd_as_0 = {11'b?????0????1};
	      wildcard bins bit_4_rd_as_1 = {11'b?????1????1};
	      wildcard bins bit_5_wr_as_0 = {11'b????0?????0};
	      wildcard bins bit_5_wr_as_1 = {11'b????1?????0};
	      wildcard bins bit_5_rd_as_0 = {11'b????0?????1};
	      wildcard bins bit_5_rd_as_1 = {11'b????1?????1};
	      wildcard bins bit_6_wr_as_0 = {11'b???0??????0};
	      wildcard bins bit_6_wr_as_1 = {11'b???1??????0};
	      wildcard bins bit_6_rd_as_0 = {11'b???0??????1};
	      wildcard bins bit_6_rd_as_1 = {11'b???1??????1};
	      wildcard bins bit_7_wr_as_0 = {11'b??0???????0};
	      wildcard bins bit_7_wr_as_1 = {11'b??1???????0};
	      wildcard bins bit_7_rd_as_0 = {11'b??0???????1};
	      wildcard bins bit_7_rd_as_1 = {11'b??1???????1};
	      wildcard bins bit_8_wr_as_0 = {11'b?0????????0};
	      wildcard bins bit_8_wr_as_1 = {11'b?1????????0};
	      wildcard bins bit_8_rd_as_0 = {11'b?0????????1};
	      wildcard bins bit_8_rd_as_1 = {11'b?1????????1};
	      wildcard bins bit_9_wr_as_0 = {11'b0?????????0};
	      wildcard bins bit_9_wr_as_1 = {11'b1?????????0};
	      wildcard bins bit_9_rd_as_0 = {11'b0?????????1};
	      wildcard bins bit_9_rd_as_1 = {11'b1?????????1};
	      option.weight = 40;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.TxDqDlyTg1_r8_p1 = uvm_reg_field::type_id::create("TxDqDlyTg1_r8_p1",,get_full_name());
      this.TxDqDlyTg1_r8_p1.configure(this, 10, 0, "RW", 0, 10'h20, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r8_p1 extends uvm_reg;
	rand uvm_reg_field DqRxVrefDac_r8_p1;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   DqRxVrefDac_r8_p1: coverpoint {m_data[8:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {10'b????????00};
	      wildcard bins bit_0_wr_as_1 = {10'b????????10};
	      wildcard bins bit_0_rd_as_0 = {10'b????????01};
	      wildcard bins bit_0_rd_as_1 = {10'b????????11};
	      wildcard bins bit_1_wr_as_0 = {10'b???????0?0};
	      wildcard bins bit_1_wr_as_1 = {10'b???????1?0};
	      wildcard bins bit_1_rd_as_0 = {10'b???????0?1};
	      wildcard bins bit_1_rd_as_1 = {10'b???????1?1};
	      wildcard bins bit_2_wr_as_0 = {10'b??????0??0};
	      wildcard bins bit_2_wr_as_1 = {10'b??????1??0};
	      wildcard bins bit_2_rd_as_0 = {10'b??????0??1};
	      wildcard bins bit_2_rd_as_1 = {10'b??????1??1};
	      wildcard bins bit_3_wr_as_0 = {10'b?????0???0};
	      wildcard bins bit_3_wr_as_1 = {10'b?????1???0};
	      wildcard bins bit_3_rd_as_0 = {10'b?????0???1};
	      wildcard bins bit_3_rd_as_1 = {10'b?????1???1};
	      wildcard bins bit_4_wr_as_0 = {10'b????0????0};
	      wildcard bins bit_4_wr_as_1 = {10'b????1????0};
	      wildcard bins bit_4_rd_as_0 = {10'b????0????1};
	      wildcard bins bit_4_rd_as_1 = {10'b????1????1};
	      wildcard bins bit_5_wr_as_0 = {10'b???0?????0};
	      wildcard bins bit_5_wr_as_1 = {10'b???1?????0};
	      wildcard bins bit_5_rd_as_0 = {10'b???0?????1};
	      wildcard bins bit_5_rd_as_1 = {10'b???1?????1};
	      wildcard bins bit_6_wr_as_0 = {10'b??0??????0};
	      wildcard bins bit_6_wr_as_1 = {10'b??1??????0};
	      wildcard bins bit_6_rd_as_0 = {10'b??0??????1};
	      wildcard bins bit_6_rd_as_1 = {10'b??1??????1};
	      wildcard bins bit_7_wr_as_0 = {10'b?0???????0};
	      wildcard bins bit_7_wr_as_1 = {10'b?1???????0};
	      wildcard bins bit_7_rd_as_0 = {10'b?0???????1};
	      wildcard bins bit_7_rd_as_1 = {10'b?1???????1};
	      wildcard bins bit_8_wr_as_0 = {10'b0????????0};
	      wildcard bins bit_8_wr_as_1 = {10'b1????????0};
	      wildcard bins bit_8_rd_as_0 = {10'b0????????1};
	      wildcard bins bit_8_rd_as_1 = {10'b1????????1};
	      option.weight = 36;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r8_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.DqRxVrefDac_r8_p1 = uvm_reg_field::type_id::create("DqRxVrefDac_r8_p1",,get_full_name());
      this.DqRxVrefDac_r8_p1.configure(this, 9, 0, "RW", 0, 9'hff, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r8_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r8_p1


class ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl1DB_p1 extends uvm_reg;
	rand uvm_reg_field PclkDCAInvertSampDB;
	rand uvm_reg_field PclkDCALcdlEn4pDB;
	rand uvm_reg_field PclkDCDMissionModeDelayDB;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   PclkDCAInvertSampDB: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PclkDCALcdlEn4pDB: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   PclkDCDMissionModeDelayDB: coverpoint {m_data[8:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {8'b??????00};
	      wildcard bins bit_0_wr_as_1 = {8'b??????10};
	      wildcard bins bit_0_rd_as_0 = {8'b??????01};
	      wildcard bins bit_0_rd_as_1 = {8'b??????11};
	      wildcard bins bit_1_wr_as_0 = {8'b?????0?0};
	      wildcard bins bit_1_wr_as_1 = {8'b?????1?0};
	      wildcard bins bit_1_rd_as_0 = {8'b?????0?1};
	      wildcard bins bit_1_rd_as_1 = {8'b?????1?1};
	      wildcard bins bit_2_wr_as_0 = {8'b????0??0};
	      wildcard bins bit_2_wr_as_1 = {8'b????1??0};
	      wildcard bins bit_2_rd_as_0 = {8'b????0??1};
	      wildcard bins bit_2_rd_as_1 = {8'b????1??1};
	      wildcard bins bit_3_wr_as_0 = {8'b???0???0};
	      wildcard bins bit_3_wr_as_1 = {8'b???1???0};
	      wildcard bins bit_3_rd_as_0 = {8'b???0???1};
	      wildcard bins bit_3_rd_as_1 = {8'b???1???1};
	      wildcard bins bit_4_wr_as_0 = {8'b??0????0};
	      wildcard bins bit_4_wr_as_1 = {8'b??1????0};
	      wildcard bins bit_4_rd_as_0 = {8'b??0????1};
	      wildcard bins bit_4_rd_as_1 = {8'b??1????1};
	      wildcard bins bit_5_wr_as_0 = {8'b?0?????0};
	      wildcard bins bit_5_wr_as_1 = {8'b?1?????0};
	      wildcard bins bit_5_rd_as_0 = {8'b?0?????1};
	      wildcard bins bit_5_rd_as_1 = {8'b?1?????1};
	      wildcard bins bit_6_wr_as_0 = {8'b0??????0};
	      wildcard bins bit_6_wr_as_1 = {8'b1??????0};
	      wildcard bins bit_6_rd_as_0 = {8'b0??????1};
	      wildcard bins bit_6_rd_as_1 = {8'b1??????1};
	      option.weight = 28;
	   }
	endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl1DB_p1");
		super.new(name, 16,build_coverage(UVM_NO_COVERAGE));
		add_coverage(build_coverage(UVM_NO_COVERAGE));
		if (has_coverage(UVM_CVR_ALL))
			cg_bits = new();
	endfunction: new
   virtual function void build();
      this.PclkDCAInvertSampDB = uvm_reg_field::type_id::create("PclkDCAInvertSampDB",,get_full_name());
      this.PclkDCAInvertSampDB.configure(this, 1, 0, "RW", 0, 1'h0, 1, 0, 0);
      this.PclkDCALcdlEn4pDB = uvm_reg_field::type_id::create("PclkDCALcdlEn4pDB",,get_full_name());
      this.PclkDCALcdlEn4pDB.configure(this, 1, 1, "RW", 0, 1'h0, 1, 0, 0);
      this.PclkDCDMissionModeDelayDB = uvm_reg_field::type_id::create("PclkDCDMissionModeDelayDB",,get_full_name());
      this.PclkDCDMissionModeDelayDB.configure(this, 7, 2, "RW", 0, 7'h4, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl1DB_p1)

`ifdef UVM_REG_PROTECTED_SAMPLE
    	 protected virtual function void sample(uvm_reg_data_t data,
    	                             uvm_reg_data_t byte_en,
    	                             bit            is_read,
    	                             uvm_reg_map    map);
`else
	 virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
`endif
	   if (get_coverage(UVM_CVR_ALL)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction
endclass : ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl1DB_p1


class ral_block_DWC_DDRPHYA_DBYTE3_p1 extends uvm_reg_block;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DFIMRL_p1 DFIMRL_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_EnableWriteLinkEcc_p1 EnableWriteLinkEcc_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxDfiClkDis_p1 DxDfiClkDis_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPClkDis_p1 DxPClkDis_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_LP5DfiDataEnLatency_p1 LP5DfiDataEnLatency_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg0_p1 PptDqsCntInvTrnTg0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg1_p1 PptDqsCntInvTrnTg1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TrackingModeCntrl_p1 TrackingModeCntrl_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r0_p1 RxClkT2UIDlyTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r0_p1 RxClkT2UIDlyTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r0_p1 RxClkC2UIDlyTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r0_p1 RxClkC2UIDlyTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg0_p1 PptWck2DqoCntInvTrnTg0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg1_p1 PptWck2DqoCntInvTrnTg1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg0_p1 TxDqsLeftEyeOffsetTg0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg1_p1 TxDqsLeftEyeOffsetTg1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg0_p1 RxEnDlyTg0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg1_p1 RxEnDlyTg1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg0_p1 TxDqsRightEyeOffsetTg0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg1_p1 TxDqsRightEyeOffsetTg1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqsPreambleControl_p1 DqsPreambleControl_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DbyteRxDqsModeCntrl_p1 DbyteRxDqsModeCntrl_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCntl1_p1 RxClkCntl1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg0_p1 TxDqsDlyTg0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg1_p1 TxDqsDlyTg1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg0_p1 TxWckDlyTg0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg1_p1 TxWckDlyTg1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxModeCtlRxReplica_p1 RxModeCtlRxReplica_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxGainCurrAdjRxReplica_p1 RxGainCurrAdjRxReplica_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxRxStandbyEn_p1 DxRxStandbyEn_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r0_p1 TxDqLeftEyeOffsetTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r0_p1 TxDqLeftEyeOffsetTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r0_p1 TxDqRightEyeOffsetTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r0_p1 TxDqRightEyeOffsetTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r0_p1 RxClkTLeftEyeOffsetTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r0_p1 RxClkTLeftEyeOffsetTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r0_p1 RxClkTRightEyeOffsetTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r0_p1 RxClkTRightEyeOffsetTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r0_p1 RxClkCLeftEyeOffsetTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r0_p1 RxClkCLeftEyeOffsetTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r0_p1 RxClkCRightEyeOffsetTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r0_p1 RxClkCRightEyeOffsetTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r0_p1 RxDigStrbDlyTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r0_p1 RxDigStrbDlyTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r0_p1 TxDqDlyTg0_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r0_p1 TxDqDlyTg1_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_SingleEndedMode_p1 SingleEndedMode_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxTrainPattern8BitMode_p1 RxTrainPattern8BitMode_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r0_p1 DqRxVrefDac_r0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbEn_p1 RxDigStrbEn_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPipeEn_p1 DxPipeEn_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCDCtrl_p1 PclkDCDCtrl_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PPTTrainSetup2_p1 PPTTrainSetup2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DMIPinPresent_p1 DMIPinPresent_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_InhibitTxRdPtrInit_p1 InhibitTxRdPtrInit_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r1_p1 RxClkT2UIDlyTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r1_p1 RxClkT2UIDlyTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r1_p1 RxClkC2UIDlyTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r1_p1 RxClkC2UIDlyTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RDqRDqsCntrl_p1 RDqRDqsCntrl_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r1_p1 TxDqLeftEyeOffsetTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r1_p1 TxDqLeftEyeOffsetTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r1_p1 TxDqRightEyeOffsetTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r1_p1 TxDqRightEyeOffsetTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r1_p1 RxClkTLeftEyeOffsetTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r1_p1 RxClkTLeftEyeOffsetTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r1_p1 RxClkTRightEyeOffsetTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r1_p1 RxClkTRightEyeOffsetTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r1_p1 RxClkCLeftEyeOffsetTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r1_p1 RxClkCLeftEyeOffsetTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r1_p1 RxClkCRightEyeOffsetTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r1_p1 RxClkCRightEyeOffsetTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r1_p1 RxDigStrbDlyTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r1_p1 RxDigStrbDlyTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r1_p1 TxDqDlyTg0_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r1_p1 TxDqDlyTg1_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r1_p1 DqRxVrefDac_r1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaRangeVal_p1 RxReplicaRangeVal_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl04_p1 RxReplicaCtl04_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r2_p1 RxClkT2UIDlyTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r2_p1 RxClkT2UIDlyTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r2_p1 RxClkC2UIDlyTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r2_p1 RxClkC2UIDlyTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r2_p1 TxDqLeftEyeOffsetTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r2_p1 TxDqLeftEyeOffsetTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r2_p1 TxDqRightEyeOffsetTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r2_p1 TxDqRightEyeOffsetTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r2_p1 RxClkTLeftEyeOffsetTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r2_p1 RxClkTLeftEyeOffsetTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r2_p1 RxClkTRightEyeOffsetTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r2_p1 RxClkTRightEyeOffsetTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r2_p1 RxClkCLeftEyeOffsetTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r2_p1 RxClkCLeftEyeOffsetTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r2_p1 RxClkCRightEyeOffsetTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r2_p1 RxClkCRightEyeOffsetTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r2_p1 RxDigStrbDlyTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r2_p1 RxDigStrbDlyTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r2_p1 TxDqDlyTg0_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r2_p1 TxDqDlyTg1_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase0_p1 RxReplicaPathPhase0_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase1_p1 RxReplicaPathPhase1_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase2_p1 RxReplicaPathPhase2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase3_p1 RxReplicaPathPhase3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase4_p1 RxReplicaPathPhase4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl01_p1 RxReplicaCtl01_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl02_p1 RxReplicaCtl02_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl03_p1 RxReplicaCtl03_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r2_p1 DqRxVrefDac_r2_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r3_p1 RxClkT2UIDlyTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r3_p1 RxClkT2UIDlyTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r3_p1 RxClkC2UIDlyTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r3_p1 RxClkC2UIDlyTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r3_p1 TxDqLeftEyeOffsetTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r3_p1 TxDqLeftEyeOffsetTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r3_p1 TxDqRightEyeOffsetTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r3_p1 TxDqRightEyeOffsetTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r3_p1 RxClkTLeftEyeOffsetTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r3_p1 RxClkTLeftEyeOffsetTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r3_p1 RxClkTRightEyeOffsetTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r3_p1 RxClkTRightEyeOffsetTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r3_p1 RxClkCLeftEyeOffsetTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r3_p1 RxClkCLeftEyeOffsetTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r3_p1 RxClkCRightEyeOffsetTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r3_p1 RxClkCRightEyeOffsetTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r3_p1 RxDigStrbDlyTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r3_p1 RxDigStrbDlyTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r3_p1 TxDqDlyTg0_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r3_p1 TxDqDlyTg1_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r3_p1 DqRxVrefDac_r3_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r4_p1 RxClkT2UIDlyTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r4_p1 RxClkT2UIDlyTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r4_p1 RxClkC2UIDlyTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r4_p1 RxClkC2UIDlyTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r4_p1 TxDqLeftEyeOffsetTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r4_p1 TxDqLeftEyeOffsetTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r4_p1 TxDqRightEyeOffsetTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r4_p1 TxDqRightEyeOffsetTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r4_p1 RxClkTLeftEyeOffsetTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r4_p1 RxClkTLeftEyeOffsetTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r4_p1 RxClkTRightEyeOffsetTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r4_p1 RxClkTRightEyeOffsetTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r4_p1 RxClkCLeftEyeOffsetTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r4_p1 RxClkCLeftEyeOffsetTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r4_p1 RxClkCRightEyeOffsetTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r4_p1 RxClkCRightEyeOffsetTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r4_p1 RxDigStrbDlyTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r4_p1 RxDigStrbDlyTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r4_p1 TxDqDlyTg0_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r4_p1 TxDqDlyTg1_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r4_p1 DqRxVrefDac_r4_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r5_p1 RxClkT2UIDlyTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r5_p1 RxClkT2UIDlyTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r5_p1 RxClkC2UIDlyTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r5_p1 RxClkC2UIDlyTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r5_p1 TxDqLeftEyeOffsetTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r5_p1 TxDqLeftEyeOffsetTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r5_p1 TxDqRightEyeOffsetTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r5_p1 TxDqRightEyeOffsetTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r5_p1 RxClkTLeftEyeOffsetTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r5_p1 RxClkTLeftEyeOffsetTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r5_p1 RxClkTRightEyeOffsetTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r5_p1 RxClkTRightEyeOffsetTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r5_p1 RxClkCLeftEyeOffsetTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r5_p1 RxClkCLeftEyeOffsetTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r5_p1 RxClkCRightEyeOffsetTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r5_p1 RxClkCRightEyeOffsetTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r5_p1 RxDigStrbDlyTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r5_p1 RxDigStrbDlyTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r5_p1 TxDqDlyTg0_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r5_p1 TxDqDlyTg1_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r5_p1 DqRxVrefDac_r5_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r6_p1 RxClkT2UIDlyTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r6_p1 RxClkT2UIDlyTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r6_p1 RxClkC2UIDlyTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r6_p1 RxClkC2UIDlyTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r6_p1 TxDqLeftEyeOffsetTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r6_p1 TxDqLeftEyeOffsetTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r6_p1 TxDqRightEyeOffsetTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r6_p1 TxDqRightEyeOffsetTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r6_p1 RxClkTLeftEyeOffsetTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r6_p1 RxClkTLeftEyeOffsetTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r6_p1 RxClkTRightEyeOffsetTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r6_p1 RxClkTRightEyeOffsetTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r6_p1 RxClkCLeftEyeOffsetTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r6_p1 RxClkCLeftEyeOffsetTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r6_p1 RxClkCRightEyeOffsetTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r6_p1 RxClkCRightEyeOffsetTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r6_p1 RxDigStrbDlyTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r6_p1 RxDigStrbDlyTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r6_p1 TxDqDlyTg0_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r6_p1 TxDqDlyTg1_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r6_p1 DqRxVrefDac_r6_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r7_p1 RxClkT2UIDlyTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r7_p1 RxClkT2UIDlyTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r7_p1 RxClkC2UIDlyTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r7_p1 RxClkC2UIDlyTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r7_p1 TxDqLeftEyeOffsetTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r7_p1 TxDqLeftEyeOffsetTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r7_p1 TxDqRightEyeOffsetTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r7_p1 TxDqRightEyeOffsetTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r7_p1 RxClkTLeftEyeOffsetTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r7_p1 RxClkTLeftEyeOffsetTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r7_p1 RxClkTRightEyeOffsetTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r7_p1 RxClkTRightEyeOffsetTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r7_p1 RxClkCLeftEyeOffsetTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r7_p1 RxClkCLeftEyeOffsetTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r7_p1 RxClkCRightEyeOffsetTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r7_p1 RxClkCRightEyeOffsetTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r7_p1 RxDigStrbDlyTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r7_p1 RxDigStrbDlyTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r7_p1 TxDqDlyTg0_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r7_p1 TxDqDlyTg1_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r7_p1 DqRxVrefDac_r7_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl0DB_p1 PclkDCAStaticCtrl0DB_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCASampDelayLCDLDB_p1 PclkDCASampDelayLCDLDB_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r8_p1 RxClkT2UIDlyTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r8_p1 RxClkT2UIDlyTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r8_p1 RxClkC2UIDlyTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r8_p1 RxClkC2UIDlyTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r8_p1 TxDqLeftEyeOffsetTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r8_p1 TxDqLeftEyeOffsetTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r8_p1 TxDqRightEyeOffsetTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r8_p1 TxDqRightEyeOffsetTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r8_p1 RxClkTLeftEyeOffsetTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r8_p1 RxClkTLeftEyeOffsetTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r8_p1 RxClkTRightEyeOffsetTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r8_p1 RxClkTRightEyeOffsetTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r8_p1 RxClkCLeftEyeOffsetTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r8_p1 RxClkCLeftEyeOffsetTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r8_p1 RxClkCRightEyeOffsetTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r8_p1 RxClkCRightEyeOffsetTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r8_p1 RxDigStrbDlyTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r8_p1 RxDigStrbDlyTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r8_p1 TxDqDlyTg0_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r8_p1 TxDqDlyTg1_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r8_p1 DqRxVrefDac_r8_p1;
	rand ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl1DB_p1 PclkDCAStaticCtrl1DB_p1;
   local uvm_reg_data_t m_offset;
	rand uvm_reg_field DFIMRL_p1_DFIMRL_p1;
	rand uvm_reg_field EnableWriteLinkEcc_p1_EnableWriteLinkEcc_p1;
	rand uvm_reg_field DxDfiClkDis_p1_DfiClkDqDis;
	rand uvm_reg_field DfiClkDqDis;
	rand uvm_reg_field DxDfiClkDis_p1_DfiClkDqsDis;
	rand uvm_reg_field DfiClkDqsDis;
	rand uvm_reg_field DxDfiClkDis_p1_DfiClkWckDis;
	rand uvm_reg_field DfiClkWckDis;
	rand uvm_reg_field DxPClkDis_p1_PClkDqDis;
	rand uvm_reg_field PClkDqDis;
	rand uvm_reg_field DxPClkDis_p1_PClkDqsDis;
	rand uvm_reg_field PClkDqsDis;
	rand uvm_reg_field DxPClkDis_p1_PClkWckDis;
	rand uvm_reg_field PClkWckDis;
	rand uvm_reg_field LP5DfiDataEnLatency_p1_LP5RLm13;
	rand uvm_reg_field LP5RLm13;
	rand uvm_reg_field PptDqsCntInvTrnTg0_p1_PptDqsCntInvTrnTg0_p1;
	rand uvm_reg_field PptDqsCntInvTrnTg1_p1_PptDqsCntInvTrnTg1_p1;
	rand uvm_reg_field TrackingModeCntrl_p1_EnWck2DqoSnoopTracking;
	rand uvm_reg_field EnWck2DqoSnoopTracking;
	rand uvm_reg_field TrackingModeCntrl_p1_Twck2dqoTrackingLimit;
	rand uvm_reg_field Twck2dqoTrackingLimit;
	rand uvm_reg_field TrackingModeCntrl_p1_ReservedTrackingModeCntrl;
	rand uvm_reg_field ReservedTrackingModeCntrl;
	rand uvm_reg_field TrackingModeCntrl_p1_Tdqs2dqTrackingLimit;
	rand uvm_reg_field Tdqs2dqTrackingLimit;
	rand uvm_reg_field TrackingModeCntrl_p1_DqsOscRunTimeSel;
	rand uvm_reg_field DqsOscRunTimeSel;
	rand uvm_reg_field TrackingModeCntrl_p1_RxDqsTrackingThreshold;
	rand uvm_reg_field RxDqsTrackingThreshold;
	rand uvm_reg_field RxClkT2UIDlyTg0_r0_p1_RxClkT2UIDlyTg0_r0_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r0_p1_RxClkT2UIDlyTg1_r0_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r0_p1_RxClkC2UIDlyTg0_r0_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r0_p1_RxClkC2UIDlyTg1_r0_p1;
	rand uvm_reg_field PptWck2DqoCntInvTrnTg0_p1_PptWck2DqoCntInvTrnTg0_p1;
	rand uvm_reg_field PptWck2DqoCntInvTrnTg1_p1_PptWck2DqoCntInvTrnTg1_p1;
	rand uvm_reg_field TxDqsLeftEyeOffsetTg0_p1_TxDqsLeftEyeOffsetTg0_p1;
	rand uvm_reg_field TxDqsLeftEyeOffsetTg1_p1_TxDqsLeftEyeOffsetTg1_p1;
	rand uvm_reg_field RxEnDlyTg0_p1_RxEnDlyTg0_p1;
	rand uvm_reg_field RxEnDlyTg1_p1_RxEnDlyTg1_p1;
	rand uvm_reg_field TxDqsRightEyeOffsetTg0_p1_TxDqsRightEyeOffsetTg0_p1;
	rand uvm_reg_field TxDqsRightEyeOffsetTg1_p1_TxDqsRightEyeOffsetTg1_p1;
	uvm_reg_field DqsPreambleControl_p1_Reserved;
	uvm_reg_field Reserved;
	rand uvm_reg_field DqsPreambleControl_p1_LP4PostambleExt;
	rand uvm_reg_field LP4PostambleExt;
	rand uvm_reg_field DqsPreambleControl_p1_WDQSEXTENSION;
	rand uvm_reg_field WDQSEXTENSION;
	rand uvm_reg_field DqsPreambleControl_p1_WCKEXTENSION;
	rand uvm_reg_field WCKEXTENSION;
	rand uvm_reg_field DqsPreambleControl_p1_DqPreOeExt;
	rand uvm_reg_field DqPreOeExt;
	rand uvm_reg_field DqsPreambleControl_p1_DqPstOeExt;
	rand uvm_reg_field DqPstOeExt;
	rand uvm_reg_field DbyteRxDqsModeCntrl_p1_RxPostambleMode;
	rand uvm_reg_field RxPostambleMode;
	rand uvm_reg_field DbyteRxDqsModeCntrl_p1_RxPreambleMode;
	rand uvm_reg_field RxPreambleMode;
	rand uvm_reg_field DbyteRxDqsModeCntrl_p1_LPDDR5RdqsEn;
	rand uvm_reg_field LPDDR5RdqsEn;
	rand uvm_reg_field DbyteRxDqsModeCntrl_p1_LPDDR5RdqsPre;
	rand uvm_reg_field LPDDR5RdqsPre;
	rand uvm_reg_field DbyteRxDqsModeCntrl_p1_LPDDR5RdqsPst;
	rand uvm_reg_field LPDDR5RdqsPst;
	rand uvm_reg_field DbyteRxDqsModeCntrl_p1_PositionDfeInit;
	rand uvm_reg_field PositionDfeInit;
	rand uvm_reg_field DbyteRxDqsModeCntrl_p1_PositionRxPhaseUpdate;
	rand uvm_reg_field PositionRxPhaseUpdate;
	rand uvm_reg_field RxClkCntl1_p1_EnRxClkCor;
	rand uvm_reg_field EnRxClkCor;
	rand uvm_reg_field TxDqsDlyTg0_p1_TxDqsDlyTg0_p1;
	rand uvm_reg_field TxDqsDlyTg1_p1_TxDqsDlyTg1_p1;
	rand uvm_reg_field TxWckDlyTg0_p1_TxWckDlyTg0_p1;
	rand uvm_reg_field TxWckDlyTg1_p1_TxWckDlyTg1_p1;
	rand uvm_reg_field RxModeCtlRxReplica_p1_RxModeCtlRxReplica_p1;
	rand uvm_reg_field RxGainCurrAdjRxReplica_p1_RxGainCurrAdjRxReplica_p1;
	rand uvm_reg_field DxRxStandbyEn_p1_DxRxStandbyEn_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r0_p1_TxDqLeftEyeOffsetTg0_r0_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r0_p1_TxDqLeftEyeOffsetTg1_r0_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r0_p1_TxDqRightEyeOffsetTg0_r0_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r0_p1_TxDqRightEyeOffsetTg1_r0_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r0_p1_RxClkTLeftEyeOffsetTg0_r0_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r0_p1_RxClkTLeftEyeOffsetTg1_r0_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r0_p1_RxClkTRightEyeOffsetTg0_r0_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r0_p1_RxClkTRightEyeOffsetTg1_r0_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r0_p1_RxClkCLeftEyeOffsetTg0_r0_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r0_p1_RxClkCLeftEyeOffsetTg1_r0_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r0_p1_RxClkCRightEyeOffsetTg0_r0_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r0_p1_RxClkCRightEyeOffsetTg1_r0_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r0_p1_RxDigStrbDlyTg0_r0_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r0_p1_RxDigStrbDlyTg1_r0_p1;
	rand uvm_reg_field TxDqDlyTg0_r0_p1_TxDqDlyTg0_r0_p1;
	rand uvm_reg_field TxDqDlyTg1_r0_p1_TxDqDlyTg1_r0_p1;
	rand uvm_reg_field SingleEndedMode_p1_SingleEndedModeReserved;
	rand uvm_reg_field SingleEndedModeReserved;
	rand uvm_reg_field SingleEndedMode_p1_SingleEndedDQS;
	rand uvm_reg_field SingleEndedDQS;
	rand uvm_reg_field SingleEndedMode_p1_SingleEndedWCK;
	rand uvm_reg_field SingleEndedWCK;
	rand uvm_reg_field RxTrainPattern8BitMode_p1_RxTrainPattern8BitMode_p1;
	rand uvm_reg_field DqRxVrefDac_r0_p1_DqRxVrefDac_r0_p1;
	rand uvm_reg_field RxDigStrbEn_p1_EnStrblssRdMode;
	rand uvm_reg_field EnStrblssRdMode;
	rand uvm_reg_field RxDigStrbEn_p1_RxReplicaPowerDownNoRDQS;
	rand uvm_reg_field RxReplicaPowerDownNoRDQS;
	rand uvm_reg_field RxDigStrbEn_p1_OdtDisDqs;
	rand uvm_reg_field OdtDisDqs;
	rand uvm_reg_field DxPipeEn_p1_DxWrPipeEn;
	rand uvm_reg_field DxWrPipeEn;
	rand uvm_reg_field DxPipeEn_p1_DxRdPipeEn;
	rand uvm_reg_field DxRdPipeEn;
	rand uvm_reg_field PclkDCDCtrl_p1_PclkDCDEn;
	rand uvm_reg_field PclkDCDEn;
	rand uvm_reg_field PclkDCDCtrl_p1_PclkDCDOffsetMode;
	rand uvm_reg_field PclkDCDOffsetMode;
	rand uvm_reg_field PPTTrainSetup2_p1_PPTTrainSetup2_p1;
	rand uvm_reg_field DMIPinPresent_p1_RdDbiEnabled;
	rand uvm_reg_field RdDbiEnabled;
	rand uvm_reg_field InhibitTxRdPtrInit_p1_InhibitTxRdPtrInit_p1;
	rand uvm_reg_field RxClkT2UIDlyTg0_r1_p1_RxClkT2UIDlyTg0_r1_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r1_p1_RxClkT2UIDlyTg1_r1_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r1_p1_RxClkC2UIDlyTg0_r1_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r1_p1_RxClkC2UIDlyTg1_r1_p1;
	rand uvm_reg_field RDqRDqsCntrl_p1_RxPubLcdlSeed;
	rand uvm_reg_field RxPubLcdlSeed;
	rand uvm_reg_field RDqRDqsCntrl_p1_RDqRDqsCntrl9;
	rand uvm_reg_field RDqRDqsCntrl9;
	rand uvm_reg_field RDqRDqsCntrl_p1_RxPubCalModeIs1UI;
	rand uvm_reg_field RxPubCalModeIs1UI;
	rand uvm_reg_field RDqRDqsCntrl_p1_RxPubCntlByPState;
	rand uvm_reg_field RxPubCntlByPState;
	rand uvm_reg_field RDqRDqsCntrl_p1_RxPubRxReplicaCalModeIs1UI;
	rand uvm_reg_field RxPubRxReplicaCalModeIs1UI;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r1_p1_TxDqLeftEyeOffsetTg0_r1_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r1_p1_TxDqLeftEyeOffsetTg1_r1_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r1_p1_TxDqRightEyeOffsetTg0_r1_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r1_p1_TxDqRightEyeOffsetTg1_r1_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r1_p1_RxClkTLeftEyeOffsetTg0_r1_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r1_p1_RxClkTLeftEyeOffsetTg1_r1_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r1_p1_RxClkTRightEyeOffsetTg0_r1_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r1_p1_RxClkTRightEyeOffsetTg1_r1_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r1_p1_RxClkCLeftEyeOffsetTg0_r1_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r1_p1_RxClkCLeftEyeOffsetTg1_r1_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r1_p1_RxClkCRightEyeOffsetTg0_r1_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r1_p1_RxClkCRightEyeOffsetTg1_r1_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r1_p1_RxDigStrbDlyTg0_r1_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r1_p1_RxDigStrbDlyTg1_r1_p1;
	rand uvm_reg_field TxDqDlyTg0_r1_p1_TxDqDlyTg0_r1_p1;
	rand uvm_reg_field TxDqDlyTg1_r1_p1_TxDqDlyTg1_r1_p1;
	rand uvm_reg_field DqRxVrefDac_r1_p1_DqRxVrefDac_r1_p1;
	rand uvm_reg_field RxReplicaRangeVal_p1_RxReplicaShortCalRangeA;
	rand uvm_reg_field RxReplicaShortCalRangeA;
	rand uvm_reg_field RxReplicaRangeVal_p1_RxReplicaShortCalRangeB;
	rand uvm_reg_field RxReplicaShortCalRangeB;
	rand uvm_reg_field RxReplicaCtl04_p1_RxReplicaTrackEn;
	rand uvm_reg_field RxReplicaTrackEn;
	rand uvm_reg_field RxReplicaCtl04_p1_RxReplicaLongCal;
	rand uvm_reg_field RxReplicaLongCal;
	rand uvm_reg_field RxReplicaCtl04_p1_RxReplicaStride;
	rand uvm_reg_field RxReplicaStride;
	rand uvm_reg_field RxReplicaCtl04_p1_RxReplicaStandby;
	rand uvm_reg_field RxReplicaStandby;
	rand uvm_reg_field RxReplicaCtl04_p1_RxReplicaPDenFSM;
	rand uvm_reg_field RxReplicaPDenFSM;
	rand uvm_reg_field RxReplicaCtl04_p1_RxReplicaPDRecoverytime;
	rand uvm_reg_field RxReplicaPDRecoverytime;
	rand uvm_reg_field RxClkT2UIDlyTg0_r2_p1_RxClkT2UIDlyTg0_r2_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r2_p1_RxClkT2UIDlyTg1_r2_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r2_p1_RxClkC2UIDlyTg0_r2_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r2_p1_RxClkC2UIDlyTg1_r2_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r2_p1_TxDqLeftEyeOffsetTg0_r2_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r2_p1_TxDqLeftEyeOffsetTg1_r2_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r2_p1_TxDqRightEyeOffsetTg0_r2_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r2_p1_TxDqRightEyeOffsetTg1_r2_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r2_p1_RxClkTLeftEyeOffsetTg0_r2_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r2_p1_RxClkTLeftEyeOffsetTg1_r2_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r2_p1_RxClkTRightEyeOffsetTg0_r2_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r2_p1_RxClkTRightEyeOffsetTg1_r2_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r2_p1_RxClkCLeftEyeOffsetTg0_r2_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r2_p1_RxClkCLeftEyeOffsetTg1_r2_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r2_p1_RxClkCRightEyeOffsetTg0_r2_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r2_p1_RxClkCRightEyeOffsetTg1_r2_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r2_p1_RxDigStrbDlyTg0_r2_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r2_p1_RxDigStrbDlyTg1_r2_p1;
	rand uvm_reg_field TxDqDlyTg0_r2_p1_TxDqDlyTg0_r2_p1;
	rand uvm_reg_field TxDqDlyTg1_r2_p1_TxDqDlyTg1_r2_p1;
	rand uvm_reg_field RxReplicaPathPhase0_p1_RxReplicaPathPhase0_p1;
	rand uvm_reg_field RxReplicaPathPhase1_p1_RxReplicaPathPhase1_p1;
	rand uvm_reg_field RxReplicaPathPhase2_p1_RxReplicaPathPhase2_p1;
	rand uvm_reg_field RxReplicaPathPhase3_p1_RxReplicaPathPhase3_p1;
	rand uvm_reg_field RxReplicaPathPhase4_p1_RxReplicaPathPhase4_p1;
	rand uvm_reg_field RxReplicaCtl01_p1_RxReplicaSelPathPhase;
	rand uvm_reg_field RxReplicaSelPathPhase;
	rand uvm_reg_field RxReplicaCtl02_p1_RxReplicaDiffLimit;
	rand uvm_reg_field RxReplicaDiffLimit;
	rand uvm_reg_field RxReplicaCtl03_p1_RxReplicaRatioTrn;
	rand uvm_reg_field RxReplicaRatioTrn;
	rand uvm_reg_field DqRxVrefDac_r2_p1_DqRxVrefDac_r2_p1;
	rand uvm_reg_field RxClkT2UIDlyTg0_r3_p1_RxClkT2UIDlyTg0_r3_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r3_p1_RxClkT2UIDlyTg1_r3_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r3_p1_RxClkC2UIDlyTg0_r3_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r3_p1_RxClkC2UIDlyTg1_r3_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r3_p1_TxDqLeftEyeOffsetTg0_r3_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r3_p1_TxDqLeftEyeOffsetTg1_r3_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r3_p1_TxDqRightEyeOffsetTg0_r3_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r3_p1_TxDqRightEyeOffsetTg1_r3_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r3_p1_RxClkTLeftEyeOffsetTg0_r3_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r3_p1_RxClkTLeftEyeOffsetTg1_r3_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r3_p1_RxClkTRightEyeOffsetTg0_r3_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r3_p1_RxClkTRightEyeOffsetTg1_r3_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r3_p1_RxClkCLeftEyeOffsetTg0_r3_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r3_p1_RxClkCLeftEyeOffsetTg1_r3_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r3_p1_RxClkCRightEyeOffsetTg0_r3_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r3_p1_RxClkCRightEyeOffsetTg1_r3_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r3_p1_RxDigStrbDlyTg0_r3_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r3_p1_RxDigStrbDlyTg1_r3_p1;
	rand uvm_reg_field TxDqDlyTg0_r3_p1_TxDqDlyTg0_r3_p1;
	rand uvm_reg_field TxDqDlyTg1_r3_p1_TxDqDlyTg1_r3_p1;
	rand uvm_reg_field DqRxVrefDac_r3_p1_DqRxVrefDac_r3_p1;
	rand uvm_reg_field RxClkT2UIDlyTg0_r4_p1_RxClkT2UIDlyTg0_r4_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r4_p1_RxClkT2UIDlyTg1_r4_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r4_p1_RxClkC2UIDlyTg0_r4_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r4_p1_RxClkC2UIDlyTg1_r4_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r4_p1_TxDqLeftEyeOffsetTg0_r4_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r4_p1_TxDqLeftEyeOffsetTg1_r4_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r4_p1_TxDqRightEyeOffsetTg0_r4_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r4_p1_TxDqRightEyeOffsetTg1_r4_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r4_p1_RxClkTLeftEyeOffsetTg0_r4_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r4_p1_RxClkTLeftEyeOffsetTg1_r4_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r4_p1_RxClkTRightEyeOffsetTg0_r4_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r4_p1_RxClkTRightEyeOffsetTg1_r4_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r4_p1_RxClkCLeftEyeOffsetTg0_r4_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r4_p1_RxClkCLeftEyeOffsetTg1_r4_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r4_p1_RxClkCRightEyeOffsetTg0_r4_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r4_p1_RxClkCRightEyeOffsetTg1_r4_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r4_p1_RxDigStrbDlyTg0_r4_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r4_p1_RxDigStrbDlyTg1_r4_p1;
	rand uvm_reg_field TxDqDlyTg0_r4_p1_TxDqDlyTg0_r4_p1;
	rand uvm_reg_field TxDqDlyTg1_r4_p1_TxDqDlyTg1_r4_p1;
	rand uvm_reg_field DqRxVrefDac_r4_p1_DqRxVrefDac_r4_p1;
	rand uvm_reg_field RxClkT2UIDlyTg0_r5_p1_RxClkT2UIDlyTg0_r5_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r5_p1_RxClkT2UIDlyTg1_r5_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r5_p1_RxClkC2UIDlyTg0_r5_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r5_p1_RxClkC2UIDlyTg1_r5_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r5_p1_TxDqLeftEyeOffsetTg0_r5_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r5_p1_TxDqLeftEyeOffsetTg1_r5_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r5_p1_TxDqRightEyeOffsetTg0_r5_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r5_p1_TxDqRightEyeOffsetTg1_r5_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r5_p1_RxClkTLeftEyeOffsetTg0_r5_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r5_p1_RxClkTLeftEyeOffsetTg1_r5_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r5_p1_RxClkTRightEyeOffsetTg0_r5_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r5_p1_RxClkTRightEyeOffsetTg1_r5_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r5_p1_RxClkCLeftEyeOffsetTg0_r5_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r5_p1_RxClkCLeftEyeOffsetTg1_r5_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r5_p1_RxClkCRightEyeOffsetTg0_r5_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r5_p1_RxClkCRightEyeOffsetTg1_r5_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r5_p1_RxDigStrbDlyTg0_r5_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r5_p1_RxDigStrbDlyTg1_r5_p1;
	rand uvm_reg_field TxDqDlyTg0_r5_p1_TxDqDlyTg0_r5_p1;
	rand uvm_reg_field TxDqDlyTg1_r5_p1_TxDqDlyTg1_r5_p1;
	rand uvm_reg_field DqRxVrefDac_r5_p1_DqRxVrefDac_r5_p1;
	rand uvm_reg_field RxClkT2UIDlyTg0_r6_p1_RxClkT2UIDlyTg0_r6_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r6_p1_RxClkT2UIDlyTg1_r6_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r6_p1_RxClkC2UIDlyTg0_r6_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r6_p1_RxClkC2UIDlyTg1_r6_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r6_p1_TxDqLeftEyeOffsetTg0_r6_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r6_p1_TxDqLeftEyeOffsetTg1_r6_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r6_p1_TxDqRightEyeOffsetTg0_r6_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r6_p1_TxDqRightEyeOffsetTg1_r6_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r6_p1_RxClkTLeftEyeOffsetTg0_r6_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r6_p1_RxClkTLeftEyeOffsetTg1_r6_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r6_p1_RxClkTRightEyeOffsetTg0_r6_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r6_p1_RxClkTRightEyeOffsetTg1_r6_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r6_p1_RxClkCLeftEyeOffsetTg0_r6_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r6_p1_RxClkCLeftEyeOffsetTg1_r6_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r6_p1_RxClkCRightEyeOffsetTg0_r6_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r6_p1_RxClkCRightEyeOffsetTg1_r6_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r6_p1_RxDigStrbDlyTg0_r6_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r6_p1_RxDigStrbDlyTg1_r6_p1;
	rand uvm_reg_field TxDqDlyTg0_r6_p1_TxDqDlyTg0_r6_p1;
	rand uvm_reg_field TxDqDlyTg1_r6_p1_TxDqDlyTg1_r6_p1;
	rand uvm_reg_field DqRxVrefDac_r6_p1_DqRxVrefDac_r6_p1;
	rand uvm_reg_field RxClkT2UIDlyTg0_r7_p1_RxClkT2UIDlyTg0_r7_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r7_p1_RxClkT2UIDlyTg1_r7_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r7_p1_RxClkC2UIDlyTg0_r7_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r7_p1_RxClkC2UIDlyTg1_r7_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r7_p1_TxDqLeftEyeOffsetTg0_r7_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r7_p1_TxDqLeftEyeOffsetTg1_r7_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r7_p1_TxDqRightEyeOffsetTg0_r7_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r7_p1_TxDqRightEyeOffsetTg1_r7_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r7_p1_RxClkTLeftEyeOffsetTg0_r7_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r7_p1_RxClkTLeftEyeOffsetTg1_r7_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r7_p1_RxClkTRightEyeOffsetTg0_r7_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r7_p1_RxClkTRightEyeOffsetTg1_r7_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r7_p1_RxClkCLeftEyeOffsetTg0_r7_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r7_p1_RxClkCLeftEyeOffsetTg1_r7_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r7_p1_RxClkCRightEyeOffsetTg0_r7_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r7_p1_RxClkCRightEyeOffsetTg1_r7_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r7_p1_RxDigStrbDlyTg0_r7_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r7_p1_RxDigStrbDlyTg1_r7_p1;
	rand uvm_reg_field TxDqDlyTg0_r7_p1_TxDqDlyTg0_r7_p1;
	rand uvm_reg_field TxDqDlyTg1_r7_p1_TxDqDlyTg1_r7_p1;
	rand uvm_reg_field DqRxVrefDac_r7_p1_DqRxVrefDac_r7_p1;
	rand uvm_reg_field PclkDCAStaticCtrl0DB_p1_PclkDCACalModeDB;
	rand uvm_reg_field PclkDCACalModeDB;
	rand uvm_reg_field PclkDCAStaticCtrl0DB_p1_PclkDCAEnDB;
	rand uvm_reg_field PclkDCAEnDB;
	rand uvm_reg_field PclkDCAStaticCtrl0DB_p1_PclkDCATxLcdlPhSelDB;
	rand uvm_reg_field PclkDCATxLcdlPhSelDB;
	rand uvm_reg_field PclkDCAStaticCtrl0DB_p1_PclkDCDSettleDB;
	rand uvm_reg_field PclkDCDSettleDB;
	rand uvm_reg_field PclkDCAStaticCtrl0DB_p1_PclkDCDSampTimeDB;
	rand uvm_reg_field PclkDCDSampTimeDB;
	rand uvm_reg_field PclkDCASampDelayLCDLDB_p1_PclkDCASampDelayLCDLDB_p1;
	rand uvm_reg_field RxClkT2UIDlyTg0_r8_p1_RxClkT2UIDlyTg0_r8_p1;
	rand uvm_reg_field RxClkT2UIDlyTg1_r8_p1_RxClkT2UIDlyTg1_r8_p1;
	rand uvm_reg_field RxClkC2UIDlyTg0_r8_p1_RxClkC2UIDlyTg0_r8_p1;
	rand uvm_reg_field RxClkC2UIDlyTg1_r8_p1_RxClkC2UIDlyTg1_r8_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg0_r8_p1_TxDqLeftEyeOffsetTg0_r8_p1;
	rand uvm_reg_field TxDqLeftEyeOffsetTg1_r8_p1_TxDqLeftEyeOffsetTg1_r8_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg0_r8_p1_TxDqRightEyeOffsetTg0_r8_p1;
	rand uvm_reg_field TxDqRightEyeOffsetTg1_r8_p1_TxDqRightEyeOffsetTg1_r8_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg0_r8_p1_RxClkTLeftEyeOffsetTg0_r8_p1;
	rand uvm_reg_field RxClkTLeftEyeOffsetTg1_r8_p1_RxClkTLeftEyeOffsetTg1_r8_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg0_r8_p1_RxClkTRightEyeOffsetTg0_r8_p1;
	rand uvm_reg_field RxClkTRightEyeOffsetTg1_r8_p1_RxClkTRightEyeOffsetTg1_r8_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg0_r8_p1_RxClkCLeftEyeOffsetTg0_r8_p1;
	rand uvm_reg_field RxClkCLeftEyeOffsetTg1_r8_p1_RxClkCLeftEyeOffsetTg1_r8_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg0_r8_p1_RxClkCRightEyeOffsetTg0_r8_p1;
	rand uvm_reg_field RxClkCRightEyeOffsetTg1_r8_p1_RxClkCRightEyeOffsetTg1_r8_p1;
	rand uvm_reg_field RxDigStrbDlyTg0_r8_p1_RxDigStrbDlyTg0_r8_p1;
	rand uvm_reg_field RxDigStrbDlyTg1_r8_p1_RxDigStrbDlyTg1_r8_p1;
	rand uvm_reg_field TxDqDlyTg0_r8_p1_TxDqDlyTg0_r8_p1;
	rand uvm_reg_field TxDqDlyTg1_r8_p1_TxDqDlyTg1_r8_p1;
	rand uvm_reg_field DqRxVrefDac_r8_p1_DqRxVrefDac_r8_p1;
	rand uvm_reg_field PclkDCAStaticCtrl1DB_p1_PclkDCAInvertSampDB;
	rand uvm_reg_field PclkDCAInvertSampDB;
	rand uvm_reg_field PclkDCAStaticCtrl1DB_p1_PclkDCALcdlEn4pDB;
	rand uvm_reg_field PclkDCALcdlEn4pDB;
	rand uvm_reg_field PclkDCAStaticCtrl1DB_p1_PclkDCDMissionModeDelayDB;
	rand uvm_reg_field PclkDCDMissionModeDelayDB;


	covergroup cg_addr (input string name);
	option.per_instance = 1;
option.name = get_name();

	DFIMRL_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h0 };
		option.weight = 1;
	}

	EnableWriteLinkEcc_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1 };
		option.weight = 1;
	}

	DxDfiClkDis_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3 };
		option.weight = 1;
	}

	DxPClkDis_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h4 };
		option.weight = 1;
	}

	LP5DfiDataEnLatency_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h8 };
		option.weight = 1;
	}

	PptDqsCntInvTrnTg0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hC };
		option.weight = 1;
	}

	PptDqsCntInvTrnTg1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hD };
		option.weight = 1;
	}

	TrackingModeCntrl_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hE };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h10 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h11 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h12 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h13 };
		option.weight = 1;
	}

	PptWck2DqoCntInvTrnTg0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h14 };
		option.weight = 1;
	}

	PptWck2DqoCntInvTrnTg1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h15 };
		option.weight = 1;
	}

	TxDqsLeftEyeOffsetTg0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h19 };
		option.weight = 1;
	}

	TxDqsLeftEyeOffsetTg1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1B };
		option.weight = 1;
	}

	RxEnDlyTg0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20 };
		option.weight = 1;
	}

	RxEnDlyTg1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h21 };
		option.weight = 1;
	}

	TxDqsRightEyeOffsetTg0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h22 };
		option.weight = 1;
	}

	TxDqsRightEyeOffsetTg1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h23 };
		option.weight = 1;
	}

	DqsPreambleControl_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h24 };
		option.weight = 1;
	}

	DbyteRxDqsModeCntrl_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h25 };
		option.weight = 1;
	}

	RxClkCntl1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h27 };
		option.weight = 1;
	}

	TxDqsDlyTg0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h28 };
		option.weight = 1;
	}

	TxDqsDlyTg1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h29 };
		option.weight = 1;
	}

	TxWckDlyTg0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2A };
		option.weight = 1;
	}

	TxWckDlyTg1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2B };
		option.weight = 1;
	}

	RxModeCtlRxReplica_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h39 };
		option.weight = 1;
	}

	RxGainCurrAdjRxReplica_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3E };
		option.weight = 1;
	}

	DxRxStandbyEn_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h5F };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h60 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h61 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h63 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h64 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h68 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h69 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h78 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h79 };
		option.weight = 1;
	}

	TxDqDlyTg0_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h7A };
		option.weight = 1;
	}

	TxDqDlyTg1_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h7B };
		option.weight = 1;
	}

	SingleEndedMode_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h7C };
		option.weight = 1;
	}

	RxTrainPattern8BitMode_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hA5 };
		option.weight = 1;
	}

	DqRxVrefDac_r0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hC8 };
		option.weight = 1;
	}

	RxDigStrbEn_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hFB };
		option.weight = 1;
	}

	DxPipeEn_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hFC };
		option.weight = 1;
	}

	PclkDCDCtrl_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h100 };
		option.weight = 1;
	}

	PPTTrainSetup2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h102 };
		option.weight = 1;
	}

	DMIPinPresent_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h108 };
		option.weight = 1;
	}

	InhibitTxRdPtrInit_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h10B };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h110 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h111 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h112 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h113 };
		option.weight = 1;
	}

	RDqRDqsCntrl_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h15F };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h160 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h161 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h163 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h164 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h168 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h169 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h16A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h16B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h16C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h16D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h16E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h16F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h178 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h179 };
		option.weight = 1;
	}

	TxDqDlyTg0_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h17A };
		option.weight = 1;
	}

	TxDqDlyTg1_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h17B };
		option.weight = 1;
	}

	DqRxVrefDac_r1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h1C8 };
		option.weight = 1;
	}

	RxReplicaRangeVal_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h209 };
		option.weight = 1;
	}

	RxReplicaCtl04_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h20F };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h210 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h211 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h212 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h213 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h260 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h261 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h263 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h264 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h268 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h269 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h26A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h26B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h26C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h26D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h26E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h26F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h278 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h279 };
		option.weight = 1;
	}

	TxDqDlyTg0_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h27A };
		option.weight = 1;
	}

	TxDqDlyTg1_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h27B };
		option.weight = 1;
	}

	RxReplicaPathPhase0_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2A0 };
		option.weight = 1;
	}

	RxReplicaPathPhase1_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2A1 };
		option.weight = 1;
	}

	RxReplicaPathPhase2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2A2 };
		option.weight = 1;
	}

	RxReplicaPathPhase3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2A3 };
		option.weight = 1;
	}

	RxReplicaPathPhase4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2A4 };
		option.weight = 1;
	}

	RxReplicaCtl01_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2AD };
		option.weight = 1;
	}

	RxReplicaCtl02_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2AE };
		option.weight = 1;
	}

	RxReplicaCtl03_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2AF };
		option.weight = 1;
	}

	DqRxVrefDac_r2_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h2C8 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h310 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h311 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h312 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h313 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h360 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h361 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h363 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h364 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h368 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h369 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h36A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h36B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h36C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h36D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h36E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h36F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h378 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h379 };
		option.weight = 1;
	}

	TxDqDlyTg0_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h37A };
		option.weight = 1;
	}

	TxDqDlyTg1_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h37B };
		option.weight = 1;
	}

	DqRxVrefDac_r3_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h3C8 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h410 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h411 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h412 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h413 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h460 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h461 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h463 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h464 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h468 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h469 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h46A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h46B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h46C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h46D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h46E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h46F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h478 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h479 };
		option.weight = 1;
	}

	TxDqDlyTg0_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h47A };
		option.weight = 1;
	}

	TxDqDlyTg1_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h47B };
		option.weight = 1;
	}

	DqRxVrefDac_r4_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h4C8 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h510 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h511 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h512 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h513 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h560 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h561 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h563 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h564 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h568 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h569 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h56A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h56B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h56C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h56D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h56E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h56F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h578 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h579 };
		option.weight = 1;
	}

	TxDqDlyTg0_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h57A };
		option.weight = 1;
	}

	TxDqDlyTg1_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h57B };
		option.weight = 1;
	}

	DqRxVrefDac_r5_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h5C8 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h610 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h611 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h612 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h613 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h660 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h661 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h663 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h664 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h668 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h669 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h66A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h66B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h66C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h66D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h66E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h66F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h678 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h679 };
		option.weight = 1;
	}

	TxDqDlyTg0_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h67A };
		option.weight = 1;
	}

	TxDqDlyTg1_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h67B };
		option.weight = 1;
	}

	DqRxVrefDac_r6_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h6C8 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h710 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h711 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h712 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h713 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h760 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h761 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h763 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h764 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h768 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h769 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h76A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h76B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h76C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h76D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h76E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h76F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h778 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h779 };
		option.weight = 1;
	}

	TxDqDlyTg0_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h77A };
		option.weight = 1;
	}

	TxDqDlyTg1_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h77B };
		option.weight = 1;
	}

	DqRxVrefDac_r7_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h7C8 };
		option.weight = 1;
	}

	PclkDCAStaticCtrl0DB_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h803 };
		option.weight = 1;
	}

	PclkDCASampDelayLCDLDB_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h80B };
		option.weight = 1;
	}

	RxClkT2UIDlyTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h810 };
		option.weight = 1;
	}

	RxClkT2UIDlyTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h811 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h812 };
		option.weight = 1;
	}

	RxClkC2UIDlyTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h813 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h860 };
		option.weight = 1;
	}

	TxDqLeftEyeOffsetTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h861 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h863 };
		option.weight = 1;
	}

	TxDqRightEyeOffsetTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h864 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h868 };
		option.weight = 1;
	}

	RxClkTLeftEyeOffsetTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h869 };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h86A };
		option.weight = 1;
	}

	RxClkTRightEyeOffsetTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h86B };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h86C };
		option.weight = 1;
	}

	RxClkCLeftEyeOffsetTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h86D };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h86E };
		option.weight = 1;
	}

	RxClkCRightEyeOffsetTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h86F };
		option.weight = 1;
	}

	RxDigStrbDlyTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h878 };
		option.weight = 1;
	}

	RxDigStrbDlyTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h879 };
		option.weight = 1;
	}

	TxDqDlyTg0_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h87A };
		option.weight = 1;
	}

	TxDqDlyTg1_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h87B };
		option.weight = 1;
	}

	DqRxVrefDac_r8_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h8C8 };
		option.weight = 1;
	}

	PclkDCAStaticCtrl1DB_p1 : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'hC03 };
		option.weight = 1;
	}
endgroup
	function new(string name = "DWC_DDRPHYA_DBYTE3_p1");
		super.new(name, build_coverage(UVM_CVR_ADDR_MAP));
		add_coverage(build_coverage(UVM_CVR_ADDR_MAP));
		if (has_coverage(UVM_CVR_ADDR_MAP))
			cg_addr = new("cg_addr");
	endfunction: new

   virtual function void build();
      this.default_map = create_map("", 0, 4, UVM_LITTLE_ENDIAN, 0);
      this.DFIMRL_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DFIMRL_p1::type_id::create("DFIMRL_p1",,get_full_name());
      if(this.DFIMRL_p1.has_coverage(UVM_CVR_ALL))
      	this.DFIMRL_p1.cg_bits.option.name = {get_name(), ".", "DFIMRL_p1_bits"};
      this.DFIMRL_p1.configure(this, null, "");
      this.DFIMRL_p1.build();
      this.default_map.add_reg(this.DFIMRL_p1, `UVM_REG_ADDR_WIDTH'h0, "RW", 0);
		this.DFIMRL_p1_DFIMRL_p1 = this.DFIMRL_p1.DFIMRL_p1;
      this.EnableWriteLinkEcc_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_EnableWriteLinkEcc_p1::type_id::create("EnableWriteLinkEcc_p1",,get_full_name());
      if(this.EnableWriteLinkEcc_p1.has_coverage(UVM_CVR_ALL))
      	this.EnableWriteLinkEcc_p1.cg_bits.option.name = {get_name(), ".", "EnableWriteLinkEcc_p1_bits"};
      this.EnableWriteLinkEcc_p1.configure(this, null, "");
      this.EnableWriteLinkEcc_p1.build();
      this.default_map.add_reg(this.EnableWriteLinkEcc_p1, `UVM_REG_ADDR_WIDTH'h1, "RW", 0);
		this.EnableWriteLinkEcc_p1_EnableWriteLinkEcc_p1 = this.EnableWriteLinkEcc_p1.EnableWriteLinkEcc_p1;
      this.DxDfiClkDis_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxDfiClkDis_p1::type_id::create("DxDfiClkDis_p1",,get_full_name());
      if(this.DxDfiClkDis_p1.has_coverage(UVM_CVR_ALL))
      	this.DxDfiClkDis_p1.cg_bits.option.name = {get_name(), ".", "DxDfiClkDis_p1_bits"};
      this.DxDfiClkDis_p1.configure(this, null, "");
      this.DxDfiClkDis_p1.build();
      this.default_map.add_reg(this.DxDfiClkDis_p1, `UVM_REG_ADDR_WIDTH'h3, "RW", 0);
		this.DxDfiClkDis_p1_DfiClkDqDis = this.DxDfiClkDis_p1.DfiClkDqDis;
		this.DfiClkDqDis = this.DxDfiClkDis_p1.DfiClkDqDis;
		this.DxDfiClkDis_p1_DfiClkDqsDis = this.DxDfiClkDis_p1.DfiClkDqsDis;
		this.DfiClkDqsDis = this.DxDfiClkDis_p1.DfiClkDqsDis;
		this.DxDfiClkDis_p1_DfiClkWckDis = this.DxDfiClkDis_p1.DfiClkWckDis;
		this.DfiClkWckDis = this.DxDfiClkDis_p1.DfiClkWckDis;
      this.DxPClkDis_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPClkDis_p1::type_id::create("DxPClkDis_p1",,get_full_name());
      if(this.DxPClkDis_p1.has_coverage(UVM_CVR_ALL))
      	this.DxPClkDis_p1.cg_bits.option.name = {get_name(), ".", "DxPClkDis_p1_bits"};
      this.DxPClkDis_p1.configure(this, null, "");
      this.DxPClkDis_p1.build();
      this.default_map.add_reg(this.DxPClkDis_p1, `UVM_REG_ADDR_WIDTH'h4, "RW", 0);
		this.DxPClkDis_p1_PClkDqDis = this.DxPClkDis_p1.PClkDqDis;
		this.PClkDqDis = this.DxPClkDis_p1.PClkDqDis;
		this.DxPClkDis_p1_PClkDqsDis = this.DxPClkDis_p1.PClkDqsDis;
		this.PClkDqsDis = this.DxPClkDis_p1.PClkDqsDis;
		this.DxPClkDis_p1_PClkWckDis = this.DxPClkDis_p1.PClkWckDis;
		this.PClkWckDis = this.DxPClkDis_p1.PClkWckDis;
      this.LP5DfiDataEnLatency_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_LP5DfiDataEnLatency_p1::type_id::create("LP5DfiDataEnLatency_p1",,get_full_name());
      if(this.LP5DfiDataEnLatency_p1.has_coverage(UVM_CVR_ALL))
      	this.LP5DfiDataEnLatency_p1.cg_bits.option.name = {get_name(), ".", "LP5DfiDataEnLatency_p1_bits"};
      this.LP5DfiDataEnLatency_p1.configure(this, null, "");
      this.LP5DfiDataEnLatency_p1.build();
      this.default_map.add_reg(this.LP5DfiDataEnLatency_p1, `UVM_REG_ADDR_WIDTH'h8, "RW", 0);
		this.LP5DfiDataEnLatency_p1_LP5RLm13 = this.LP5DfiDataEnLatency_p1.LP5RLm13;
		this.LP5RLm13 = this.LP5DfiDataEnLatency_p1.LP5RLm13;
      this.PptDqsCntInvTrnTg0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg0_p1::type_id::create("PptDqsCntInvTrnTg0_p1",,get_full_name());
      if(this.PptDqsCntInvTrnTg0_p1.has_coverage(UVM_CVR_ALL))
      	this.PptDqsCntInvTrnTg0_p1.cg_bits.option.name = {get_name(), ".", "PptDqsCntInvTrnTg0_p1_bits"};
      this.PptDqsCntInvTrnTg0_p1.configure(this, null, "");
      this.PptDqsCntInvTrnTg0_p1.build();
      this.default_map.add_reg(this.PptDqsCntInvTrnTg0_p1, `UVM_REG_ADDR_WIDTH'hC, "RW", 0);
		this.PptDqsCntInvTrnTg0_p1_PptDqsCntInvTrnTg0_p1 = this.PptDqsCntInvTrnTg0_p1.PptDqsCntInvTrnTg0_p1;
      this.PptDqsCntInvTrnTg1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptDqsCntInvTrnTg1_p1::type_id::create("PptDqsCntInvTrnTg1_p1",,get_full_name());
      if(this.PptDqsCntInvTrnTg1_p1.has_coverage(UVM_CVR_ALL))
      	this.PptDqsCntInvTrnTg1_p1.cg_bits.option.name = {get_name(), ".", "PptDqsCntInvTrnTg1_p1_bits"};
      this.PptDqsCntInvTrnTg1_p1.configure(this, null, "");
      this.PptDqsCntInvTrnTg1_p1.build();
      this.default_map.add_reg(this.PptDqsCntInvTrnTg1_p1, `UVM_REG_ADDR_WIDTH'hD, "RW", 0);
		this.PptDqsCntInvTrnTg1_p1_PptDqsCntInvTrnTg1_p1 = this.PptDqsCntInvTrnTg1_p1.PptDqsCntInvTrnTg1_p1;
      this.TrackingModeCntrl_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TrackingModeCntrl_p1::type_id::create("TrackingModeCntrl_p1",,get_full_name());
      if(this.TrackingModeCntrl_p1.has_coverage(UVM_CVR_ALL))
      	this.TrackingModeCntrl_p1.cg_bits.option.name = {get_name(), ".", "TrackingModeCntrl_p1_bits"};
      this.TrackingModeCntrl_p1.configure(this, null, "");
      this.TrackingModeCntrl_p1.build();
      this.default_map.add_reg(this.TrackingModeCntrl_p1, `UVM_REG_ADDR_WIDTH'hE, "RW", 0);
		this.TrackingModeCntrl_p1_EnWck2DqoSnoopTracking = this.TrackingModeCntrl_p1.EnWck2DqoSnoopTracking;
		this.EnWck2DqoSnoopTracking = this.TrackingModeCntrl_p1.EnWck2DqoSnoopTracking;
		this.TrackingModeCntrl_p1_Twck2dqoTrackingLimit = this.TrackingModeCntrl_p1.Twck2dqoTrackingLimit;
		this.Twck2dqoTrackingLimit = this.TrackingModeCntrl_p1.Twck2dqoTrackingLimit;
		this.TrackingModeCntrl_p1_ReservedTrackingModeCntrl = this.TrackingModeCntrl_p1.ReservedTrackingModeCntrl;
		this.ReservedTrackingModeCntrl = this.TrackingModeCntrl_p1.ReservedTrackingModeCntrl;
		this.TrackingModeCntrl_p1_Tdqs2dqTrackingLimit = this.TrackingModeCntrl_p1.Tdqs2dqTrackingLimit;
		this.Tdqs2dqTrackingLimit = this.TrackingModeCntrl_p1.Tdqs2dqTrackingLimit;
		this.TrackingModeCntrl_p1_DqsOscRunTimeSel = this.TrackingModeCntrl_p1.DqsOscRunTimeSel;
		this.DqsOscRunTimeSel = this.TrackingModeCntrl_p1.DqsOscRunTimeSel;
		this.TrackingModeCntrl_p1_RxDqsTrackingThreshold = this.TrackingModeCntrl_p1.RxDqsTrackingThreshold;
		this.RxDqsTrackingThreshold = this.TrackingModeCntrl_p1.RxDqsTrackingThreshold;
      this.RxClkT2UIDlyTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r0_p1::type_id::create("RxClkT2UIDlyTg0_r0_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r0_p1_bits"};
      this.RxClkT2UIDlyTg0_r0_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r0_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h10, "RW", 0);
		this.RxClkT2UIDlyTg0_r0_p1_RxClkT2UIDlyTg0_r0_p1 = this.RxClkT2UIDlyTg0_r0_p1.RxClkT2UIDlyTg0_r0_p1;
      this.RxClkT2UIDlyTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r0_p1::type_id::create("RxClkT2UIDlyTg1_r0_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r0_p1_bits"};
      this.RxClkT2UIDlyTg1_r0_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r0_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h11, "RW", 0);
		this.RxClkT2UIDlyTg1_r0_p1_RxClkT2UIDlyTg1_r0_p1 = this.RxClkT2UIDlyTg1_r0_p1.RxClkT2UIDlyTg1_r0_p1;
      this.RxClkC2UIDlyTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r0_p1::type_id::create("RxClkC2UIDlyTg0_r0_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r0_p1_bits"};
      this.RxClkC2UIDlyTg0_r0_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r0_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h12, "RW", 0);
		this.RxClkC2UIDlyTg0_r0_p1_RxClkC2UIDlyTg0_r0_p1 = this.RxClkC2UIDlyTg0_r0_p1.RxClkC2UIDlyTg0_r0_p1;
      this.RxClkC2UIDlyTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r0_p1::type_id::create("RxClkC2UIDlyTg1_r0_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r0_p1_bits"};
      this.RxClkC2UIDlyTg1_r0_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r0_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h13, "RW", 0);
		this.RxClkC2UIDlyTg1_r0_p1_RxClkC2UIDlyTg1_r0_p1 = this.RxClkC2UIDlyTg1_r0_p1.RxClkC2UIDlyTg1_r0_p1;
      this.PptWck2DqoCntInvTrnTg0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg0_p1::type_id::create("PptWck2DqoCntInvTrnTg0_p1",,get_full_name());
      if(this.PptWck2DqoCntInvTrnTg0_p1.has_coverage(UVM_CVR_ALL))
      	this.PptWck2DqoCntInvTrnTg0_p1.cg_bits.option.name = {get_name(), ".", "PptWck2DqoCntInvTrnTg0_p1_bits"};
      this.PptWck2DqoCntInvTrnTg0_p1.configure(this, null, "");
      this.PptWck2DqoCntInvTrnTg0_p1.build();
      this.default_map.add_reg(this.PptWck2DqoCntInvTrnTg0_p1, `UVM_REG_ADDR_WIDTH'h14, "RW", 0);
		this.PptWck2DqoCntInvTrnTg0_p1_PptWck2DqoCntInvTrnTg0_p1 = this.PptWck2DqoCntInvTrnTg0_p1.PptWck2DqoCntInvTrnTg0_p1;
      this.PptWck2DqoCntInvTrnTg1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PptWck2DqoCntInvTrnTg1_p1::type_id::create("PptWck2DqoCntInvTrnTg1_p1",,get_full_name());
      if(this.PptWck2DqoCntInvTrnTg1_p1.has_coverage(UVM_CVR_ALL))
      	this.PptWck2DqoCntInvTrnTg1_p1.cg_bits.option.name = {get_name(), ".", "PptWck2DqoCntInvTrnTg1_p1_bits"};
      this.PptWck2DqoCntInvTrnTg1_p1.configure(this, null, "");
      this.PptWck2DqoCntInvTrnTg1_p1.build();
      this.default_map.add_reg(this.PptWck2DqoCntInvTrnTg1_p1, `UVM_REG_ADDR_WIDTH'h15, "RW", 0);
		this.PptWck2DqoCntInvTrnTg1_p1_PptWck2DqoCntInvTrnTg1_p1 = this.PptWck2DqoCntInvTrnTg1_p1.PptWck2DqoCntInvTrnTg1_p1;
      this.TxDqsLeftEyeOffsetTg0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg0_p1::type_id::create("TxDqsLeftEyeOffsetTg0_p1",,get_full_name());
      if(this.TxDqsLeftEyeOffsetTg0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqsLeftEyeOffsetTg0_p1.cg_bits.option.name = {get_name(), ".", "TxDqsLeftEyeOffsetTg0_p1_bits"};
      this.TxDqsLeftEyeOffsetTg0_p1.configure(this, null, "");
      this.TxDqsLeftEyeOffsetTg0_p1.build();
      this.default_map.add_reg(this.TxDqsLeftEyeOffsetTg0_p1, `UVM_REG_ADDR_WIDTH'h19, "RW", 0);
		this.TxDqsLeftEyeOffsetTg0_p1_TxDqsLeftEyeOffsetTg0_p1 = this.TxDqsLeftEyeOffsetTg0_p1.TxDqsLeftEyeOffsetTg0_p1;
      this.TxDqsLeftEyeOffsetTg1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsLeftEyeOffsetTg1_p1::type_id::create("TxDqsLeftEyeOffsetTg1_p1",,get_full_name());
      if(this.TxDqsLeftEyeOffsetTg1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqsLeftEyeOffsetTg1_p1.cg_bits.option.name = {get_name(), ".", "TxDqsLeftEyeOffsetTg1_p1_bits"};
      this.TxDqsLeftEyeOffsetTg1_p1.configure(this, null, "");
      this.TxDqsLeftEyeOffsetTg1_p1.build();
      this.default_map.add_reg(this.TxDqsLeftEyeOffsetTg1_p1, `UVM_REG_ADDR_WIDTH'h1B, "RW", 0);
		this.TxDqsLeftEyeOffsetTg1_p1_TxDqsLeftEyeOffsetTg1_p1 = this.TxDqsLeftEyeOffsetTg1_p1.TxDqsLeftEyeOffsetTg1_p1;
      this.RxEnDlyTg0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg0_p1::type_id::create("RxEnDlyTg0_p1",,get_full_name());
      if(this.RxEnDlyTg0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxEnDlyTg0_p1.cg_bits.option.name = {get_name(), ".", "RxEnDlyTg0_p1_bits"};
      this.RxEnDlyTg0_p1.configure(this, null, "");
      this.RxEnDlyTg0_p1.build();
      this.default_map.add_reg(this.RxEnDlyTg0_p1, `UVM_REG_ADDR_WIDTH'h20, "RW", 0);
		this.RxEnDlyTg0_p1_RxEnDlyTg0_p1 = this.RxEnDlyTg0_p1.RxEnDlyTg0_p1;
      this.RxEnDlyTg1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxEnDlyTg1_p1::type_id::create("RxEnDlyTg1_p1",,get_full_name());
      if(this.RxEnDlyTg1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxEnDlyTg1_p1.cg_bits.option.name = {get_name(), ".", "RxEnDlyTg1_p1_bits"};
      this.RxEnDlyTg1_p1.configure(this, null, "");
      this.RxEnDlyTg1_p1.build();
      this.default_map.add_reg(this.RxEnDlyTg1_p1, `UVM_REG_ADDR_WIDTH'h21, "RW", 0);
		this.RxEnDlyTg1_p1_RxEnDlyTg1_p1 = this.RxEnDlyTg1_p1.RxEnDlyTg1_p1;
      this.TxDqsRightEyeOffsetTg0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg0_p1::type_id::create("TxDqsRightEyeOffsetTg0_p1",,get_full_name());
      if(this.TxDqsRightEyeOffsetTg0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqsRightEyeOffsetTg0_p1.cg_bits.option.name = {get_name(), ".", "TxDqsRightEyeOffsetTg0_p1_bits"};
      this.TxDqsRightEyeOffsetTg0_p1.configure(this, null, "");
      this.TxDqsRightEyeOffsetTg0_p1.build();
      this.default_map.add_reg(this.TxDqsRightEyeOffsetTg0_p1, `UVM_REG_ADDR_WIDTH'h22, "RW", 0);
		this.TxDqsRightEyeOffsetTg0_p1_TxDqsRightEyeOffsetTg0_p1 = this.TxDqsRightEyeOffsetTg0_p1.TxDqsRightEyeOffsetTg0_p1;
      this.TxDqsRightEyeOffsetTg1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsRightEyeOffsetTg1_p1::type_id::create("TxDqsRightEyeOffsetTg1_p1",,get_full_name());
      if(this.TxDqsRightEyeOffsetTg1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqsRightEyeOffsetTg1_p1.cg_bits.option.name = {get_name(), ".", "TxDqsRightEyeOffsetTg1_p1_bits"};
      this.TxDqsRightEyeOffsetTg1_p1.configure(this, null, "");
      this.TxDqsRightEyeOffsetTg1_p1.build();
      this.default_map.add_reg(this.TxDqsRightEyeOffsetTg1_p1, `UVM_REG_ADDR_WIDTH'h23, "RW", 0);
		this.TxDqsRightEyeOffsetTg1_p1_TxDqsRightEyeOffsetTg1_p1 = this.TxDqsRightEyeOffsetTg1_p1.TxDqsRightEyeOffsetTg1_p1;
      this.DqsPreambleControl_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqsPreambleControl_p1::type_id::create("DqsPreambleControl_p1",,get_full_name());
      if(this.DqsPreambleControl_p1.has_coverage(UVM_CVR_ALL))
      	this.DqsPreambleControl_p1.cg_bits.option.name = {get_name(), ".", "DqsPreambleControl_p1_bits"};
      this.DqsPreambleControl_p1.configure(this, null, "");
      this.DqsPreambleControl_p1.build();
      this.default_map.add_reg(this.DqsPreambleControl_p1, `UVM_REG_ADDR_WIDTH'h24, "RW", 0);
		this.DqsPreambleControl_p1_Reserved = this.DqsPreambleControl_p1.Reserved;
		this.Reserved = this.DqsPreambleControl_p1.Reserved;
		this.DqsPreambleControl_p1_LP4PostambleExt = this.DqsPreambleControl_p1.LP4PostambleExt;
		this.LP4PostambleExt = this.DqsPreambleControl_p1.LP4PostambleExt;
		this.DqsPreambleControl_p1_WDQSEXTENSION = this.DqsPreambleControl_p1.WDQSEXTENSION;
		this.WDQSEXTENSION = this.DqsPreambleControl_p1.WDQSEXTENSION;
		this.DqsPreambleControl_p1_WCKEXTENSION = this.DqsPreambleControl_p1.WCKEXTENSION;
		this.WCKEXTENSION = this.DqsPreambleControl_p1.WCKEXTENSION;
		this.DqsPreambleControl_p1_DqPreOeExt = this.DqsPreambleControl_p1.DqPreOeExt;
		this.DqPreOeExt = this.DqsPreambleControl_p1.DqPreOeExt;
		this.DqsPreambleControl_p1_DqPstOeExt = this.DqsPreambleControl_p1.DqPstOeExt;
		this.DqPstOeExt = this.DqsPreambleControl_p1.DqPstOeExt;
      this.DbyteRxDqsModeCntrl_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DbyteRxDqsModeCntrl_p1::type_id::create("DbyteRxDqsModeCntrl_p1",,get_full_name());
      if(this.DbyteRxDqsModeCntrl_p1.has_coverage(UVM_CVR_ALL))
      	this.DbyteRxDqsModeCntrl_p1.cg_bits.option.name = {get_name(), ".", "DbyteRxDqsModeCntrl_p1_bits"};
      this.DbyteRxDqsModeCntrl_p1.configure(this, null, "");
      this.DbyteRxDqsModeCntrl_p1.build();
      this.default_map.add_reg(this.DbyteRxDqsModeCntrl_p1, `UVM_REG_ADDR_WIDTH'h25, "RW", 0);
		this.DbyteRxDqsModeCntrl_p1_RxPostambleMode = this.DbyteRxDqsModeCntrl_p1.RxPostambleMode;
		this.RxPostambleMode = this.DbyteRxDqsModeCntrl_p1.RxPostambleMode;
		this.DbyteRxDqsModeCntrl_p1_RxPreambleMode = this.DbyteRxDqsModeCntrl_p1.RxPreambleMode;
		this.RxPreambleMode = this.DbyteRxDqsModeCntrl_p1.RxPreambleMode;
		this.DbyteRxDqsModeCntrl_p1_LPDDR5RdqsEn = this.DbyteRxDqsModeCntrl_p1.LPDDR5RdqsEn;
		this.LPDDR5RdqsEn = this.DbyteRxDqsModeCntrl_p1.LPDDR5RdqsEn;
		this.DbyteRxDqsModeCntrl_p1_LPDDR5RdqsPre = this.DbyteRxDqsModeCntrl_p1.LPDDR5RdqsPre;
		this.LPDDR5RdqsPre = this.DbyteRxDqsModeCntrl_p1.LPDDR5RdqsPre;
		this.DbyteRxDqsModeCntrl_p1_LPDDR5RdqsPst = this.DbyteRxDqsModeCntrl_p1.LPDDR5RdqsPst;
		this.LPDDR5RdqsPst = this.DbyteRxDqsModeCntrl_p1.LPDDR5RdqsPst;
		this.DbyteRxDqsModeCntrl_p1_PositionDfeInit = this.DbyteRxDqsModeCntrl_p1.PositionDfeInit;
		this.PositionDfeInit = this.DbyteRxDqsModeCntrl_p1.PositionDfeInit;
		this.DbyteRxDqsModeCntrl_p1_PositionRxPhaseUpdate = this.DbyteRxDqsModeCntrl_p1.PositionRxPhaseUpdate;
		this.PositionRxPhaseUpdate = this.DbyteRxDqsModeCntrl_p1.PositionRxPhaseUpdate;
      this.RxClkCntl1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCntl1_p1::type_id::create("RxClkCntl1_p1",,get_full_name());
      if(this.RxClkCntl1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCntl1_p1.cg_bits.option.name = {get_name(), ".", "RxClkCntl1_p1_bits"};
      this.RxClkCntl1_p1.configure(this, null, "");
      this.RxClkCntl1_p1.build();
      this.default_map.add_reg(this.RxClkCntl1_p1, `UVM_REG_ADDR_WIDTH'h27, "RW", 0);
		this.RxClkCntl1_p1_EnRxClkCor = this.RxClkCntl1_p1.EnRxClkCor;
		this.EnRxClkCor = this.RxClkCntl1_p1.EnRxClkCor;
      this.TxDqsDlyTg0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg0_p1::type_id::create("TxDqsDlyTg0_p1",,get_full_name());
      if(this.TxDqsDlyTg0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqsDlyTg0_p1.cg_bits.option.name = {get_name(), ".", "TxDqsDlyTg0_p1_bits"};
      this.TxDqsDlyTg0_p1.configure(this, null, "");
      this.TxDqsDlyTg0_p1.build();
      this.default_map.add_reg(this.TxDqsDlyTg0_p1, `UVM_REG_ADDR_WIDTH'h28, "RW", 0);
		this.TxDqsDlyTg0_p1_TxDqsDlyTg0_p1 = this.TxDqsDlyTg0_p1.TxDqsDlyTg0_p1;
      this.TxDqsDlyTg1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqsDlyTg1_p1::type_id::create("TxDqsDlyTg1_p1",,get_full_name());
      if(this.TxDqsDlyTg1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqsDlyTg1_p1.cg_bits.option.name = {get_name(), ".", "TxDqsDlyTg1_p1_bits"};
      this.TxDqsDlyTg1_p1.configure(this, null, "");
      this.TxDqsDlyTg1_p1.build();
      this.default_map.add_reg(this.TxDqsDlyTg1_p1, `UVM_REG_ADDR_WIDTH'h29, "RW", 0);
		this.TxDqsDlyTg1_p1_TxDqsDlyTg1_p1 = this.TxDqsDlyTg1_p1.TxDqsDlyTg1_p1;
      this.TxWckDlyTg0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg0_p1::type_id::create("TxWckDlyTg0_p1",,get_full_name());
      if(this.TxWckDlyTg0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxWckDlyTg0_p1.cg_bits.option.name = {get_name(), ".", "TxWckDlyTg0_p1_bits"};
      this.TxWckDlyTg0_p1.configure(this, null, "");
      this.TxWckDlyTg0_p1.build();
      this.default_map.add_reg(this.TxWckDlyTg0_p1, `UVM_REG_ADDR_WIDTH'h2A, "RW", 0);
		this.TxWckDlyTg0_p1_TxWckDlyTg0_p1 = this.TxWckDlyTg0_p1.TxWckDlyTg0_p1;
      this.TxWckDlyTg1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxWckDlyTg1_p1::type_id::create("TxWckDlyTg1_p1",,get_full_name());
      if(this.TxWckDlyTg1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxWckDlyTg1_p1.cg_bits.option.name = {get_name(), ".", "TxWckDlyTg1_p1_bits"};
      this.TxWckDlyTg1_p1.configure(this, null, "");
      this.TxWckDlyTg1_p1.build();
      this.default_map.add_reg(this.TxWckDlyTg1_p1, `UVM_REG_ADDR_WIDTH'h2B, "RW", 0);
		this.TxWckDlyTg1_p1_TxWckDlyTg1_p1 = this.TxWckDlyTg1_p1.TxWckDlyTg1_p1;
      this.RxModeCtlRxReplica_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxModeCtlRxReplica_p1::type_id::create("RxModeCtlRxReplica_p1",,get_full_name());
      if(this.RxModeCtlRxReplica_p1.has_coverage(UVM_CVR_ALL))
      	this.RxModeCtlRxReplica_p1.cg_bits.option.name = {get_name(), ".", "RxModeCtlRxReplica_p1_bits"};
      this.RxModeCtlRxReplica_p1.configure(this, null, "");
      this.RxModeCtlRxReplica_p1.build();
      this.default_map.add_reg(this.RxModeCtlRxReplica_p1, `UVM_REG_ADDR_WIDTH'h39, "RW", 0);
		this.RxModeCtlRxReplica_p1_RxModeCtlRxReplica_p1 = this.RxModeCtlRxReplica_p1.RxModeCtlRxReplica_p1;
      this.RxGainCurrAdjRxReplica_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxGainCurrAdjRxReplica_p1::type_id::create("RxGainCurrAdjRxReplica_p1",,get_full_name());
      if(this.RxGainCurrAdjRxReplica_p1.has_coverage(UVM_CVR_ALL))
      	this.RxGainCurrAdjRxReplica_p1.cg_bits.option.name = {get_name(), ".", "RxGainCurrAdjRxReplica_p1_bits"};
      this.RxGainCurrAdjRxReplica_p1.configure(this, null, "");
      this.RxGainCurrAdjRxReplica_p1.build();
      this.default_map.add_reg(this.RxGainCurrAdjRxReplica_p1, `UVM_REG_ADDR_WIDTH'h3E, "RW", 0);
		this.RxGainCurrAdjRxReplica_p1_RxGainCurrAdjRxReplica_p1 = this.RxGainCurrAdjRxReplica_p1.RxGainCurrAdjRxReplica_p1;
      this.DxRxStandbyEn_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxRxStandbyEn_p1::type_id::create("DxRxStandbyEn_p1",,get_full_name());
      if(this.DxRxStandbyEn_p1.has_coverage(UVM_CVR_ALL))
      	this.DxRxStandbyEn_p1.cg_bits.option.name = {get_name(), ".", "DxRxStandbyEn_p1_bits"};
      this.DxRxStandbyEn_p1.configure(this, null, "");
      this.DxRxStandbyEn_p1.build();
      this.default_map.add_reg(this.DxRxStandbyEn_p1, `UVM_REG_ADDR_WIDTH'h5F, "RW", 0);
		this.DxRxStandbyEn_p1_DxRxStandbyEn_p1 = this.DxRxStandbyEn_p1.DxRxStandbyEn_p1;
      this.TxDqLeftEyeOffsetTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r0_p1::type_id::create("TxDqLeftEyeOffsetTg0_r0_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r0_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r0_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r0_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h60, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r0_p1_TxDqLeftEyeOffsetTg0_r0_p1 = this.TxDqLeftEyeOffsetTg0_r0_p1.TxDqLeftEyeOffsetTg0_r0_p1;
      this.TxDqLeftEyeOffsetTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r0_p1::type_id::create("TxDqLeftEyeOffsetTg1_r0_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r0_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r0_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r0_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h61, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r0_p1_TxDqLeftEyeOffsetTg1_r0_p1 = this.TxDqLeftEyeOffsetTg1_r0_p1.TxDqLeftEyeOffsetTg1_r0_p1;
      this.TxDqRightEyeOffsetTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r0_p1::type_id::create("TxDqRightEyeOffsetTg0_r0_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r0_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r0_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r0_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h63, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r0_p1_TxDqRightEyeOffsetTg0_r0_p1 = this.TxDqRightEyeOffsetTg0_r0_p1.TxDqRightEyeOffsetTg0_r0_p1;
      this.TxDqRightEyeOffsetTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r0_p1::type_id::create("TxDqRightEyeOffsetTg1_r0_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r0_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r0_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r0_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h64, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r0_p1_TxDqRightEyeOffsetTg1_r0_p1 = this.TxDqRightEyeOffsetTg1_r0_p1.TxDqRightEyeOffsetTg1_r0_p1;
      this.RxClkTLeftEyeOffsetTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r0_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r0_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r0_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r0_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r0_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h68, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r0_p1_RxClkTLeftEyeOffsetTg0_r0_p1 = this.RxClkTLeftEyeOffsetTg0_r0_p1.RxClkTLeftEyeOffsetTg0_r0_p1;
      this.RxClkTLeftEyeOffsetTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r0_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r0_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r0_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r0_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r0_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h69, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r0_p1_RxClkTLeftEyeOffsetTg1_r0_p1 = this.RxClkTLeftEyeOffsetTg1_r0_p1.RxClkTLeftEyeOffsetTg1_r0_p1;
      this.RxClkTRightEyeOffsetTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r0_p1::type_id::create("RxClkTRightEyeOffsetTg0_r0_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r0_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r0_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r0_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h6A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r0_p1_RxClkTRightEyeOffsetTg0_r0_p1 = this.RxClkTRightEyeOffsetTg0_r0_p1.RxClkTRightEyeOffsetTg0_r0_p1;
      this.RxClkTRightEyeOffsetTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r0_p1::type_id::create("RxClkTRightEyeOffsetTg1_r0_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r0_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r0_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r0_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h6B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r0_p1_RxClkTRightEyeOffsetTg1_r0_p1 = this.RxClkTRightEyeOffsetTg1_r0_p1.RxClkTRightEyeOffsetTg1_r0_p1;
      this.RxClkCLeftEyeOffsetTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r0_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r0_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r0_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r0_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r0_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h6C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r0_p1_RxClkCLeftEyeOffsetTg0_r0_p1 = this.RxClkCLeftEyeOffsetTg0_r0_p1.RxClkCLeftEyeOffsetTg0_r0_p1;
      this.RxClkCLeftEyeOffsetTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r0_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r0_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r0_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r0_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r0_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h6D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r0_p1_RxClkCLeftEyeOffsetTg1_r0_p1 = this.RxClkCLeftEyeOffsetTg1_r0_p1.RxClkCLeftEyeOffsetTg1_r0_p1;
      this.RxClkCRightEyeOffsetTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r0_p1::type_id::create("RxClkCRightEyeOffsetTg0_r0_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r0_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r0_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r0_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h6E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r0_p1_RxClkCRightEyeOffsetTg0_r0_p1 = this.RxClkCRightEyeOffsetTg0_r0_p1.RxClkCRightEyeOffsetTg0_r0_p1;
      this.RxClkCRightEyeOffsetTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r0_p1::type_id::create("RxClkCRightEyeOffsetTg1_r0_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r0_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r0_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r0_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h6F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r0_p1_RxClkCRightEyeOffsetTg1_r0_p1 = this.RxClkCRightEyeOffsetTg1_r0_p1.RxClkCRightEyeOffsetTg1_r0_p1;
      this.RxDigStrbDlyTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r0_p1::type_id::create("RxDigStrbDlyTg0_r0_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r0_p1_bits"};
      this.RxDigStrbDlyTg0_r0_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r0_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h78, "RW", 0);
		this.RxDigStrbDlyTg0_r0_p1_RxDigStrbDlyTg0_r0_p1 = this.RxDigStrbDlyTg0_r0_p1.RxDigStrbDlyTg0_r0_p1;
      this.RxDigStrbDlyTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r0_p1::type_id::create("RxDigStrbDlyTg1_r0_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r0_p1_bits"};
      this.RxDigStrbDlyTg1_r0_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r0_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h79, "RW", 0);
		this.RxDigStrbDlyTg1_r0_p1_RxDigStrbDlyTg1_r0_p1 = this.RxDigStrbDlyTg1_r0_p1.RxDigStrbDlyTg1_r0_p1;
      this.TxDqDlyTg0_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r0_p1::type_id::create("TxDqDlyTg0_r0_p1",,get_full_name());
      if(this.TxDqDlyTg0_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r0_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r0_p1_bits"};
      this.TxDqDlyTg0_r0_p1.configure(this, null, "");
      this.TxDqDlyTg0_r0_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r0_p1, `UVM_REG_ADDR_WIDTH'h7A, "RW", 0);
		this.TxDqDlyTg0_r0_p1_TxDqDlyTg0_r0_p1 = this.TxDqDlyTg0_r0_p1.TxDqDlyTg0_r0_p1;
      this.TxDqDlyTg1_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r0_p1::type_id::create("TxDqDlyTg1_r0_p1",,get_full_name());
      if(this.TxDqDlyTg1_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r0_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r0_p1_bits"};
      this.TxDqDlyTg1_r0_p1.configure(this, null, "");
      this.TxDqDlyTg1_r0_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r0_p1, `UVM_REG_ADDR_WIDTH'h7B, "RW", 0);
		this.TxDqDlyTg1_r0_p1_TxDqDlyTg1_r0_p1 = this.TxDqDlyTg1_r0_p1.TxDqDlyTg1_r0_p1;
      this.SingleEndedMode_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_SingleEndedMode_p1::type_id::create("SingleEndedMode_p1",,get_full_name());
      if(this.SingleEndedMode_p1.has_coverage(UVM_CVR_ALL))
      	this.SingleEndedMode_p1.cg_bits.option.name = {get_name(), ".", "SingleEndedMode_p1_bits"};
      this.SingleEndedMode_p1.configure(this, null, "");
      this.SingleEndedMode_p1.build();
      this.default_map.add_reg(this.SingleEndedMode_p1, `UVM_REG_ADDR_WIDTH'h7C, "RW", 0);
		this.SingleEndedMode_p1_SingleEndedModeReserved = this.SingleEndedMode_p1.SingleEndedModeReserved;
		this.SingleEndedModeReserved = this.SingleEndedMode_p1.SingleEndedModeReserved;
		this.SingleEndedMode_p1_SingleEndedDQS = this.SingleEndedMode_p1.SingleEndedDQS;
		this.SingleEndedDQS = this.SingleEndedMode_p1.SingleEndedDQS;
		this.SingleEndedMode_p1_SingleEndedWCK = this.SingleEndedMode_p1.SingleEndedWCK;
		this.SingleEndedWCK = this.SingleEndedMode_p1.SingleEndedWCK;
      this.RxTrainPattern8BitMode_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxTrainPattern8BitMode_p1::type_id::create("RxTrainPattern8BitMode_p1",,get_full_name());
      if(this.RxTrainPattern8BitMode_p1.has_coverage(UVM_CVR_ALL))
      	this.RxTrainPattern8BitMode_p1.cg_bits.option.name = {get_name(), ".", "RxTrainPattern8BitMode_p1_bits"};
      this.RxTrainPattern8BitMode_p1.configure(this, null, "");
      this.RxTrainPattern8BitMode_p1.build();
      this.default_map.add_reg(this.RxTrainPattern8BitMode_p1, `UVM_REG_ADDR_WIDTH'hA5, "RW", 0);
		this.RxTrainPattern8BitMode_p1_RxTrainPattern8BitMode_p1 = this.RxTrainPattern8BitMode_p1.RxTrainPattern8BitMode_p1;
      this.DqRxVrefDac_r0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r0_p1::type_id::create("DqRxVrefDac_r0_p1",,get_full_name());
      if(this.DqRxVrefDac_r0_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r0_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r0_p1_bits"};
      this.DqRxVrefDac_r0_p1.configure(this, null, "");
      this.DqRxVrefDac_r0_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r0_p1, `UVM_REG_ADDR_WIDTH'hC8, "RW", 0);
		this.DqRxVrefDac_r0_p1_DqRxVrefDac_r0_p1 = this.DqRxVrefDac_r0_p1.DqRxVrefDac_r0_p1;
      this.RxDigStrbEn_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbEn_p1::type_id::create("RxDigStrbEn_p1",,get_full_name());
      if(this.RxDigStrbEn_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbEn_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbEn_p1_bits"};
      this.RxDigStrbEn_p1.configure(this, null, "");
      this.RxDigStrbEn_p1.build();
      this.default_map.add_reg(this.RxDigStrbEn_p1, `UVM_REG_ADDR_WIDTH'hFB, "RW", 0);
		this.RxDigStrbEn_p1_EnStrblssRdMode = this.RxDigStrbEn_p1.EnStrblssRdMode;
		this.EnStrblssRdMode = this.RxDigStrbEn_p1.EnStrblssRdMode;
		this.RxDigStrbEn_p1_RxReplicaPowerDownNoRDQS = this.RxDigStrbEn_p1.RxReplicaPowerDownNoRDQS;
		this.RxReplicaPowerDownNoRDQS = this.RxDigStrbEn_p1.RxReplicaPowerDownNoRDQS;
		this.RxDigStrbEn_p1_OdtDisDqs = this.RxDigStrbEn_p1.OdtDisDqs;
		this.OdtDisDqs = this.RxDigStrbEn_p1.OdtDisDqs;
      this.DxPipeEn_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DxPipeEn_p1::type_id::create("DxPipeEn_p1",,get_full_name());
      if(this.DxPipeEn_p1.has_coverage(UVM_CVR_ALL))
      	this.DxPipeEn_p1.cg_bits.option.name = {get_name(), ".", "DxPipeEn_p1_bits"};
      this.DxPipeEn_p1.configure(this, null, "");
      this.DxPipeEn_p1.build();
      this.default_map.add_reg(this.DxPipeEn_p1, `UVM_REG_ADDR_WIDTH'hFC, "RW", 0);
		this.DxPipeEn_p1_DxWrPipeEn = this.DxPipeEn_p1.DxWrPipeEn;
		this.DxWrPipeEn = this.DxPipeEn_p1.DxWrPipeEn;
		this.DxPipeEn_p1_DxRdPipeEn = this.DxPipeEn_p1.DxRdPipeEn;
		this.DxRdPipeEn = this.DxPipeEn_p1.DxRdPipeEn;
      this.PclkDCDCtrl_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCDCtrl_p1::type_id::create("PclkDCDCtrl_p1",,get_full_name());
      if(this.PclkDCDCtrl_p1.has_coverage(UVM_CVR_ALL))
      	this.PclkDCDCtrl_p1.cg_bits.option.name = {get_name(), ".", "PclkDCDCtrl_p1_bits"};
      this.PclkDCDCtrl_p1.configure(this, null, "");
      this.PclkDCDCtrl_p1.build();
      this.default_map.add_reg(this.PclkDCDCtrl_p1, `UVM_REG_ADDR_WIDTH'h100, "RW", 0);
		this.PclkDCDCtrl_p1_PclkDCDEn = this.PclkDCDCtrl_p1.PclkDCDEn;
		this.PclkDCDEn = this.PclkDCDCtrl_p1.PclkDCDEn;
		this.PclkDCDCtrl_p1_PclkDCDOffsetMode = this.PclkDCDCtrl_p1.PclkDCDOffsetMode;
		this.PclkDCDOffsetMode = this.PclkDCDCtrl_p1.PclkDCDOffsetMode;
      this.PPTTrainSetup2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PPTTrainSetup2_p1::type_id::create("PPTTrainSetup2_p1",,get_full_name());
      if(this.PPTTrainSetup2_p1.has_coverage(UVM_CVR_ALL))
      	this.PPTTrainSetup2_p1.cg_bits.option.name = {get_name(), ".", "PPTTrainSetup2_p1_bits"};
      this.PPTTrainSetup2_p1.configure(this, null, "");
      this.PPTTrainSetup2_p1.build();
      this.default_map.add_reg(this.PPTTrainSetup2_p1, `UVM_REG_ADDR_WIDTH'h102, "RW", 0);
		this.PPTTrainSetup2_p1_PPTTrainSetup2_p1 = this.PPTTrainSetup2_p1.PPTTrainSetup2_p1;
      this.DMIPinPresent_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DMIPinPresent_p1::type_id::create("DMIPinPresent_p1",,get_full_name());
      if(this.DMIPinPresent_p1.has_coverage(UVM_CVR_ALL))
      	this.DMIPinPresent_p1.cg_bits.option.name = {get_name(), ".", "DMIPinPresent_p1_bits"};
      this.DMIPinPresent_p1.configure(this, null, "");
      this.DMIPinPresent_p1.build();
      this.default_map.add_reg(this.DMIPinPresent_p1, `UVM_REG_ADDR_WIDTH'h108, "RW", 0);
		this.DMIPinPresent_p1_RdDbiEnabled = this.DMIPinPresent_p1.RdDbiEnabled;
		this.RdDbiEnabled = this.DMIPinPresent_p1.RdDbiEnabled;
      this.InhibitTxRdPtrInit_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_InhibitTxRdPtrInit_p1::type_id::create("InhibitTxRdPtrInit_p1",,get_full_name());
      if(this.InhibitTxRdPtrInit_p1.has_coverage(UVM_CVR_ALL))
      	this.InhibitTxRdPtrInit_p1.cg_bits.option.name = {get_name(), ".", "InhibitTxRdPtrInit_p1_bits"};
      this.InhibitTxRdPtrInit_p1.configure(this, null, "");
      this.InhibitTxRdPtrInit_p1.build();
      this.default_map.add_reg(this.InhibitTxRdPtrInit_p1, `UVM_REG_ADDR_WIDTH'h10B, "RW", 0);
		this.InhibitTxRdPtrInit_p1_InhibitTxRdPtrInit_p1 = this.InhibitTxRdPtrInit_p1.InhibitTxRdPtrInit_p1;
      this.RxClkT2UIDlyTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r1_p1::type_id::create("RxClkT2UIDlyTg0_r1_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r1_p1_bits"};
      this.RxClkT2UIDlyTg0_r1_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r1_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h110, "RW", 0);
		this.RxClkT2UIDlyTg0_r1_p1_RxClkT2UIDlyTg0_r1_p1 = this.RxClkT2UIDlyTg0_r1_p1.RxClkT2UIDlyTg0_r1_p1;
      this.RxClkT2UIDlyTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r1_p1::type_id::create("RxClkT2UIDlyTg1_r1_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r1_p1_bits"};
      this.RxClkT2UIDlyTg1_r1_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r1_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h111, "RW", 0);
		this.RxClkT2UIDlyTg1_r1_p1_RxClkT2UIDlyTg1_r1_p1 = this.RxClkT2UIDlyTg1_r1_p1.RxClkT2UIDlyTg1_r1_p1;
      this.RxClkC2UIDlyTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r1_p1::type_id::create("RxClkC2UIDlyTg0_r1_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r1_p1_bits"};
      this.RxClkC2UIDlyTg0_r1_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r1_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h112, "RW", 0);
		this.RxClkC2UIDlyTg0_r1_p1_RxClkC2UIDlyTg0_r1_p1 = this.RxClkC2UIDlyTg0_r1_p1.RxClkC2UIDlyTg0_r1_p1;
      this.RxClkC2UIDlyTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r1_p1::type_id::create("RxClkC2UIDlyTg1_r1_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r1_p1_bits"};
      this.RxClkC2UIDlyTg1_r1_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r1_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h113, "RW", 0);
		this.RxClkC2UIDlyTg1_r1_p1_RxClkC2UIDlyTg1_r1_p1 = this.RxClkC2UIDlyTg1_r1_p1.RxClkC2UIDlyTg1_r1_p1;
      this.RDqRDqsCntrl_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RDqRDqsCntrl_p1::type_id::create("RDqRDqsCntrl_p1",,get_full_name());
      if(this.RDqRDqsCntrl_p1.has_coverage(UVM_CVR_ALL))
      	this.RDqRDqsCntrl_p1.cg_bits.option.name = {get_name(), ".", "RDqRDqsCntrl_p1_bits"};
      this.RDqRDqsCntrl_p1.configure(this, null, "");
      this.RDqRDqsCntrl_p1.build();
      this.default_map.add_reg(this.RDqRDqsCntrl_p1, `UVM_REG_ADDR_WIDTH'h15F, "RW", 0);
		this.RDqRDqsCntrl_p1_RxPubLcdlSeed = this.RDqRDqsCntrl_p1.RxPubLcdlSeed;
		this.RxPubLcdlSeed = this.RDqRDqsCntrl_p1.RxPubLcdlSeed;
		this.RDqRDqsCntrl_p1_RDqRDqsCntrl9 = this.RDqRDqsCntrl_p1.RDqRDqsCntrl9;
		this.RDqRDqsCntrl9 = this.RDqRDqsCntrl_p1.RDqRDqsCntrl9;
		this.RDqRDqsCntrl_p1_RxPubCalModeIs1UI = this.RDqRDqsCntrl_p1.RxPubCalModeIs1UI;
		this.RxPubCalModeIs1UI = this.RDqRDqsCntrl_p1.RxPubCalModeIs1UI;
		this.RDqRDqsCntrl_p1_RxPubCntlByPState = this.RDqRDqsCntrl_p1.RxPubCntlByPState;
		this.RxPubCntlByPState = this.RDqRDqsCntrl_p1.RxPubCntlByPState;
		this.RDqRDqsCntrl_p1_RxPubRxReplicaCalModeIs1UI = this.RDqRDqsCntrl_p1.RxPubRxReplicaCalModeIs1UI;
		this.RxPubRxReplicaCalModeIs1UI = this.RDqRDqsCntrl_p1.RxPubRxReplicaCalModeIs1UI;
      this.TxDqLeftEyeOffsetTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r1_p1::type_id::create("TxDqLeftEyeOffsetTg0_r1_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r1_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r1_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r1_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h160, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r1_p1_TxDqLeftEyeOffsetTg0_r1_p1 = this.TxDqLeftEyeOffsetTg0_r1_p1.TxDqLeftEyeOffsetTg0_r1_p1;
      this.TxDqLeftEyeOffsetTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r1_p1::type_id::create("TxDqLeftEyeOffsetTg1_r1_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r1_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r1_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r1_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h161, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r1_p1_TxDqLeftEyeOffsetTg1_r1_p1 = this.TxDqLeftEyeOffsetTg1_r1_p1.TxDqLeftEyeOffsetTg1_r1_p1;
      this.TxDqRightEyeOffsetTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r1_p1::type_id::create("TxDqRightEyeOffsetTg0_r1_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r1_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r1_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r1_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h163, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r1_p1_TxDqRightEyeOffsetTg0_r1_p1 = this.TxDqRightEyeOffsetTg0_r1_p1.TxDqRightEyeOffsetTg0_r1_p1;
      this.TxDqRightEyeOffsetTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r1_p1::type_id::create("TxDqRightEyeOffsetTg1_r1_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r1_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r1_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r1_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h164, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r1_p1_TxDqRightEyeOffsetTg1_r1_p1 = this.TxDqRightEyeOffsetTg1_r1_p1.TxDqRightEyeOffsetTg1_r1_p1;
      this.RxClkTLeftEyeOffsetTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r1_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r1_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r1_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r1_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r1_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h168, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r1_p1_RxClkTLeftEyeOffsetTg0_r1_p1 = this.RxClkTLeftEyeOffsetTg0_r1_p1.RxClkTLeftEyeOffsetTg0_r1_p1;
      this.RxClkTLeftEyeOffsetTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r1_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r1_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r1_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r1_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r1_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h169, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r1_p1_RxClkTLeftEyeOffsetTg1_r1_p1 = this.RxClkTLeftEyeOffsetTg1_r1_p1.RxClkTLeftEyeOffsetTg1_r1_p1;
      this.RxClkTRightEyeOffsetTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r1_p1::type_id::create("RxClkTRightEyeOffsetTg0_r1_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r1_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r1_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r1_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h16A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r1_p1_RxClkTRightEyeOffsetTg0_r1_p1 = this.RxClkTRightEyeOffsetTg0_r1_p1.RxClkTRightEyeOffsetTg0_r1_p1;
      this.RxClkTRightEyeOffsetTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r1_p1::type_id::create("RxClkTRightEyeOffsetTg1_r1_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r1_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r1_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r1_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h16B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r1_p1_RxClkTRightEyeOffsetTg1_r1_p1 = this.RxClkTRightEyeOffsetTg1_r1_p1.RxClkTRightEyeOffsetTg1_r1_p1;
      this.RxClkCLeftEyeOffsetTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r1_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r1_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r1_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r1_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r1_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h16C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r1_p1_RxClkCLeftEyeOffsetTg0_r1_p1 = this.RxClkCLeftEyeOffsetTg0_r1_p1.RxClkCLeftEyeOffsetTg0_r1_p1;
      this.RxClkCLeftEyeOffsetTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r1_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r1_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r1_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r1_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r1_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h16D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r1_p1_RxClkCLeftEyeOffsetTg1_r1_p1 = this.RxClkCLeftEyeOffsetTg1_r1_p1.RxClkCLeftEyeOffsetTg1_r1_p1;
      this.RxClkCRightEyeOffsetTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r1_p1::type_id::create("RxClkCRightEyeOffsetTg0_r1_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r1_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r1_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r1_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h16E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r1_p1_RxClkCRightEyeOffsetTg0_r1_p1 = this.RxClkCRightEyeOffsetTg0_r1_p1.RxClkCRightEyeOffsetTg0_r1_p1;
      this.RxClkCRightEyeOffsetTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r1_p1::type_id::create("RxClkCRightEyeOffsetTg1_r1_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r1_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r1_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r1_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h16F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r1_p1_RxClkCRightEyeOffsetTg1_r1_p1 = this.RxClkCRightEyeOffsetTg1_r1_p1.RxClkCRightEyeOffsetTg1_r1_p1;
      this.RxDigStrbDlyTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r1_p1::type_id::create("RxDigStrbDlyTg0_r1_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r1_p1_bits"};
      this.RxDigStrbDlyTg0_r1_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r1_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h178, "RW", 0);
		this.RxDigStrbDlyTg0_r1_p1_RxDigStrbDlyTg0_r1_p1 = this.RxDigStrbDlyTg0_r1_p1.RxDigStrbDlyTg0_r1_p1;
      this.RxDigStrbDlyTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r1_p1::type_id::create("RxDigStrbDlyTg1_r1_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r1_p1_bits"};
      this.RxDigStrbDlyTg1_r1_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r1_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h179, "RW", 0);
		this.RxDigStrbDlyTg1_r1_p1_RxDigStrbDlyTg1_r1_p1 = this.RxDigStrbDlyTg1_r1_p1.RxDigStrbDlyTg1_r1_p1;
      this.TxDqDlyTg0_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r1_p1::type_id::create("TxDqDlyTg0_r1_p1",,get_full_name());
      if(this.TxDqDlyTg0_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r1_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r1_p1_bits"};
      this.TxDqDlyTg0_r1_p1.configure(this, null, "");
      this.TxDqDlyTg0_r1_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r1_p1, `UVM_REG_ADDR_WIDTH'h17A, "RW", 0);
		this.TxDqDlyTg0_r1_p1_TxDqDlyTg0_r1_p1 = this.TxDqDlyTg0_r1_p1.TxDqDlyTg0_r1_p1;
      this.TxDqDlyTg1_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r1_p1::type_id::create("TxDqDlyTg1_r1_p1",,get_full_name());
      if(this.TxDqDlyTg1_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r1_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r1_p1_bits"};
      this.TxDqDlyTg1_r1_p1.configure(this, null, "");
      this.TxDqDlyTg1_r1_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r1_p1, `UVM_REG_ADDR_WIDTH'h17B, "RW", 0);
		this.TxDqDlyTg1_r1_p1_TxDqDlyTg1_r1_p1 = this.TxDqDlyTg1_r1_p1.TxDqDlyTg1_r1_p1;
      this.DqRxVrefDac_r1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r1_p1::type_id::create("DqRxVrefDac_r1_p1",,get_full_name());
      if(this.DqRxVrefDac_r1_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r1_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r1_p1_bits"};
      this.DqRxVrefDac_r1_p1.configure(this, null, "");
      this.DqRxVrefDac_r1_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r1_p1, `UVM_REG_ADDR_WIDTH'h1C8, "RW", 0);
		this.DqRxVrefDac_r1_p1_DqRxVrefDac_r1_p1 = this.DqRxVrefDac_r1_p1.DqRxVrefDac_r1_p1;
      this.RxReplicaRangeVal_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaRangeVal_p1::type_id::create("RxReplicaRangeVal_p1",,get_full_name());
      if(this.RxReplicaRangeVal_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaRangeVal_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaRangeVal_p1_bits"};
      this.RxReplicaRangeVal_p1.configure(this, null, "");
      this.RxReplicaRangeVal_p1.build();
      this.default_map.add_reg(this.RxReplicaRangeVal_p1, `UVM_REG_ADDR_WIDTH'h209, "RW", 0);
		this.RxReplicaRangeVal_p1_RxReplicaShortCalRangeA = this.RxReplicaRangeVal_p1.RxReplicaShortCalRangeA;
		this.RxReplicaShortCalRangeA = this.RxReplicaRangeVal_p1.RxReplicaShortCalRangeA;
		this.RxReplicaRangeVal_p1_RxReplicaShortCalRangeB = this.RxReplicaRangeVal_p1.RxReplicaShortCalRangeB;
		this.RxReplicaShortCalRangeB = this.RxReplicaRangeVal_p1.RxReplicaShortCalRangeB;
      this.RxReplicaCtl04_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl04_p1::type_id::create("RxReplicaCtl04_p1",,get_full_name());
      if(this.RxReplicaCtl04_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaCtl04_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaCtl04_p1_bits"};
      this.RxReplicaCtl04_p1.configure(this, null, "");
      this.RxReplicaCtl04_p1.build();
      this.default_map.add_reg(this.RxReplicaCtl04_p1, `UVM_REG_ADDR_WIDTH'h20F, "RW", 0);
		this.RxReplicaCtl04_p1_RxReplicaTrackEn = this.RxReplicaCtl04_p1.RxReplicaTrackEn;
		this.RxReplicaTrackEn = this.RxReplicaCtl04_p1.RxReplicaTrackEn;
		this.RxReplicaCtl04_p1_RxReplicaLongCal = this.RxReplicaCtl04_p1.RxReplicaLongCal;
		this.RxReplicaLongCal = this.RxReplicaCtl04_p1.RxReplicaLongCal;
		this.RxReplicaCtl04_p1_RxReplicaStride = this.RxReplicaCtl04_p1.RxReplicaStride;
		this.RxReplicaStride = this.RxReplicaCtl04_p1.RxReplicaStride;
		this.RxReplicaCtl04_p1_RxReplicaStandby = this.RxReplicaCtl04_p1.RxReplicaStandby;
		this.RxReplicaStandby = this.RxReplicaCtl04_p1.RxReplicaStandby;
		this.RxReplicaCtl04_p1_RxReplicaPDenFSM = this.RxReplicaCtl04_p1.RxReplicaPDenFSM;
		this.RxReplicaPDenFSM = this.RxReplicaCtl04_p1.RxReplicaPDenFSM;
		this.RxReplicaCtl04_p1_RxReplicaPDRecoverytime = this.RxReplicaCtl04_p1.RxReplicaPDRecoverytime;
		this.RxReplicaPDRecoverytime = this.RxReplicaCtl04_p1.RxReplicaPDRecoverytime;
      this.RxClkT2UIDlyTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r2_p1::type_id::create("RxClkT2UIDlyTg0_r2_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r2_p1_bits"};
      this.RxClkT2UIDlyTg0_r2_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r2_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h210, "RW", 0);
		this.RxClkT2UIDlyTg0_r2_p1_RxClkT2UIDlyTg0_r2_p1 = this.RxClkT2UIDlyTg0_r2_p1.RxClkT2UIDlyTg0_r2_p1;
      this.RxClkT2UIDlyTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r2_p1::type_id::create("RxClkT2UIDlyTg1_r2_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r2_p1_bits"};
      this.RxClkT2UIDlyTg1_r2_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r2_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h211, "RW", 0);
		this.RxClkT2UIDlyTg1_r2_p1_RxClkT2UIDlyTg1_r2_p1 = this.RxClkT2UIDlyTg1_r2_p1.RxClkT2UIDlyTg1_r2_p1;
      this.RxClkC2UIDlyTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r2_p1::type_id::create("RxClkC2UIDlyTg0_r2_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r2_p1_bits"};
      this.RxClkC2UIDlyTg0_r2_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r2_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h212, "RW", 0);
		this.RxClkC2UIDlyTg0_r2_p1_RxClkC2UIDlyTg0_r2_p1 = this.RxClkC2UIDlyTg0_r2_p1.RxClkC2UIDlyTg0_r2_p1;
      this.RxClkC2UIDlyTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r2_p1::type_id::create("RxClkC2UIDlyTg1_r2_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r2_p1_bits"};
      this.RxClkC2UIDlyTg1_r2_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r2_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h213, "RW", 0);
		this.RxClkC2UIDlyTg1_r2_p1_RxClkC2UIDlyTg1_r2_p1 = this.RxClkC2UIDlyTg1_r2_p1.RxClkC2UIDlyTg1_r2_p1;
      this.TxDqLeftEyeOffsetTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r2_p1::type_id::create("TxDqLeftEyeOffsetTg0_r2_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r2_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r2_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r2_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h260, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r2_p1_TxDqLeftEyeOffsetTg0_r2_p1 = this.TxDqLeftEyeOffsetTg0_r2_p1.TxDqLeftEyeOffsetTg0_r2_p1;
      this.TxDqLeftEyeOffsetTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r2_p1::type_id::create("TxDqLeftEyeOffsetTg1_r2_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r2_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r2_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r2_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h261, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r2_p1_TxDqLeftEyeOffsetTg1_r2_p1 = this.TxDqLeftEyeOffsetTg1_r2_p1.TxDqLeftEyeOffsetTg1_r2_p1;
      this.TxDqRightEyeOffsetTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r2_p1::type_id::create("TxDqRightEyeOffsetTg0_r2_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r2_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r2_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r2_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h263, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r2_p1_TxDqRightEyeOffsetTg0_r2_p1 = this.TxDqRightEyeOffsetTg0_r2_p1.TxDqRightEyeOffsetTg0_r2_p1;
      this.TxDqRightEyeOffsetTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r2_p1::type_id::create("TxDqRightEyeOffsetTg1_r2_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r2_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r2_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r2_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h264, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r2_p1_TxDqRightEyeOffsetTg1_r2_p1 = this.TxDqRightEyeOffsetTg1_r2_p1.TxDqRightEyeOffsetTg1_r2_p1;
      this.RxClkTLeftEyeOffsetTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r2_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r2_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r2_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r2_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r2_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h268, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r2_p1_RxClkTLeftEyeOffsetTg0_r2_p1 = this.RxClkTLeftEyeOffsetTg0_r2_p1.RxClkTLeftEyeOffsetTg0_r2_p1;
      this.RxClkTLeftEyeOffsetTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r2_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r2_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r2_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r2_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r2_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h269, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r2_p1_RxClkTLeftEyeOffsetTg1_r2_p1 = this.RxClkTLeftEyeOffsetTg1_r2_p1.RxClkTLeftEyeOffsetTg1_r2_p1;
      this.RxClkTRightEyeOffsetTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r2_p1::type_id::create("RxClkTRightEyeOffsetTg0_r2_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r2_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r2_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r2_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h26A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r2_p1_RxClkTRightEyeOffsetTg0_r2_p1 = this.RxClkTRightEyeOffsetTg0_r2_p1.RxClkTRightEyeOffsetTg0_r2_p1;
      this.RxClkTRightEyeOffsetTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r2_p1::type_id::create("RxClkTRightEyeOffsetTg1_r2_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r2_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r2_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r2_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h26B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r2_p1_RxClkTRightEyeOffsetTg1_r2_p1 = this.RxClkTRightEyeOffsetTg1_r2_p1.RxClkTRightEyeOffsetTg1_r2_p1;
      this.RxClkCLeftEyeOffsetTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r2_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r2_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r2_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r2_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r2_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h26C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r2_p1_RxClkCLeftEyeOffsetTg0_r2_p1 = this.RxClkCLeftEyeOffsetTg0_r2_p1.RxClkCLeftEyeOffsetTg0_r2_p1;
      this.RxClkCLeftEyeOffsetTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r2_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r2_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r2_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r2_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r2_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h26D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r2_p1_RxClkCLeftEyeOffsetTg1_r2_p1 = this.RxClkCLeftEyeOffsetTg1_r2_p1.RxClkCLeftEyeOffsetTg1_r2_p1;
      this.RxClkCRightEyeOffsetTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r2_p1::type_id::create("RxClkCRightEyeOffsetTg0_r2_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r2_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r2_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r2_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h26E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r2_p1_RxClkCRightEyeOffsetTg0_r2_p1 = this.RxClkCRightEyeOffsetTg0_r2_p1.RxClkCRightEyeOffsetTg0_r2_p1;
      this.RxClkCRightEyeOffsetTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r2_p1::type_id::create("RxClkCRightEyeOffsetTg1_r2_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r2_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r2_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r2_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h26F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r2_p1_RxClkCRightEyeOffsetTg1_r2_p1 = this.RxClkCRightEyeOffsetTg1_r2_p1.RxClkCRightEyeOffsetTg1_r2_p1;
      this.RxDigStrbDlyTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r2_p1::type_id::create("RxDigStrbDlyTg0_r2_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r2_p1_bits"};
      this.RxDigStrbDlyTg0_r2_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r2_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h278, "RW", 0);
		this.RxDigStrbDlyTg0_r2_p1_RxDigStrbDlyTg0_r2_p1 = this.RxDigStrbDlyTg0_r2_p1.RxDigStrbDlyTg0_r2_p1;
      this.RxDigStrbDlyTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r2_p1::type_id::create("RxDigStrbDlyTg1_r2_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r2_p1_bits"};
      this.RxDigStrbDlyTg1_r2_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r2_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h279, "RW", 0);
		this.RxDigStrbDlyTg1_r2_p1_RxDigStrbDlyTg1_r2_p1 = this.RxDigStrbDlyTg1_r2_p1.RxDigStrbDlyTg1_r2_p1;
      this.TxDqDlyTg0_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r2_p1::type_id::create("TxDqDlyTg0_r2_p1",,get_full_name());
      if(this.TxDqDlyTg0_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r2_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r2_p1_bits"};
      this.TxDqDlyTg0_r2_p1.configure(this, null, "");
      this.TxDqDlyTg0_r2_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r2_p1, `UVM_REG_ADDR_WIDTH'h27A, "RW", 0);
		this.TxDqDlyTg0_r2_p1_TxDqDlyTg0_r2_p1 = this.TxDqDlyTg0_r2_p1.TxDqDlyTg0_r2_p1;
      this.TxDqDlyTg1_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r2_p1::type_id::create("TxDqDlyTg1_r2_p1",,get_full_name());
      if(this.TxDqDlyTg1_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r2_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r2_p1_bits"};
      this.TxDqDlyTg1_r2_p1.configure(this, null, "");
      this.TxDqDlyTg1_r2_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r2_p1, `UVM_REG_ADDR_WIDTH'h27B, "RW", 0);
		this.TxDqDlyTg1_r2_p1_TxDqDlyTg1_r2_p1 = this.TxDqDlyTg1_r2_p1.TxDqDlyTg1_r2_p1;
      this.RxReplicaPathPhase0_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase0_p1::type_id::create("RxReplicaPathPhase0_p1",,get_full_name());
      if(this.RxReplicaPathPhase0_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaPathPhase0_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaPathPhase0_p1_bits"};
      this.RxReplicaPathPhase0_p1.configure(this, null, "");
      this.RxReplicaPathPhase0_p1.build();
      this.default_map.add_reg(this.RxReplicaPathPhase0_p1, `UVM_REG_ADDR_WIDTH'h2A0, "RW", 0);
		this.RxReplicaPathPhase0_p1_RxReplicaPathPhase0_p1 = this.RxReplicaPathPhase0_p1.RxReplicaPathPhase0_p1;
      this.RxReplicaPathPhase1_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase1_p1::type_id::create("RxReplicaPathPhase1_p1",,get_full_name());
      if(this.RxReplicaPathPhase1_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaPathPhase1_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaPathPhase1_p1_bits"};
      this.RxReplicaPathPhase1_p1.configure(this, null, "");
      this.RxReplicaPathPhase1_p1.build();
      this.default_map.add_reg(this.RxReplicaPathPhase1_p1, `UVM_REG_ADDR_WIDTH'h2A1, "RW", 0);
		this.RxReplicaPathPhase1_p1_RxReplicaPathPhase1_p1 = this.RxReplicaPathPhase1_p1.RxReplicaPathPhase1_p1;
      this.RxReplicaPathPhase2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase2_p1::type_id::create("RxReplicaPathPhase2_p1",,get_full_name());
      if(this.RxReplicaPathPhase2_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaPathPhase2_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaPathPhase2_p1_bits"};
      this.RxReplicaPathPhase2_p1.configure(this, null, "");
      this.RxReplicaPathPhase2_p1.build();
      this.default_map.add_reg(this.RxReplicaPathPhase2_p1, `UVM_REG_ADDR_WIDTH'h2A2, "RW", 0);
		this.RxReplicaPathPhase2_p1_RxReplicaPathPhase2_p1 = this.RxReplicaPathPhase2_p1.RxReplicaPathPhase2_p1;
      this.RxReplicaPathPhase3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase3_p1::type_id::create("RxReplicaPathPhase3_p1",,get_full_name());
      if(this.RxReplicaPathPhase3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaPathPhase3_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaPathPhase3_p1_bits"};
      this.RxReplicaPathPhase3_p1.configure(this, null, "");
      this.RxReplicaPathPhase3_p1.build();
      this.default_map.add_reg(this.RxReplicaPathPhase3_p1, `UVM_REG_ADDR_WIDTH'h2A3, "RW", 0);
		this.RxReplicaPathPhase3_p1_RxReplicaPathPhase3_p1 = this.RxReplicaPathPhase3_p1.RxReplicaPathPhase3_p1;
      this.RxReplicaPathPhase4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaPathPhase4_p1::type_id::create("RxReplicaPathPhase4_p1",,get_full_name());
      if(this.RxReplicaPathPhase4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaPathPhase4_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaPathPhase4_p1_bits"};
      this.RxReplicaPathPhase4_p1.configure(this, null, "");
      this.RxReplicaPathPhase4_p1.build();
      this.default_map.add_reg(this.RxReplicaPathPhase4_p1, `UVM_REG_ADDR_WIDTH'h2A4, "RW", 0);
		this.RxReplicaPathPhase4_p1_RxReplicaPathPhase4_p1 = this.RxReplicaPathPhase4_p1.RxReplicaPathPhase4_p1;
      this.RxReplicaCtl01_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl01_p1::type_id::create("RxReplicaCtl01_p1",,get_full_name());
      if(this.RxReplicaCtl01_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaCtl01_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaCtl01_p1_bits"};
      this.RxReplicaCtl01_p1.configure(this, null, "");
      this.RxReplicaCtl01_p1.build();
      this.default_map.add_reg(this.RxReplicaCtl01_p1, `UVM_REG_ADDR_WIDTH'h2AD, "RW", 0);
		this.RxReplicaCtl01_p1_RxReplicaSelPathPhase = this.RxReplicaCtl01_p1.RxReplicaSelPathPhase;
		this.RxReplicaSelPathPhase = this.RxReplicaCtl01_p1.RxReplicaSelPathPhase;
      this.RxReplicaCtl02_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl02_p1::type_id::create("RxReplicaCtl02_p1",,get_full_name());
      if(this.RxReplicaCtl02_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaCtl02_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaCtl02_p1_bits"};
      this.RxReplicaCtl02_p1.configure(this, null, "");
      this.RxReplicaCtl02_p1.build();
      this.default_map.add_reg(this.RxReplicaCtl02_p1, `UVM_REG_ADDR_WIDTH'h2AE, "RW", 0);
		this.RxReplicaCtl02_p1_RxReplicaDiffLimit = this.RxReplicaCtl02_p1.RxReplicaDiffLimit;
		this.RxReplicaDiffLimit = this.RxReplicaCtl02_p1.RxReplicaDiffLimit;
      this.RxReplicaCtl03_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxReplicaCtl03_p1::type_id::create("RxReplicaCtl03_p1",,get_full_name());
      if(this.RxReplicaCtl03_p1.has_coverage(UVM_CVR_ALL))
      	this.RxReplicaCtl03_p1.cg_bits.option.name = {get_name(), ".", "RxReplicaCtl03_p1_bits"};
      this.RxReplicaCtl03_p1.configure(this, null, "");
      this.RxReplicaCtl03_p1.build();
      this.default_map.add_reg(this.RxReplicaCtl03_p1, `UVM_REG_ADDR_WIDTH'h2AF, "RW", 0);
		this.RxReplicaCtl03_p1_RxReplicaRatioTrn = this.RxReplicaCtl03_p1.RxReplicaRatioTrn;
		this.RxReplicaRatioTrn = this.RxReplicaCtl03_p1.RxReplicaRatioTrn;
      this.DqRxVrefDac_r2_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r2_p1::type_id::create("DqRxVrefDac_r2_p1",,get_full_name());
      if(this.DqRxVrefDac_r2_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r2_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r2_p1_bits"};
      this.DqRxVrefDac_r2_p1.configure(this, null, "");
      this.DqRxVrefDac_r2_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r2_p1, `UVM_REG_ADDR_WIDTH'h2C8, "RW", 0);
		this.DqRxVrefDac_r2_p1_DqRxVrefDac_r2_p1 = this.DqRxVrefDac_r2_p1.DqRxVrefDac_r2_p1;
      this.RxClkT2UIDlyTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r3_p1::type_id::create("RxClkT2UIDlyTg0_r3_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r3_p1_bits"};
      this.RxClkT2UIDlyTg0_r3_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r3_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h310, "RW", 0);
		this.RxClkT2UIDlyTg0_r3_p1_RxClkT2UIDlyTg0_r3_p1 = this.RxClkT2UIDlyTg0_r3_p1.RxClkT2UIDlyTg0_r3_p1;
      this.RxClkT2UIDlyTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r3_p1::type_id::create("RxClkT2UIDlyTg1_r3_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r3_p1_bits"};
      this.RxClkT2UIDlyTg1_r3_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r3_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h311, "RW", 0);
		this.RxClkT2UIDlyTg1_r3_p1_RxClkT2UIDlyTg1_r3_p1 = this.RxClkT2UIDlyTg1_r3_p1.RxClkT2UIDlyTg1_r3_p1;
      this.RxClkC2UIDlyTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r3_p1::type_id::create("RxClkC2UIDlyTg0_r3_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r3_p1_bits"};
      this.RxClkC2UIDlyTg0_r3_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r3_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h312, "RW", 0);
		this.RxClkC2UIDlyTg0_r3_p1_RxClkC2UIDlyTg0_r3_p1 = this.RxClkC2UIDlyTg0_r3_p1.RxClkC2UIDlyTg0_r3_p1;
      this.RxClkC2UIDlyTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r3_p1::type_id::create("RxClkC2UIDlyTg1_r3_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r3_p1_bits"};
      this.RxClkC2UIDlyTg1_r3_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r3_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h313, "RW", 0);
		this.RxClkC2UIDlyTg1_r3_p1_RxClkC2UIDlyTg1_r3_p1 = this.RxClkC2UIDlyTg1_r3_p1.RxClkC2UIDlyTg1_r3_p1;
      this.TxDqLeftEyeOffsetTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r3_p1::type_id::create("TxDqLeftEyeOffsetTg0_r3_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r3_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r3_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r3_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h360, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r3_p1_TxDqLeftEyeOffsetTg0_r3_p1 = this.TxDqLeftEyeOffsetTg0_r3_p1.TxDqLeftEyeOffsetTg0_r3_p1;
      this.TxDqLeftEyeOffsetTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r3_p1::type_id::create("TxDqLeftEyeOffsetTg1_r3_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r3_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r3_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r3_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h361, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r3_p1_TxDqLeftEyeOffsetTg1_r3_p1 = this.TxDqLeftEyeOffsetTg1_r3_p1.TxDqLeftEyeOffsetTg1_r3_p1;
      this.TxDqRightEyeOffsetTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r3_p1::type_id::create("TxDqRightEyeOffsetTg0_r3_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r3_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r3_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r3_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h363, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r3_p1_TxDqRightEyeOffsetTg0_r3_p1 = this.TxDqRightEyeOffsetTg0_r3_p1.TxDqRightEyeOffsetTg0_r3_p1;
      this.TxDqRightEyeOffsetTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r3_p1::type_id::create("TxDqRightEyeOffsetTg1_r3_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r3_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r3_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r3_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h364, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r3_p1_TxDqRightEyeOffsetTg1_r3_p1 = this.TxDqRightEyeOffsetTg1_r3_p1.TxDqRightEyeOffsetTg1_r3_p1;
      this.RxClkTLeftEyeOffsetTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r3_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r3_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r3_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r3_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r3_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h368, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r3_p1_RxClkTLeftEyeOffsetTg0_r3_p1 = this.RxClkTLeftEyeOffsetTg0_r3_p1.RxClkTLeftEyeOffsetTg0_r3_p1;
      this.RxClkTLeftEyeOffsetTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r3_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r3_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r3_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r3_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r3_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h369, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r3_p1_RxClkTLeftEyeOffsetTg1_r3_p1 = this.RxClkTLeftEyeOffsetTg1_r3_p1.RxClkTLeftEyeOffsetTg1_r3_p1;
      this.RxClkTRightEyeOffsetTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r3_p1::type_id::create("RxClkTRightEyeOffsetTg0_r3_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r3_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r3_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r3_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h36A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r3_p1_RxClkTRightEyeOffsetTg0_r3_p1 = this.RxClkTRightEyeOffsetTg0_r3_p1.RxClkTRightEyeOffsetTg0_r3_p1;
      this.RxClkTRightEyeOffsetTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r3_p1::type_id::create("RxClkTRightEyeOffsetTg1_r3_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r3_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r3_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r3_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h36B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r3_p1_RxClkTRightEyeOffsetTg1_r3_p1 = this.RxClkTRightEyeOffsetTg1_r3_p1.RxClkTRightEyeOffsetTg1_r3_p1;
      this.RxClkCLeftEyeOffsetTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r3_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r3_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r3_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r3_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r3_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h36C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r3_p1_RxClkCLeftEyeOffsetTg0_r3_p1 = this.RxClkCLeftEyeOffsetTg0_r3_p1.RxClkCLeftEyeOffsetTg0_r3_p1;
      this.RxClkCLeftEyeOffsetTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r3_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r3_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r3_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r3_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r3_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h36D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r3_p1_RxClkCLeftEyeOffsetTg1_r3_p1 = this.RxClkCLeftEyeOffsetTg1_r3_p1.RxClkCLeftEyeOffsetTg1_r3_p1;
      this.RxClkCRightEyeOffsetTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r3_p1::type_id::create("RxClkCRightEyeOffsetTg0_r3_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r3_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r3_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r3_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h36E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r3_p1_RxClkCRightEyeOffsetTg0_r3_p1 = this.RxClkCRightEyeOffsetTg0_r3_p1.RxClkCRightEyeOffsetTg0_r3_p1;
      this.RxClkCRightEyeOffsetTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r3_p1::type_id::create("RxClkCRightEyeOffsetTg1_r3_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r3_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r3_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r3_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h36F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r3_p1_RxClkCRightEyeOffsetTg1_r3_p1 = this.RxClkCRightEyeOffsetTg1_r3_p1.RxClkCRightEyeOffsetTg1_r3_p1;
      this.RxDigStrbDlyTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r3_p1::type_id::create("RxDigStrbDlyTg0_r3_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r3_p1_bits"};
      this.RxDigStrbDlyTg0_r3_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r3_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h378, "RW", 0);
		this.RxDigStrbDlyTg0_r3_p1_RxDigStrbDlyTg0_r3_p1 = this.RxDigStrbDlyTg0_r3_p1.RxDigStrbDlyTg0_r3_p1;
      this.RxDigStrbDlyTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r3_p1::type_id::create("RxDigStrbDlyTg1_r3_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r3_p1_bits"};
      this.RxDigStrbDlyTg1_r3_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r3_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h379, "RW", 0);
		this.RxDigStrbDlyTg1_r3_p1_RxDigStrbDlyTg1_r3_p1 = this.RxDigStrbDlyTg1_r3_p1.RxDigStrbDlyTg1_r3_p1;
      this.TxDqDlyTg0_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r3_p1::type_id::create("TxDqDlyTg0_r3_p1",,get_full_name());
      if(this.TxDqDlyTg0_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r3_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r3_p1_bits"};
      this.TxDqDlyTg0_r3_p1.configure(this, null, "");
      this.TxDqDlyTg0_r3_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r3_p1, `UVM_REG_ADDR_WIDTH'h37A, "RW", 0);
		this.TxDqDlyTg0_r3_p1_TxDqDlyTg0_r3_p1 = this.TxDqDlyTg0_r3_p1.TxDqDlyTg0_r3_p1;
      this.TxDqDlyTg1_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r3_p1::type_id::create("TxDqDlyTg1_r3_p1",,get_full_name());
      if(this.TxDqDlyTg1_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r3_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r3_p1_bits"};
      this.TxDqDlyTg1_r3_p1.configure(this, null, "");
      this.TxDqDlyTg1_r3_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r3_p1, `UVM_REG_ADDR_WIDTH'h37B, "RW", 0);
		this.TxDqDlyTg1_r3_p1_TxDqDlyTg1_r3_p1 = this.TxDqDlyTg1_r3_p1.TxDqDlyTg1_r3_p1;
      this.DqRxVrefDac_r3_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r3_p1::type_id::create("DqRxVrefDac_r3_p1",,get_full_name());
      if(this.DqRxVrefDac_r3_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r3_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r3_p1_bits"};
      this.DqRxVrefDac_r3_p1.configure(this, null, "");
      this.DqRxVrefDac_r3_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r3_p1, `UVM_REG_ADDR_WIDTH'h3C8, "RW", 0);
		this.DqRxVrefDac_r3_p1_DqRxVrefDac_r3_p1 = this.DqRxVrefDac_r3_p1.DqRxVrefDac_r3_p1;
      this.RxClkT2UIDlyTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r4_p1::type_id::create("RxClkT2UIDlyTg0_r4_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r4_p1_bits"};
      this.RxClkT2UIDlyTg0_r4_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r4_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h410, "RW", 0);
		this.RxClkT2UIDlyTg0_r4_p1_RxClkT2UIDlyTg0_r4_p1 = this.RxClkT2UIDlyTg0_r4_p1.RxClkT2UIDlyTg0_r4_p1;
      this.RxClkT2UIDlyTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r4_p1::type_id::create("RxClkT2UIDlyTg1_r4_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r4_p1_bits"};
      this.RxClkT2UIDlyTg1_r4_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r4_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h411, "RW", 0);
		this.RxClkT2UIDlyTg1_r4_p1_RxClkT2UIDlyTg1_r4_p1 = this.RxClkT2UIDlyTg1_r4_p1.RxClkT2UIDlyTg1_r4_p1;
      this.RxClkC2UIDlyTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r4_p1::type_id::create("RxClkC2UIDlyTg0_r4_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r4_p1_bits"};
      this.RxClkC2UIDlyTg0_r4_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r4_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h412, "RW", 0);
		this.RxClkC2UIDlyTg0_r4_p1_RxClkC2UIDlyTg0_r4_p1 = this.RxClkC2UIDlyTg0_r4_p1.RxClkC2UIDlyTg0_r4_p1;
      this.RxClkC2UIDlyTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r4_p1::type_id::create("RxClkC2UIDlyTg1_r4_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r4_p1_bits"};
      this.RxClkC2UIDlyTg1_r4_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r4_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h413, "RW", 0);
		this.RxClkC2UIDlyTg1_r4_p1_RxClkC2UIDlyTg1_r4_p1 = this.RxClkC2UIDlyTg1_r4_p1.RxClkC2UIDlyTg1_r4_p1;
      this.TxDqLeftEyeOffsetTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r4_p1::type_id::create("TxDqLeftEyeOffsetTg0_r4_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r4_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r4_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r4_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h460, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r4_p1_TxDqLeftEyeOffsetTg0_r4_p1 = this.TxDqLeftEyeOffsetTg0_r4_p1.TxDqLeftEyeOffsetTg0_r4_p1;
      this.TxDqLeftEyeOffsetTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r4_p1::type_id::create("TxDqLeftEyeOffsetTg1_r4_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r4_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r4_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r4_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h461, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r4_p1_TxDqLeftEyeOffsetTg1_r4_p1 = this.TxDqLeftEyeOffsetTg1_r4_p1.TxDqLeftEyeOffsetTg1_r4_p1;
      this.TxDqRightEyeOffsetTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r4_p1::type_id::create("TxDqRightEyeOffsetTg0_r4_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r4_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r4_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r4_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h463, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r4_p1_TxDqRightEyeOffsetTg0_r4_p1 = this.TxDqRightEyeOffsetTg0_r4_p1.TxDqRightEyeOffsetTg0_r4_p1;
      this.TxDqRightEyeOffsetTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r4_p1::type_id::create("TxDqRightEyeOffsetTg1_r4_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r4_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r4_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r4_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h464, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r4_p1_TxDqRightEyeOffsetTg1_r4_p1 = this.TxDqRightEyeOffsetTg1_r4_p1.TxDqRightEyeOffsetTg1_r4_p1;
      this.RxClkTLeftEyeOffsetTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r4_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r4_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r4_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r4_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r4_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h468, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r4_p1_RxClkTLeftEyeOffsetTg0_r4_p1 = this.RxClkTLeftEyeOffsetTg0_r4_p1.RxClkTLeftEyeOffsetTg0_r4_p1;
      this.RxClkTLeftEyeOffsetTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r4_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r4_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r4_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r4_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r4_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h469, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r4_p1_RxClkTLeftEyeOffsetTg1_r4_p1 = this.RxClkTLeftEyeOffsetTg1_r4_p1.RxClkTLeftEyeOffsetTg1_r4_p1;
      this.RxClkTRightEyeOffsetTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r4_p1::type_id::create("RxClkTRightEyeOffsetTg0_r4_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r4_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r4_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r4_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h46A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r4_p1_RxClkTRightEyeOffsetTg0_r4_p1 = this.RxClkTRightEyeOffsetTg0_r4_p1.RxClkTRightEyeOffsetTg0_r4_p1;
      this.RxClkTRightEyeOffsetTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r4_p1::type_id::create("RxClkTRightEyeOffsetTg1_r4_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r4_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r4_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r4_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h46B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r4_p1_RxClkTRightEyeOffsetTg1_r4_p1 = this.RxClkTRightEyeOffsetTg1_r4_p1.RxClkTRightEyeOffsetTg1_r4_p1;
      this.RxClkCLeftEyeOffsetTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r4_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r4_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r4_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r4_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r4_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h46C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r4_p1_RxClkCLeftEyeOffsetTg0_r4_p1 = this.RxClkCLeftEyeOffsetTg0_r4_p1.RxClkCLeftEyeOffsetTg0_r4_p1;
      this.RxClkCLeftEyeOffsetTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r4_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r4_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r4_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r4_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r4_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h46D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r4_p1_RxClkCLeftEyeOffsetTg1_r4_p1 = this.RxClkCLeftEyeOffsetTg1_r4_p1.RxClkCLeftEyeOffsetTg1_r4_p1;
      this.RxClkCRightEyeOffsetTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r4_p1::type_id::create("RxClkCRightEyeOffsetTg0_r4_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r4_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r4_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r4_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h46E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r4_p1_RxClkCRightEyeOffsetTg0_r4_p1 = this.RxClkCRightEyeOffsetTg0_r4_p1.RxClkCRightEyeOffsetTg0_r4_p1;
      this.RxClkCRightEyeOffsetTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r4_p1::type_id::create("RxClkCRightEyeOffsetTg1_r4_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r4_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r4_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r4_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h46F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r4_p1_RxClkCRightEyeOffsetTg1_r4_p1 = this.RxClkCRightEyeOffsetTg1_r4_p1.RxClkCRightEyeOffsetTg1_r4_p1;
      this.RxDigStrbDlyTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r4_p1::type_id::create("RxDigStrbDlyTg0_r4_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r4_p1_bits"};
      this.RxDigStrbDlyTg0_r4_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r4_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h478, "RW", 0);
		this.RxDigStrbDlyTg0_r4_p1_RxDigStrbDlyTg0_r4_p1 = this.RxDigStrbDlyTg0_r4_p1.RxDigStrbDlyTg0_r4_p1;
      this.RxDigStrbDlyTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r4_p1::type_id::create("RxDigStrbDlyTg1_r4_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r4_p1_bits"};
      this.RxDigStrbDlyTg1_r4_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r4_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h479, "RW", 0);
		this.RxDigStrbDlyTg1_r4_p1_RxDigStrbDlyTg1_r4_p1 = this.RxDigStrbDlyTg1_r4_p1.RxDigStrbDlyTg1_r4_p1;
      this.TxDqDlyTg0_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r4_p1::type_id::create("TxDqDlyTg0_r4_p1",,get_full_name());
      if(this.TxDqDlyTg0_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r4_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r4_p1_bits"};
      this.TxDqDlyTg0_r4_p1.configure(this, null, "");
      this.TxDqDlyTg0_r4_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r4_p1, `UVM_REG_ADDR_WIDTH'h47A, "RW", 0);
		this.TxDqDlyTg0_r4_p1_TxDqDlyTg0_r4_p1 = this.TxDqDlyTg0_r4_p1.TxDqDlyTg0_r4_p1;
      this.TxDqDlyTg1_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r4_p1::type_id::create("TxDqDlyTg1_r4_p1",,get_full_name());
      if(this.TxDqDlyTg1_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r4_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r4_p1_bits"};
      this.TxDqDlyTg1_r4_p1.configure(this, null, "");
      this.TxDqDlyTg1_r4_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r4_p1, `UVM_REG_ADDR_WIDTH'h47B, "RW", 0);
		this.TxDqDlyTg1_r4_p1_TxDqDlyTg1_r4_p1 = this.TxDqDlyTg1_r4_p1.TxDqDlyTg1_r4_p1;
      this.DqRxVrefDac_r4_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r4_p1::type_id::create("DqRxVrefDac_r4_p1",,get_full_name());
      if(this.DqRxVrefDac_r4_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r4_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r4_p1_bits"};
      this.DqRxVrefDac_r4_p1.configure(this, null, "");
      this.DqRxVrefDac_r4_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r4_p1, `UVM_REG_ADDR_WIDTH'h4C8, "RW", 0);
		this.DqRxVrefDac_r4_p1_DqRxVrefDac_r4_p1 = this.DqRxVrefDac_r4_p1.DqRxVrefDac_r4_p1;
      this.RxClkT2UIDlyTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r5_p1::type_id::create("RxClkT2UIDlyTg0_r5_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r5_p1_bits"};
      this.RxClkT2UIDlyTg0_r5_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r5_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h510, "RW", 0);
		this.RxClkT2UIDlyTg0_r5_p1_RxClkT2UIDlyTg0_r5_p1 = this.RxClkT2UIDlyTg0_r5_p1.RxClkT2UIDlyTg0_r5_p1;
      this.RxClkT2UIDlyTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r5_p1::type_id::create("RxClkT2UIDlyTg1_r5_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r5_p1_bits"};
      this.RxClkT2UIDlyTg1_r5_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r5_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h511, "RW", 0);
		this.RxClkT2UIDlyTg1_r5_p1_RxClkT2UIDlyTg1_r5_p1 = this.RxClkT2UIDlyTg1_r5_p1.RxClkT2UIDlyTg1_r5_p1;
      this.RxClkC2UIDlyTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r5_p1::type_id::create("RxClkC2UIDlyTg0_r5_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r5_p1_bits"};
      this.RxClkC2UIDlyTg0_r5_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r5_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h512, "RW", 0);
		this.RxClkC2UIDlyTg0_r5_p1_RxClkC2UIDlyTg0_r5_p1 = this.RxClkC2UIDlyTg0_r5_p1.RxClkC2UIDlyTg0_r5_p1;
      this.RxClkC2UIDlyTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r5_p1::type_id::create("RxClkC2UIDlyTg1_r5_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r5_p1_bits"};
      this.RxClkC2UIDlyTg1_r5_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r5_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h513, "RW", 0);
		this.RxClkC2UIDlyTg1_r5_p1_RxClkC2UIDlyTg1_r5_p1 = this.RxClkC2UIDlyTg1_r5_p1.RxClkC2UIDlyTg1_r5_p1;
      this.TxDqLeftEyeOffsetTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r5_p1::type_id::create("TxDqLeftEyeOffsetTg0_r5_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r5_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r5_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r5_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h560, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r5_p1_TxDqLeftEyeOffsetTg0_r5_p1 = this.TxDqLeftEyeOffsetTg0_r5_p1.TxDqLeftEyeOffsetTg0_r5_p1;
      this.TxDqLeftEyeOffsetTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r5_p1::type_id::create("TxDqLeftEyeOffsetTg1_r5_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r5_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r5_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r5_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h561, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r5_p1_TxDqLeftEyeOffsetTg1_r5_p1 = this.TxDqLeftEyeOffsetTg1_r5_p1.TxDqLeftEyeOffsetTg1_r5_p1;
      this.TxDqRightEyeOffsetTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r5_p1::type_id::create("TxDqRightEyeOffsetTg0_r5_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r5_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r5_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r5_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h563, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r5_p1_TxDqRightEyeOffsetTg0_r5_p1 = this.TxDqRightEyeOffsetTg0_r5_p1.TxDqRightEyeOffsetTg0_r5_p1;
      this.TxDqRightEyeOffsetTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r5_p1::type_id::create("TxDqRightEyeOffsetTg1_r5_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r5_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r5_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r5_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h564, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r5_p1_TxDqRightEyeOffsetTg1_r5_p1 = this.TxDqRightEyeOffsetTg1_r5_p1.TxDqRightEyeOffsetTg1_r5_p1;
      this.RxClkTLeftEyeOffsetTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r5_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r5_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r5_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r5_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r5_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h568, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r5_p1_RxClkTLeftEyeOffsetTg0_r5_p1 = this.RxClkTLeftEyeOffsetTg0_r5_p1.RxClkTLeftEyeOffsetTg0_r5_p1;
      this.RxClkTLeftEyeOffsetTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r5_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r5_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r5_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r5_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r5_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h569, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r5_p1_RxClkTLeftEyeOffsetTg1_r5_p1 = this.RxClkTLeftEyeOffsetTg1_r5_p1.RxClkTLeftEyeOffsetTg1_r5_p1;
      this.RxClkTRightEyeOffsetTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r5_p1::type_id::create("RxClkTRightEyeOffsetTg0_r5_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r5_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r5_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r5_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h56A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r5_p1_RxClkTRightEyeOffsetTg0_r5_p1 = this.RxClkTRightEyeOffsetTg0_r5_p1.RxClkTRightEyeOffsetTg0_r5_p1;
      this.RxClkTRightEyeOffsetTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r5_p1::type_id::create("RxClkTRightEyeOffsetTg1_r5_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r5_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r5_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r5_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h56B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r5_p1_RxClkTRightEyeOffsetTg1_r5_p1 = this.RxClkTRightEyeOffsetTg1_r5_p1.RxClkTRightEyeOffsetTg1_r5_p1;
      this.RxClkCLeftEyeOffsetTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r5_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r5_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r5_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r5_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r5_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h56C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r5_p1_RxClkCLeftEyeOffsetTg0_r5_p1 = this.RxClkCLeftEyeOffsetTg0_r5_p1.RxClkCLeftEyeOffsetTg0_r5_p1;
      this.RxClkCLeftEyeOffsetTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r5_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r5_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r5_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r5_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r5_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h56D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r5_p1_RxClkCLeftEyeOffsetTg1_r5_p1 = this.RxClkCLeftEyeOffsetTg1_r5_p1.RxClkCLeftEyeOffsetTg1_r5_p1;
      this.RxClkCRightEyeOffsetTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r5_p1::type_id::create("RxClkCRightEyeOffsetTg0_r5_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r5_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r5_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r5_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h56E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r5_p1_RxClkCRightEyeOffsetTg0_r5_p1 = this.RxClkCRightEyeOffsetTg0_r5_p1.RxClkCRightEyeOffsetTg0_r5_p1;
      this.RxClkCRightEyeOffsetTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r5_p1::type_id::create("RxClkCRightEyeOffsetTg1_r5_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r5_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r5_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r5_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h56F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r5_p1_RxClkCRightEyeOffsetTg1_r5_p1 = this.RxClkCRightEyeOffsetTg1_r5_p1.RxClkCRightEyeOffsetTg1_r5_p1;
      this.RxDigStrbDlyTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r5_p1::type_id::create("RxDigStrbDlyTg0_r5_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r5_p1_bits"};
      this.RxDigStrbDlyTg0_r5_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r5_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h578, "RW", 0);
		this.RxDigStrbDlyTg0_r5_p1_RxDigStrbDlyTg0_r5_p1 = this.RxDigStrbDlyTg0_r5_p1.RxDigStrbDlyTg0_r5_p1;
      this.RxDigStrbDlyTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r5_p1::type_id::create("RxDigStrbDlyTg1_r5_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r5_p1_bits"};
      this.RxDigStrbDlyTg1_r5_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r5_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h579, "RW", 0);
		this.RxDigStrbDlyTg1_r5_p1_RxDigStrbDlyTg1_r5_p1 = this.RxDigStrbDlyTg1_r5_p1.RxDigStrbDlyTg1_r5_p1;
      this.TxDqDlyTg0_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r5_p1::type_id::create("TxDqDlyTg0_r5_p1",,get_full_name());
      if(this.TxDqDlyTg0_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r5_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r5_p1_bits"};
      this.TxDqDlyTg0_r5_p1.configure(this, null, "");
      this.TxDqDlyTg0_r5_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r5_p1, `UVM_REG_ADDR_WIDTH'h57A, "RW", 0);
		this.TxDqDlyTg0_r5_p1_TxDqDlyTg0_r5_p1 = this.TxDqDlyTg0_r5_p1.TxDqDlyTg0_r5_p1;
      this.TxDqDlyTg1_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r5_p1::type_id::create("TxDqDlyTg1_r5_p1",,get_full_name());
      if(this.TxDqDlyTg1_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r5_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r5_p1_bits"};
      this.TxDqDlyTg1_r5_p1.configure(this, null, "");
      this.TxDqDlyTg1_r5_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r5_p1, `UVM_REG_ADDR_WIDTH'h57B, "RW", 0);
		this.TxDqDlyTg1_r5_p1_TxDqDlyTg1_r5_p1 = this.TxDqDlyTg1_r5_p1.TxDqDlyTg1_r5_p1;
      this.DqRxVrefDac_r5_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r5_p1::type_id::create("DqRxVrefDac_r5_p1",,get_full_name());
      if(this.DqRxVrefDac_r5_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r5_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r5_p1_bits"};
      this.DqRxVrefDac_r5_p1.configure(this, null, "");
      this.DqRxVrefDac_r5_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r5_p1, `UVM_REG_ADDR_WIDTH'h5C8, "RW", 0);
		this.DqRxVrefDac_r5_p1_DqRxVrefDac_r5_p1 = this.DqRxVrefDac_r5_p1.DqRxVrefDac_r5_p1;
      this.RxClkT2UIDlyTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r6_p1::type_id::create("RxClkT2UIDlyTg0_r6_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r6_p1_bits"};
      this.RxClkT2UIDlyTg0_r6_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r6_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h610, "RW", 0);
		this.RxClkT2UIDlyTg0_r6_p1_RxClkT2UIDlyTg0_r6_p1 = this.RxClkT2UIDlyTg0_r6_p1.RxClkT2UIDlyTg0_r6_p1;
      this.RxClkT2UIDlyTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r6_p1::type_id::create("RxClkT2UIDlyTg1_r6_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r6_p1_bits"};
      this.RxClkT2UIDlyTg1_r6_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r6_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h611, "RW", 0);
		this.RxClkT2UIDlyTg1_r6_p1_RxClkT2UIDlyTg1_r6_p1 = this.RxClkT2UIDlyTg1_r6_p1.RxClkT2UIDlyTg1_r6_p1;
      this.RxClkC2UIDlyTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r6_p1::type_id::create("RxClkC2UIDlyTg0_r6_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r6_p1_bits"};
      this.RxClkC2UIDlyTg0_r6_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r6_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h612, "RW", 0);
		this.RxClkC2UIDlyTg0_r6_p1_RxClkC2UIDlyTg0_r6_p1 = this.RxClkC2UIDlyTg0_r6_p1.RxClkC2UIDlyTg0_r6_p1;
      this.RxClkC2UIDlyTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r6_p1::type_id::create("RxClkC2UIDlyTg1_r6_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r6_p1_bits"};
      this.RxClkC2UIDlyTg1_r6_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r6_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h613, "RW", 0);
		this.RxClkC2UIDlyTg1_r6_p1_RxClkC2UIDlyTg1_r6_p1 = this.RxClkC2UIDlyTg1_r6_p1.RxClkC2UIDlyTg1_r6_p1;
      this.TxDqLeftEyeOffsetTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r6_p1::type_id::create("TxDqLeftEyeOffsetTg0_r6_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r6_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r6_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r6_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h660, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r6_p1_TxDqLeftEyeOffsetTg0_r6_p1 = this.TxDqLeftEyeOffsetTg0_r6_p1.TxDqLeftEyeOffsetTg0_r6_p1;
      this.TxDqLeftEyeOffsetTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r6_p1::type_id::create("TxDqLeftEyeOffsetTg1_r6_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r6_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r6_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r6_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h661, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r6_p1_TxDqLeftEyeOffsetTg1_r6_p1 = this.TxDqLeftEyeOffsetTg1_r6_p1.TxDqLeftEyeOffsetTg1_r6_p1;
      this.TxDqRightEyeOffsetTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r6_p1::type_id::create("TxDqRightEyeOffsetTg0_r6_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r6_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r6_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r6_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h663, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r6_p1_TxDqRightEyeOffsetTg0_r6_p1 = this.TxDqRightEyeOffsetTg0_r6_p1.TxDqRightEyeOffsetTg0_r6_p1;
      this.TxDqRightEyeOffsetTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r6_p1::type_id::create("TxDqRightEyeOffsetTg1_r6_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r6_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r6_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r6_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h664, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r6_p1_TxDqRightEyeOffsetTg1_r6_p1 = this.TxDqRightEyeOffsetTg1_r6_p1.TxDqRightEyeOffsetTg1_r6_p1;
      this.RxClkTLeftEyeOffsetTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r6_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r6_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r6_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r6_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r6_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h668, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r6_p1_RxClkTLeftEyeOffsetTg0_r6_p1 = this.RxClkTLeftEyeOffsetTg0_r6_p1.RxClkTLeftEyeOffsetTg0_r6_p1;
      this.RxClkTLeftEyeOffsetTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r6_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r6_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r6_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r6_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r6_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h669, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r6_p1_RxClkTLeftEyeOffsetTg1_r6_p1 = this.RxClkTLeftEyeOffsetTg1_r6_p1.RxClkTLeftEyeOffsetTg1_r6_p1;
      this.RxClkTRightEyeOffsetTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r6_p1::type_id::create("RxClkTRightEyeOffsetTg0_r6_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r6_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r6_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r6_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h66A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r6_p1_RxClkTRightEyeOffsetTg0_r6_p1 = this.RxClkTRightEyeOffsetTg0_r6_p1.RxClkTRightEyeOffsetTg0_r6_p1;
      this.RxClkTRightEyeOffsetTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r6_p1::type_id::create("RxClkTRightEyeOffsetTg1_r6_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r6_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r6_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r6_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h66B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r6_p1_RxClkTRightEyeOffsetTg1_r6_p1 = this.RxClkTRightEyeOffsetTg1_r6_p1.RxClkTRightEyeOffsetTg1_r6_p1;
      this.RxClkCLeftEyeOffsetTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r6_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r6_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r6_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r6_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r6_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h66C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r6_p1_RxClkCLeftEyeOffsetTg0_r6_p1 = this.RxClkCLeftEyeOffsetTg0_r6_p1.RxClkCLeftEyeOffsetTg0_r6_p1;
      this.RxClkCLeftEyeOffsetTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r6_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r6_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r6_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r6_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r6_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h66D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r6_p1_RxClkCLeftEyeOffsetTg1_r6_p1 = this.RxClkCLeftEyeOffsetTg1_r6_p1.RxClkCLeftEyeOffsetTg1_r6_p1;
      this.RxClkCRightEyeOffsetTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r6_p1::type_id::create("RxClkCRightEyeOffsetTg0_r6_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r6_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r6_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r6_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h66E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r6_p1_RxClkCRightEyeOffsetTg0_r6_p1 = this.RxClkCRightEyeOffsetTg0_r6_p1.RxClkCRightEyeOffsetTg0_r6_p1;
      this.RxClkCRightEyeOffsetTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r6_p1::type_id::create("RxClkCRightEyeOffsetTg1_r6_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r6_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r6_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r6_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h66F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r6_p1_RxClkCRightEyeOffsetTg1_r6_p1 = this.RxClkCRightEyeOffsetTg1_r6_p1.RxClkCRightEyeOffsetTg1_r6_p1;
      this.RxDigStrbDlyTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r6_p1::type_id::create("RxDigStrbDlyTg0_r6_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r6_p1_bits"};
      this.RxDigStrbDlyTg0_r6_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r6_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h678, "RW", 0);
		this.RxDigStrbDlyTg0_r6_p1_RxDigStrbDlyTg0_r6_p1 = this.RxDigStrbDlyTg0_r6_p1.RxDigStrbDlyTg0_r6_p1;
      this.RxDigStrbDlyTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r6_p1::type_id::create("RxDigStrbDlyTg1_r6_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r6_p1_bits"};
      this.RxDigStrbDlyTg1_r6_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r6_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h679, "RW", 0);
		this.RxDigStrbDlyTg1_r6_p1_RxDigStrbDlyTg1_r6_p1 = this.RxDigStrbDlyTg1_r6_p1.RxDigStrbDlyTg1_r6_p1;
      this.TxDqDlyTg0_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r6_p1::type_id::create("TxDqDlyTg0_r6_p1",,get_full_name());
      if(this.TxDqDlyTg0_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r6_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r6_p1_bits"};
      this.TxDqDlyTg0_r6_p1.configure(this, null, "");
      this.TxDqDlyTg0_r6_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r6_p1, `UVM_REG_ADDR_WIDTH'h67A, "RW", 0);
		this.TxDqDlyTg0_r6_p1_TxDqDlyTg0_r6_p1 = this.TxDqDlyTg0_r6_p1.TxDqDlyTg0_r6_p1;
      this.TxDqDlyTg1_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r6_p1::type_id::create("TxDqDlyTg1_r6_p1",,get_full_name());
      if(this.TxDqDlyTg1_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r6_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r6_p1_bits"};
      this.TxDqDlyTg1_r6_p1.configure(this, null, "");
      this.TxDqDlyTg1_r6_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r6_p1, `UVM_REG_ADDR_WIDTH'h67B, "RW", 0);
		this.TxDqDlyTg1_r6_p1_TxDqDlyTg1_r6_p1 = this.TxDqDlyTg1_r6_p1.TxDqDlyTg1_r6_p1;
      this.DqRxVrefDac_r6_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r6_p1::type_id::create("DqRxVrefDac_r6_p1",,get_full_name());
      if(this.DqRxVrefDac_r6_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r6_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r6_p1_bits"};
      this.DqRxVrefDac_r6_p1.configure(this, null, "");
      this.DqRxVrefDac_r6_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r6_p1, `UVM_REG_ADDR_WIDTH'h6C8, "RW", 0);
		this.DqRxVrefDac_r6_p1_DqRxVrefDac_r6_p1 = this.DqRxVrefDac_r6_p1.DqRxVrefDac_r6_p1;
      this.RxClkT2UIDlyTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r7_p1::type_id::create("RxClkT2UIDlyTg0_r7_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r7_p1_bits"};
      this.RxClkT2UIDlyTg0_r7_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r7_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h710, "RW", 0);
		this.RxClkT2UIDlyTg0_r7_p1_RxClkT2UIDlyTg0_r7_p1 = this.RxClkT2UIDlyTg0_r7_p1.RxClkT2UIDlyTg0_r7_p1;
      this.RxClkT2UIDlyTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r7_p1::type_id::create("RxClkT2UIDlyTg1_r7_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r7_p1_bits"};
      this.RxClkT2UIDlyTg1_r7_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r7_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h711, "RW", 0);
		this.RxClkT2UIDlyTg1_r7_p1_RxClkT2UIDlyTg1_r7_p1 = this.RxClkT2UIDlyTg1_r7_p1.RxClkT2UIDlyTg1_r7_p1;
      this.RxClkC2UIDlyTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r7_p1::type_id::create("RxClkC2UIDlyTg0_r7_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r7_p1_bits"};
      this.RxClkC2UIDlyTg0_r7_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r7_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h712, "RW", 0);
		this.RxClkC2UIDlyTg0_r7_p1_RxClkC2UIDlyTg0_r7_p1 = this.RxClkC2UIDlyTg0_r7_p1.RxClkC2UIDlyTg0_r7_p1;
      this.RxClkC2UIDlyTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r7_p1::type_id::create("RxClkC2UIDlyTg1_r7_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r7_p1_bits"};
      this.RxClkC2UIDlyTg1_r7_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r7_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h713, "RW", 0);
		this.RxClkC2UIDlyTg1_r7_p1_RxClkC2UIDlyTg1_r7_p1 = this.RxClkC2UIDlyTg1_r7_p1.RxClkC2UIDlyTg1_r7_p1;
      this.TxDqLeftEyeOffsetTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r7_p1::type_id::create("TxDqLeftEyeOffsetTg0_r7_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r7_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r7_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r7_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h760, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r7_p1_TxDqLeftEyeOffsetTg0_r7_p1 = this.TxDqLeftEyeOffsetTg0_r7_p1.TxDqLeftEyeOffsetTg0_r7_p1;
      this.TxDqLeftEyeOffsetTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r7_p1::type_id::create("TxDqLeftEyeOffsetTg1_r7_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r7_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r7_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r7_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h761, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r7_p1_TxDqLeftEyeOffsetTg1_r7_p1 = this.TxDqLeftEyeOffsetTg1_r7_p1.TxDqLeftEyeOffsetTg1_r7_p1;
      this.TxDqRightEyeOffsetTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r7_p1::type_id::create("TxDqRightEyeOffsetTg0_r7_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r7_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r7_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r7_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h763, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r7_p1_TxDqRightEyeOffsetTg0_r7_p1 = this.TxDqRightEyeOffsetTg0_r7_p1.TxDqRightEyeOffsetTg0_r7_p1;
      this.TxDqRightEyeOffsetTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r7_p1::type_id::create("TxDqRightEyeOffsetTg1_r7_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r7_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r7_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r7_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h764, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r7_p1_TxDqRightEyeOffsetTg1_r7_p1 = this.TxDqRightEyeOffsetTg1_r7_p1.TxDqRightEyeOffsetTg1_r7_p1;
      this.RxClkTLeftEyeOffsetTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r7_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r7_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r7_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r7_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r7_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h768, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r7_p1_RxClkTLeftEyeOffsetTg0_r7_p1 = this.RxClkTLeftEyeOffsetTg0_r7_p1.RxClkTLeftEyeOffsetTg0_r7_p1;
      this.RxClkTLeftEyeOffsetTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r7_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r7_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r7_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r7_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r7_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h769, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r7_p1_RxClkTLeftEyeOffsetTg1_r7_p1 = this.RxClkTLeftEyeOffsetTg1_r7_p1.RxClkTLeftEyeOffsetTg1_r7_p1;
      this.RxClkTRightEyeOffsetTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r7_p1::type_id::create("RxClkTRightEyeOffsetTg0_r7_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r7_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r7_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r7_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h76A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r7_p1_RxClkTRightEyeOffsetTg0_r7_p1 = this.RxClkTRightEyeOffsetTg0_r7_p1.RxClkTRightEyeOffsetTg0_r7_p1;
      this.RxClkTRightEyeOffsetTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r7_p1::type_id::create("RxClkTRightEyeOffsetTg1_r7_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r7_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r7_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r7_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h76B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r7_p1_RxClkTRightEyeOffsetTg1_r7_p1 = this.RxClkTRightEyeOffsetTg1_r7_p1.RxClkTRightEyeOffsetTg1_r7_p1;
      this.RxClkCLeftEyeOffsetTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r7_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r7_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r7_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r7_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r7_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h76C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r7_p1_RxClkCLeftEyeOffsetTg0_r7_p1 = this.RxClkCLeftEyeOffsetTg0_r7_p1.RxClkCLeftEyeOffsetTg0_r7_p1;
      this.RxClkCLeftEyeOffsetTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r7_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r7_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r7_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r7_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r7_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h76D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r7_p1_RxClkCLeftEyeOffsetTg1_r7_p1 = this.RxClkCLeftEyeOffsetTg1_r7_p1.RxClkCLeftEyeOffsetTg1_r7_p1;
      this.RxClkCRightEyeOffsetTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r7_p1::type_id::create("RxClkCRightEyeOffsetTg0_r7_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r7_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r7_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r7_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h76E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r7_p1_RxClkCRightEyeOffsetTg0_r7_p1 = this.RxClkCRightEyeOffsetTg0_r7_p1.RxClkCRightEyeOffsetTg0_r7_p1;
      this.RxClkCRightEyeOffsetTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r7_p1::type_id::create("RxClkCRightEyeOffsetTg1_r7_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r7_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r7_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r7_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h76F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r7_p1_RxClkCRightEyeOffsetTg1_r7_p1 = this.RxClkCRightEyeOffsetTg1_r7_p1.RxClkCRightEyeOffsetTg1_r7_p1;
      this.RxDigStrbDlyTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r7_p1::type_id::create("RxDigStrbDlyTg0_r7_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r7_p1_bits"};
      this.RxDigStrbDlyTg0_r7_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r7_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h778, "RW", 0);
		this.RxDigStrbDlyTg0_r7_p1_RxDigStrbDlyTg0_r7_p1 = this.RxDigStrbDlyTg0_r7_p1.RxDigStrbDlyTg0_r7_p1;
      this.RxDigStrbDlyTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r7_p1::type_id::create("RxDigStrbDlyTg1_r7_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r7_p1_bits"};
      this.RxDigStrbDlyTg1_r7_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r7_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h779, "RW", 0);
		this.RxDigStrbDlyTg1_r7_p1_RxDigStrbDlyTg1_r7_p1 = this.RxDigStrbDlyTg1_r7_p1.RxDigStrbDlyTg1_r7_p1;
      this.TxDqDlyTg0_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r7_p1::type_id::create("TxDqDlyTg0_r7_p1",,get_full_name());
      if(this.TxDqDlyTg0_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r7_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r7_p1_bits"};
      this.TxDqDlyTg0_r7_p1.configure(this, null, "");
      this.TxDqDlyTg0_r7_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r7_p1, `UVM_REG_ADDR_WIDTH'h77A, "RW", 0);
		this.TxDqDlyTg0_r7_p1_TxDqDlyTg0_r7_p1 = this.TxDqDlyTg0_r7_p1.TxDqDlyTg0_r7_p1;
      this.TxDqDlyTg1_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r7_p1::type_id::create("TxDqDlyTg1_r7_p1",,get_full_name());
      if(this.TxDqDlyTg1_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r7_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r7_p1_bits"};
      this.TxDqDlyTg1_r7_p1.configure(this, null, "");
      this.TxDqDlyTg1_r7_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r7_p1, `UVM_REG_ADDR_WIDTH'h77B, "RW", 0);
		this.TxDqDlyTg1_r7_p1_TxDqDlyTg1_r7_p1 = this.TxDqDlyTg1_r7_p1.TxDqDlyTg1_r7_p1;
      this.DqRxVrefDac_r7_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r7_p1::type_id::create("DqRxVrefDac_r7_p1",,get_full_name());
      if(this.DqRxVrefDac_r7_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r7_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r7_p1_bits"};
      this.DqRxVrefDac_r7_p1.configure(this, null, "");
      this.DqRxVrefDac_r7_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r7_p1, `UVM_REG_ADDR_WIDTH'h7C8, "RW", 0);
		this.DqRxVrefDac_r7_p1_DqRxVrefDac_r7_p1 = this.DqRxVrefDac_r7_p1.DqRxVrefDac_r7_p1;
      this.PclkDCAStaticCtrl0DB_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl0DB_p1::type_id::create("PclkDCAStaticCtrl0DB_p1",,get_full_name());
      if(this.PclkDCAStaticCtrl0DB_p1.has_coverage(UVM_CVR_ALL))
      	this.PclkDCAStaticCtrl0DB_p1.cg_bits.option.name = {get_name(), ".", "PclkDCAStaticCtrl0DB_p1_bits"};
      this.PclkDCAStaticCtrl0DB_p1.configure(this, null, "");
      this.PclkDCAStaticCtrl0DB_p1.build();
      this.default_map.add_reg(this.PclkDCAStaticCtrl0DB_p1, `UVM_REG_ADDR_WIDTH'h803, "RW", 0);
		this.PclkDCAStaticCtrl0DB_p1_PclkDCACalModeDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCACalModeDB;
		this.PclkDCACalModeDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCACalModeDB;
		this.PclkDCAStaticCtrl0DB_p1_PclkDCAEnDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCAEnDB;
		this.PclkDCAEnDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCAEnDB;
		this.PclkDCAStaticCtrl0DB_p1_PclkDCATxLcdlPhSelDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCATxLcdlPhSelDB;
		this.PclkDCATxLcdlPhSelDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCATxLcdlPhSelDB;
		this.PclkDCAStaticCtrl0DB_p1_PclkDCDSettleDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCDSettleDB;
		this.PclkDCDSettleDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCDSettleDB;
		this.PclkDCAStaticCtrl0DB_p1_PclkDCDSampTimeDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCDSampTimeDB;
		this.PclkDCDSampTimeDB = this.PclkDCAStaticCtrl0DB_p1.PclkDCDSampTimeDB;
      this.PclkDCASampDelayLCDLDB_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCASampDelayLCDLDB_p1::type_id::create("PclkDCASampDelayLCDLDB_p1",,get_full_name());
      if(this.PclkDCASampDelayLCDLDB_p1.has_coverage(UVM_CVR_ALL))
      	this.PclkDCASampDelayLCDLDB_p1.cg_bits.option.name = {get_name(), ".", "PclkDCASampDelayLCDLDB_p1_bits"};
      this.PclkDCASampDelayLCDLDB_p1.configure(this, null, "");
      this.PclkDCASampDelayLCDLDB_p1.build();
      this.default_map.add_reg(this.PclkDCASampDelayLCDLDB_p1, `UVM_REG_ADDR_WIDTH'h80B, "RW", 0);
		this.PclkDCASampDelayLCDLDB_p1_PclkDCASampDelayLCDLDB_p1 = this.PclkDCASampDelayLCDLDB_p1.PclkDCASampDelayLCDLDB_p1;
      this.RxClkT2UIDlyTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg0_r8_p1::type_id::create("RxClkT2UIDlyTg0_r8_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg0_r8_p1_bits"};
      this.RxClkT2UIDlyTg0_r8_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg0_r8_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h810, "RW", 0);
		this.RxClkT2UIDlyTg0_r8_p1_RxClkT2UIDlyTg0_r8_p1 = this.RxClkT2UIDlyTg0_r8_p1.RxClkT2UIDlyTg0_r8_p1;
      this.RxClkT2UIDlyTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkT2UIDlyTg1_r8_p1::type_id::create("RxClkT2UIDlyTg1_r8_p1",,get_full_name());
      if(this.RxClkT2UIDlyTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkT2UIDlyTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkT2UIDlyTg1_r8_p1_bits"};
      this.RxClkT2UIDlyTg1_r8_p1.configure(this, null, "");
      this.RxClkT2UIDlyTg1_r8_p1.build();
      this.default_map.add_reg(this.RxClkT2UIDlyTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h811, "RW", 0);
		this.RxClkT2UIDlyTg1_r8_p1_RxClkT2UIDlyTg1_r8_p1 = this.RxClkT2UIDlyTg1_r8_p1.RxClkT2UIDlyTg1_r8_p1;
      this.RxClkC2UIDlyTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg0_r8_p1::type_id::create("RxClkC2UIDlyTg0_r8_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg0_r8_p1_bits"};
      this.RxClkC2UIDlyTg0_r8_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg0_r8_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h812, "RW", 0);
		this.RxClkC2UIDlyTg0_r8_p1_RxClkC2UIDlyTg0_r8_p1 = this.RxClkC2UIDlyTg0_r8_p1.RxClkC2UIDlyTg0_r8_p1;
      this.RxClkC2UIDlyTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkC2UIDlyTg1_r8_p1::type_id::create("RxClkC2UIDlyTg1_r8_p1",,get_full_name());
      if(this.RxClkC2UIDlyTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkC2UIDlyTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkC2UIDlyTg1_r8_p1_bits"};
      this.RxClkC2UIDlyTg1_r8_p1.configure(this, null, "");
      this.RxClkC2UIDlyTg1_r8_p1.build();
      this.default_map.add_reg(this.RxClkC2UIDlyTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h813, "RW", 0);
		this.RxClkC2UIDlyTg1_r8_p1_RxClkC2UIDlyTg1_r8_p1 = this.RxClkC2UIDlyTg1_r8_p1.RxClkC2UIDlyTg1_r8_p1;
      this.TxDqLeftEyeOffsetTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg0_r8_p1::type_id::create("TxDqLeftEyeOffsetTg0_r8_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg0_r8_p1_bits"};
      this.TxDqLeftEyeOffsetTg0_r8_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg0_r8_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h860, "RW", 0);
		this.TxDqLeftEyeOffsetTg0_r8_p1_TxDqLeftEyeOffsetTg0_r8_p1 = this.TxDqLeftEyeOffsetTg0_r8_p1.TxDqLeftEyeOffsetTg0_r8_p1;
      this.TxDqLeftEyeOffsetTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqLeftEyeOffsetTg1_r8_p1::type_id::create("TxDqLeftEyeOffsetTg1_r8_p1",,get_full_name());
      if(this.TxDqLeftEyeOffsetTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqLeftEyeOffsetTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "TxDqLeftEyeOffsetTg1_r8_p1_bits"};
      this.TxDqLeftEyeOffsetTg1_r8_p1.configure(this, null, "");
      this.TxDqLeftEyeOffsetTg1_r8_p1.build();
      this.default_map.add_reg(this.TxDqLeftEyeOffsetTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h861, "RW", 0);
		this.TxDqLeftEyeOffsetTg1_r8_p1_TxDqLeftEyeOffsetTg1_r8_p1 = this.TxDqLeftEyeOffsetTg1_r8_p1.TxDqLeftEyeOffsetTg1_r8_p1;
      this.TxDqRightEyeOffsetTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg0_r8_p1::type_id::create("TxDqRightEyeOffsetTg0_r8_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg0_r8_p1_bits"};
      this.TxDqRightEyeOffsetTg0_r8_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg0_r8_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h863, "RW", 0);
		this.TxDqRightEyeOffsetTg0_r8_p1_TxDqRightEyeOffsetTg0_r8_p1 = this.TxDqRightEyeOffsetTg0_r8_p1.TxDqRightEyeOffsetTg0_r8_p1;
      this.TxDqRightEyeOffsetTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqRightEyeOffsetTg1_r8_p1::type_id::create("TxDqRightEyeOffsetTg1_r8_p1",,get_full_name());
      if(this.TxDqRightEyeOffsetTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqRightEyeOffsetTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "TxDqRightEyeOffsetTg1_r8_p1_bits"};
      this.TxDqRightEyeOffsetTg1_r8_p1.configure(this, null, "");
      this.TxDqRightEyeOffsetTg1_r8_p1.build();
      this.default_map.add_reg(this.TxDqRightEyeOffsetTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h864, "RW", 0);
		this.TxDqRightEyeOffsetTg1_r8_p1_TxDqRightEyeOffsetTg1_r8_p1 = this.TxDqRightEyeOffsetTg1_r8_p1.TxDqRightEyeOffsetTg1_r8_p1;
      this.RxClkTLeftEyeOffsetTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg0_r8_p1::type_id::create("RxClkTLeftEyeOffsetTg0_r8_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg0_r8_p1_bits"};
      this.RxClkTLeftEyeOffsetTg0_r8_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg0_r8_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h868, "RW", 0);
		this.RxClkTLeftEyeOffsetTg0_r8_p1_RxClkTLeftEyeOffsetTg0_r8_p1 = this.RxClkTLeftEyeOffsetTg0_r8_p1.RxClkTLeftEyeOffsetTg0_r8_p1;
      this.RxClkTLeftEyeOffsetTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTLeftEyeOffsetTg1_r8_p1::type_id::create("RxClkTLeftEyeOffsetTg1_r8_p1",,get_full_name());
      if(this.RxClkTLeftEyeOffsetTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTLeftEyeOffsetTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkTLeftEyeOffsetTg1_r8_p1_bits"};
      this.RxClkTLeftEyeOffsetTg1_r8_p1.configure(this, null, "");
      this.RxClkTLeftEyeOffsetTg1_r8_p1.build();
      this.default_map.add_reg(this.RxClkTLeftEyeOffsetTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h869, "RW", 0);
		this.RxClkTLeftEyeOffsetTg1_r8_p1_RxClkTLeftEyeOffsetTg1_r8_p1 = this.RxClkTLeftEyeOffsetTg1_r8_p1.RxClkTLeftEyeOffsetTg1_r8_p1;
      this.RxClkTRightEyeOffsetTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg0_r8_p1::type_id::create("RxClkTRightEyeOffsetTg0_r8_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg0_r8_p1_bits"};
      this.RxClkTRightEyeOffsetTg0_r8_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg0_r8_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h86A, "RW", 0);
		this.RxClkTRightEyeOffsetTg0_r8_p1_RxClkTRightEyeOffsetTg0_r8_p1 = this.RxClkTRightEyeOffsetTg0_r8_p1.RxClkTRightEyeOffsetTg0_r8_p1;
      this.RxClkTRightEyeOffsetTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkTRightEyeOffsetTg1_r8_p1::type_id::create("RxClkTRightEyeOffsetTg1_r8_p1",,get_full_name());
      if(this.RxClkTRightEyeOffsetTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkTRightEyeOffsetTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkTRightEyeOffsetTg1_r8_p1_bits"};
      this.RxClkTRightEyeOffsetTg1_r8_p1.configure(this, null, "");
      this.RxClkTRightEyeOffsetTg1_r8_p1.build();
      this.default_map.add_reg(this.RxClkTRightEyeOffsetTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h86B, "RW", 0);
		this.RxClkTRightEyeOffsetTg1_r8_p1_RxClkTRightEyeOffsetTg1_r8_p1 = this.RxClkTRightEyeOffsetTg1_r8_p1.RxClkTRightEyeOffsetTg1_r8_p1;
      this.RxClkCLeftEyeOffsetTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg0_r8_p1::type_id::create("RxClkCLeftEyeOffsetTg0_r8_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg0_r8_p1_bits"};
      this.RxClkCLeftEyeOffsetTg0_r8_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg0_r8_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h86C, "RW", 0);
		this.RxClkCLeftEyeOffsetTg0_r8_p1_RxClkCLeftEyeOffsetTg0_r8_p1 = this.RxClkCLeftEyeOffsetTg0_r8_p1.RxClkCLeftEyeOffsetTg0_r8_p1;
      this.RxClkCLeftEyeOffsetTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCLeftEyeOffsetTg1_r8_p1::type_id::create("RxClkCLeftEyeOffsetTg1_r8_p1",,get_full_name());
      if(this.RxClkCLeftEyeOffsetTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCLeftEyeOffsetTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkCLeftEyeOffsetTg1_r8_p1_bits"};
      this.RxClkCLeftEyeOffsetTg1_r8_p1.configure(this, null, "");
      this.RxClkCLeftEyeOffsetTg1_r8_p1.build();
      this.default_map.add_reg(this.RxClkCLeftEyeOffsetTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h86D, "RW", 0);
		this.RxClkCLeftEyeOffsetTg1_r8_p1_RxClkCLeftEyeOffsetTg1_r8_p1 = this.RxClkCLeftEyeOffsetTg1_r8_p1.RxClkCLeftEyeOffsetTg1_r8_p1;
      this.RxClkCRightEyeOffsetTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg0_r8_p1::type_id::create("RxClkCRightEyeOffsetTg0_r8_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg0_r8_p1_bits"};
      this.RxClkCRightEyeOffsetTg0_r8_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg0_r8_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h86E, "RW", 0);
		this.RxClkCRightEyeOffsetTg0_r8_p1_RxClkCRightEyeOffsetTg0_r8_p1 = this.RxClkCRightEyeOffsetTg0_r8_p1.RxClkCRightEyeOffsetTg0_r8_p1;
      this.RxClkCRightEyeOffsetTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxClkCRightEyeOffsetTg1_r8_p1::type_id::create("RxClkCRightEyeOffsetTg1_r8_p1",,get_full_name());
      if(this.RxClkCRightEyeOffsetTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxClkCRightEyeOffsetTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "RxClkCRightEyeOffsetTg1_r8_p1_bits"};
      this.RxClkCRightEyeOffsetTg1_r8_p1.configure(this, null, "");
      this.RxClkCRightEyeOffsetTg1_r8_p1.build();
      this.default_map.add_reg(this.RxClkCRightEyeOffsetTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h86F, "RW", 0);
		this.RxClkCRightEyeOffsetTg1_r8_p1_RxClkCRightEyeOffsetTg1_r8_p1 = this.RxClkCRightEyeOffsetTg1_r8_p1.RxClkCRightEyeOffsetTg1_r8_p1;
      this.RxDigStrbDlyTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg0_r8_p1::type_id::create("RxDigStrbDlyTg0_r8_p1",,get_full_name());
      if(this.RxDigStrbDlyTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg0_r8_p1_bits"};
      this.RxDigStrbDlyTg0_r8_p1.configure(this, null, "");
      this.RxDigStrbDlyTg0_r8_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h878, "RW", 0);
		this.RxDigStrbDlyTg0_r8_p1_RxDigStrbDlyTg0_r8_p1 = this.RxDigStrbDlyTg0_r8_p1.RxDigStrbDlyTg0_r8_p1;
      this.RxDigStrbDlyTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_RxDigStrbDlyTg1_r8_p1::type_id::create("RxDigStrbDlyTg1_r8_p1",,get_full_name());
      if(this.RxDigStrbDlyTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.RxDigStrbDlyTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "RxDigStrbDlyTg1_r8_p1_bits"};
      this.RxDigStrbDlyTg1_r8_p1.configure(this, null, "");
      this.RxDigStrbDlyTg1_r8_p1.build();
      this.default_map.add_reg(this.RxDigStrbDlyTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h879, "RW", 0);
		this.RxDigStrbDlyTg1_r8_p1_RxDigStrbDlyTg1_r8_p1 = this.RxDigStrbDlyTg1_r8_p1.RxDigStrbDlyTg1_r8_p1;
      this.TxDqDlyTg0_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg0_r8_p1::type_id::create("TxDqDlyTg0_r8_p1",,get_full_name());
      if(this.TxDqDlyTg0_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg0_r8_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg0_r8_p1_bits"};
      this.TxDqDlyTg0_r8_p1.configure(this, null, "");
      this.TxDqDlyTg0_r8_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg0_r8_p1, `UVM_REG_ADDR_WIDTH'h87A, "RW", 0);
		this.TxDqDlyTg0_r8_p1_TxDqDlyTg0_r8_p1 = this.TxDqDlyTg0_r8_p1.TxDqDlyTg0_r8_p1;
      this.TxDqDlyTg1_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_TxDqDlyTg1_r8_p1::type_id::create("TxDqDlyTg1_r8_p1",,get_full_name());
      if(this.TxDqDlyTg1_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.TxDqDlyTg1_r8_p1.cg_bits.option.name = {get_name(), ".", "TxDqDlyTg1_r8_p1_bits"};
      this.TxDqDlyTg1_r8_p1.configure(this, null, "");
      this.TxDqDlyTg1_r8_p1.build();
      this.default_map.add_reg(this.TxDqDlyTg1_r8_p1, `UVM_REG_ADDR_WIDTH'h87B, "RW", 0);
		this.TxDqDlyTg1_r8_p1_TxDqDlyTg1_r8_p1 = this.TxDqDlyTg1_r8_p1.TxDqDlyTg1_r8_p1;
      this.DqRxVrefDac_r8_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_DqRxVrefDac_r8_p1::type_id::create("DqRxVrefDac_r8_p1",,get_full_name());
      if(this.DqRxVrefDac_r8_p1.has_coverage(UVM_CVR_ALL))
      	this.DqRxVrefDac_r8_p1.cg_bits.option.name = {get_name(), ".", "DqRxVrefDac_r8_p1_bits"};
      this.DqRxVrefDac_r8_p1.configure(this, null, "");
      this.DqRxVrefDac_r8_p1.build();
      this.default_map.add_reg(this.DqRxVrefDac_r8_p1, `UVM_REG_ADDR_WIDTH'h8C8, "RW", 0);
		this.DqRxVrefDac_r8_p1_DqRxVrefDac_r8_p1 = this.DqRxVrefDac_r8_p1.DqRxVrefDac_r8_p1;
      this.PclkDCAStaticCtrl1DB_p1 = ral_reg_DWC_DDRPHYA_DBYTE3_p1_PclkDCAStaticCtrl1DB_p1::type_id::create("PclkDCAStaticCtrl1DB_p1",,get_full_name());
      if(this.PclkDCAStaticCtrl1DB_p1.has_coverage(UVM_CVR_ALL))
      	this.PclkDCAStaticCtrl1DB_p1.cg_bits.option.name = {get_name(), ".", "PclkDCAStaticCtrl1DB_p1_bits"};
      this.PclkDCAStaticCtrl1DB_p1.configure(this, null, "");
      this.PclkDCAStaticCtrl1DB_p1.build();
      this.default_map.add_reg(this.PclkDCAStaticCtrl1DB_p1, `UVM_REG_ADDR_WIDTH'hC03, "RW", 0);
		this.PclkDCAStaticCtrl1DB_p1_PclkDCAInvertSampDB = this.PclkDCAStaticCtrl1DB_p1.PclkDCAInvertSampDB;
		this.PclkDCAInvertSampDB = this.PclkDCAStaticCtrl1DB_p1.PclkDCAInvertSampDB;
		this.PclkDCAStaticCtrl1DB_p1_PclkDCALcdlEn4pDB = this.PclkDCAStaticCtrl1DB_p1.PclkDCALcdlEn4pDB;
		this.PclkDCALcdlEn4pDB = this.PclkDCAStaticCtrl1DB_p1.PclkDCALcdlEn4pDB;
		this.PclkDCAStaticCtrl1DB_p1_PclkDCDMissionModeDelayDB = this.PclkDCAStaticCtrl1DB_p1.PclkDCDMissionModeDelayDB;
		this.PclkDCDMissionModeDelayDB = this.PclkDCAStaticCtrl1DB_p1.PclkDCDMissionModeDelayDB;
   endfunction : build

	`uvm_object_utils(ral_block_DWC_DDRPHYA_DBYTE3_p1)


function void sample(uvm_reg_addr_t offset,
                     bit            is_read,
                     uvm_reg_map    map);
  if (get_coverage(UVM_CVR_ADDR_MAP)) begin
    m_offset = offset;
    cg_addr.sample();
  end
endfunction
endclass : ral_block_DWC_DDRPHYA_DBYTE3_p1


endpackage
`endif
