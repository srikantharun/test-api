// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_soc
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_soc (
    input  wire                                     i_apu_aon_clk,
    input  wire                                     i_apu_aon_rst_n,
    input  chip_pkg::chip_axi_addr_t                i_apu_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_apu_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_apu_init_lt_axi_s_arcache,
    input  logic[9:0]                               i_apu_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_apu_init_lt_axi_s_arlen,
    input  logic                                    i_apu_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_apu_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_apu_init_lt_axi_s_arqos,
    output logic                                    o_apu_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_apu_init_lt_axi_s_arsize,
    input  logic                                    i_apu_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                i_apu_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_apu_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_apu_init_lt_axi_s_awcache,
    input  logic[9:0]                               i_apu_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_apu_init_lt_axi_s_awlen,
    input  logic                                    i_apu_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_apu_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_apu_init_lt_axi_s_awqos,
    output logic                                    o_apu_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_apu_init_lt_axi_s_awsize,
    input  logic                                    i_apu_init_lt_axi_s_awvalid,
    output logic[9:0]                               o_apu_init_lt_axi_s_bid,
    input  logic                                    i_apu_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_apu_init_lt_axi_s_bresp,
    output logic                                    o_apu_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t             o_apu_init_lt_axi_s_rdata,
    output logic[9:0]                               o_apu_init_lt_axi_s_rid,
    output logic                                    o_apu_init_lt_axi_s_rlast,
    input  logic                                    i_apu_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_apu_init_lt_axi_s_rresp,
    output logic                                    o_apu_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_apu_init_lt_axi_s_wdata,
    input  logic                                    i_apu_init_lt_axi_s_wlast,
    output logic                                    o_apu_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t            i_apu_init_lt_axi_s_wstrb,
    input  logic                                    i_apu_init_lt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_apu_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_apu_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_apu_init_mt_axi_s_arcache,
    input  logic[8:0]                               i_apu_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_apu_init_mt_axi_s_arlen,
    input  logic                                    i_apu_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_apu_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_apu_init_mt_axi_s_arqos,
    output logic                                    o_apu_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_apu_init_mt_axi_s_arsize,
    input  logic                                    i_apu_init_mt_axi_s_arvalid,
    output apu_pkg::apu_axi_mt_data_t               o_apu_init_mt_axi_s_rdata,
    output logic[8:0]                               o_apu_init_mt_axi_s_rid,
    output logic                                    o_apu_init_mt_axi_s_rlast,
    input  logic                                    i_apu_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_apu_init_mt_axi_s_rresp,
    output logic                                    o_apu_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_apu_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_apu_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_apu_init_mt_axi_s_awcache,
    input  logic[8:0]                               i_apu_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_apu_init_mt_axi_s_awlen,
    input  logic                                    i_apu_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_apu_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_apu_init_mt_axi_s_awqos,
    output logic                                    o_apu_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_apu_init_mt_axi_s_awsize,
    input  logic                                    i_apu_init_mt_axi_s_awvalid,
    output logic[8:0]                               o_apu_init_mt_axi_s_bid,
    input  logic                                    i_apu_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_apu_init_mt_axi_s_bresp,
    output logic                                    o_apu_init_mt_axi_s_bvalid,
    input  apu_pkg::apu_axi_mt_data_t               i_apu_init_mt_axi_s_wdata,
    input  logic                                    i_apu_init_mt_axi_s_wlast,
    output logic                                    o_apu_init_mt_axi_s_wready,
    input  apu_pkg::apu_axi_mt_wstrb_t              i_apu_init_mt_axi_s_wstrb,
    input  logic                                    i_apu_init_mt_axi_s_wvalid,
    output logic                                    o_apu_pwr_idle_val,
    output logic                                    o_apu_pwr_idle_ack,
    input  logic                                    i_apu_pwr_idle_req,
    output chip_pkg::chip_axi_addr_t                o_apu_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_apu_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_apu_targ_lt_axi_m_arcache,
    output logic[7:0]                               o_apu_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_apu_targ_lt_axi_m_arlen,
    output logic                                    o_apu_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_apu_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_apu_targ_lt_axi_m_arqos,
    input  logic                                    i_apu_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_apu_targ_lt_axi_m_arsize,
    output logic                                    o_apu_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_apu_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_apu_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_apu_targ_lt_axi_m_awcache,
    output logic[7:0]                               o_apu_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_apu_targ_lt_axi_m_awlen,
    output logic                                    o_apu_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_apu_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_apu_targ_lt_axi_m_awqos,
    input  logic                                    i_apu_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_apu_targ_lt_axi_m_awsize,
    output logic                                    o_apu_targ_lt_axi_m_awvalid,
    input  logic[7:0]                               i_apu_targ_lt_axi_m_bid,
    output logic                                    o_apu_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_apu_targ_lt_axi_m_bresp,
    input  logic                                    i_apu_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_apu_targ_lt_axi_m_rdata,
    input  logic[7:0]                               i_apu_targ_lt_axi_m_rid,
    input  logic                                    i_apu_targ_lt_axi_m_rlast,
    output logic                                    o_apu_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_apu_targ_lt_axi_m_rresp,
    input  logic                                    i_apu_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_apu_targ_lt_axi_m_wdata,
    output logic                                    o_apu_targ_lt_axi_m_wlast,
    input  logic                                    i_apu_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_apu_targ_lt_axi_m_wstrb,
    output logic                                    o_apu_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_apu_targ_syscfg_apb_m_paddr,
    output logic                                    o_apu_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_apu_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_apu_targ_syscfg_apb_m_prdata,
    input  logic                                    i_apu_targ_syscfg_apb_m_pready,
    output logic                                    o_apu_targ_syscfg_apb_m_psel,
    input  logic                                    i_apu_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_apu_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_apu_targ_syscfg_apb_m_pwdata,
    output logic                                    o_apu_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_apu_x_clk,
    input  wire                                     i_apu_x_clken,
    input  wire                                     i_apu_x_rst_n,
    input  wire                                     i_dcd_aon_clk,
    input  wire                                     i_dcd_aon_rst_n,
    input  wire                                     i_dcd_codec_clk,
    input  wire                                     i_dcd_codec_clken,
    input  wire                                     i_dcd_codec_rst_n,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_0_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_0_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_0_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_0_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_0_init_mt_axi_s_arlen,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_0_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_0_init_mt_axi_s_arqos,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_0_init_mt_axi_s_arsize,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_arvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_data_t    o_dcd_dec_0_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_0_init_mt_axi_s_rid,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_rlast,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_0_init_mt_axi_s_rresp,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_0_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_0_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_0_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_0_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_0_init_mt_axi_s_awlen,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_0_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_0_init_mt_axi_s_awqos,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_0_init_mt_axi_s_awsize,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_0_init_mt_axi_s_bid,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_0_init_mt_axi_s_bresp,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_bvalid,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_data_t    i_dcd_dec_0_init_mt_axi_s_wdata,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_wlast,
    output logic                                    o_dcd_dec_0_init_mt_axi_s_wready,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_strb_t    i_dcd_dec_0_init_mt_axi_s_wstrb,
    input  logic                                    i_dcd_dec_0_init_mt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_1_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_1_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_1_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_1_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_1_init_mt_axi_s_arlen,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_1_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_1_init_mt_axi_s_arqos,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_1_init_mt_axi_s_arsize,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_arvalid,
    output dcd_pkg::dcd_dec_1_init_mt_axi_data_t    o_dcd_dec_1_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_1_init_mt_axi_s_rid,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_rlast,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_1_init_mt_axi_s_rresp,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_1_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_1_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_1_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_1_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_1_init_mt_axi_s_awlen,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_1_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_1_init_mt_axi_s_awqos,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_1_init_mt_axi_s_awsize,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_1_init_mt_axi_s_bid,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_1_init_mt_axi_s_bresp,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_bvalid,
    input  dcd_pkg::dcd_dec_1_init_mt_axi_data_t    i_dcd_dec_1_init_mt_axi_s_wdata,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_wlast,
    output logic                                    o_dcd_dec_1_init_mt_axi_s_wready,
    input  dcd_pkg::dcd_dec_1_init_mt_axi_strb_t    i_dcd_dec_1_init_mt_axi_s_wstrb,
    input  logic                                    i_dcd_dec_1_init_mt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_2_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_2_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_2_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_2_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_2_init_mt_axi_s_arlen,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_2_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_2_init_mt_axi_s_arqos,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_2_init_mt_axi_s_arsize,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_arvalid,
    output logic [127:0]                            o_dcd_dec_2_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_2_init_mt_axi_s_rid,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_rlast,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_2_init_mt_axi_s_rresp,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_dec_2_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_dcd_dec_2_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_dcd_dec_2_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t      i_dcd_dec_2_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_dcd_dec_2_init_mt_axi_s_awlen,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_dcd_dec_2_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_dcd_dec_2_init_mt_axi_s_awqos,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_dcd_dec_2_init_mt_axi_s_awsize,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t      o_dcd_dec_2_init_mt_axi_s_bid,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_dcd_dec_2_init_mt_axi_s_bresp,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_bvalid,
    input  logic [127:0]                            i_dcd_dec_2_init_mt_axi_s_wdata,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_wlast,
    output logic                                    o_dcd_dec_2_init_mt_axi_s_wready,
    input  logic [15:0]                             i_dcd_dec_2_init_mt_axi_s_wstrb,
    input  logic                                    i_dcd_dec_2_init_mt_axi_s_wvalid,
    input  wire                                     i_dcd_mcu_clk,
    input  wire                                     i_dcd_mcu_clken,
    input  chip_pkg::chip_axi_addr_t                i_dcd_mcu_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_dcd_mcu_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_dcd_mcu_init_lt_axi_s_arcache,
    input  dcd_pkg::dcd_mcu_init_lt_axi_id_t        i_dcd_mcu_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_dcd_mcu_init_lt_axi_s_arlen,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_dcd_mcu_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_dcd_mcu_init_lt_axi_s_arqos,
    output logic                                    o_dcd_mcu_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_dcd_mcu_init_lt_axi_s_arsize,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_arvalid,
    output dcd_pkg::dcd_mcu_init_lt_axi_data_t      o_dcd_mcu_init_lt_axi_s_rdata,
    output dcd_pkg::dcd_mcu_init_lt_axi_id_t        o_dcd_mcu_init_lt_axi_s_rid,
    output logic                                    o_dcd_mcu_init_lt_axi_s_rlast,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_dcd_mcu_init_lt_axi_s_rresp,
    output logic                                    o_dcd_mcu_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_dcd_mcu_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_dcd_mcu_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_dcd_mcu_init_lt_axi_s_awcache,
    input  dcd_pkg::dcd_mcu_init_lt_axi_id_t        i_dcd_mcu_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_dcd_mcu_init_lt_axi_s_awlen,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_dcd_mcu_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_dcd_mcu_init_lt_axi_s_awqos,
    output logic                                    o_dcd_mcu_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_dcd_mcu_init_lt_axi_s_awsize,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_awvalid,
    output dcd_pkg::dcd_mcu_init_lt_axi_id_t        o_dcd_mcu_init_lt_axi_s_bid,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_dcd_mcu_init_lt_axi_s_bresp,
    output logic                                    o_dcd_mcu_init_lt_axi_s_bvalid,
    input  dcd_pkg::dcd_mcu_init_lt_axi_data_t      i_dcd_mcu_init_lt_axi_s_wdata,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_wlast,
    output logic                                    o_dcd_mcu_init_lt_axi_s_wready,
    input  dcd_pkg::dcd_mcu_init_lt_axi_strb_t      i_dcd_mcu_init_lt_axi_s_wstrb,
    input  logic                                    i_dcd_mcu_init_lt_axi_s_wvalid,
    output logic                                    o_dcd_mcu_pwr_idle_val,
    output logic                                    o_dcd_mcu_pwr_idle_ack,
    input  logic                                    i_dcd_mcu_pwr_idle_req,
    input  wire                                     i_dcd_mcu_rst_n,
    output logic                                    o_dcd_pwr_idle_val,
    output logic                                    o_dcd_pwr_idle_ack,
    input  logic                                    i_dcd_pwr_idle_req,
    output dcd_pkg::dcd_targ_cfg_apb_addr_t         o_dcd_targ_cfg_apb_m_paddr,
    output logic                                    o_dcd_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_dcd_targ_cfg_apb_m_pprot,
    input  dcd_pkg::dcd_targ_cfg_apb_data_t         i_dcd_targ_cfg_apb_m_prdata,
    input  logic                                    i_dcd_targ_cfg_apb_m_pready,
    output logic                                    o_dcd_targ_cfg_apb_m_psel,
    input  logic                                    i_dcd_targ_cfg_apb_m_pslverr,
    output dcd_pkg::dcd_targ_cfg_apb_strb_t         o_dcd_targ_cfg_apb_m_pstrb,
    output dcd_pkg::dcd_targ_cfg_apb_data_t         o_dcd_targ_cfg_apb_m_pwdata,
    output logic                                    o_dcd_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_syscfg_addr_t             o_dcd_targ_syscfg_apb_m_paddr,
    output logic                                    o_dcd_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_dcd_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_dcd_targ_syscfg_apb_m_prdata,
    input  logic                                    i_dcd_targ_syscfg_apb_m_pready,
    output logic                                    o_dcd_targ_syscfg_apb_m_psel,
    input  logic                                    i_dcd_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_dcd_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_dcd_targ_syscfg_apb_m_pwdata,
    output logic                                    o_dcd_targ_syscfg_apb_m_pwrite,
    input  logic [686:0]                            i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld,
    output logic [108:0]                            o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld,
    input  logic [686:0]                            i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld,
    output logic [108:0]                            o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld,
    input  logic [146:0]                            i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld,
    output logic [686:0]                            o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld,
    input  logic [146:0]                            i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld,
    output logic [686:0]                            o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld,
    input  logic [182:0]                            i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data,
    input  logic                                    i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head,
    output logic                                    o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy,
    input  logic                                    i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail,
    input  logic                                    i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld,
    output logic [182:0]                            o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data,
    output logic                                    o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head,
    input  logic                                    i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy,
    output logic                                    o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail,
    output logic                                    o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld,
    input  logic [182:0]                            i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data,
    input  logic                                    i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head,
    output logic                                    o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy,
    input  logic                                    i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail,
    input  logic                                    i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld,
    output logic [182:0]                            o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data,
    output logic                                    o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head,
    input  logic                                    i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy,
    output logic                                    o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail,
    output logic                                    o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld,
    output logic [398:0]                            o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld,
    input  logic [398:0]                            i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld,
    output logic [398:0]                            o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld,
    input  logic [398:0]                            i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld,
    output logic [398:0]                            o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld,
    input  logic [398:0]                            i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld,
    output logic [398:0]                            o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld,
    input  logic [398:0]                            i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld,
    output logic [182:0]                            o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld,
    input  logic [182:0]                            i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld,
    output logic [686:0]                            o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld,
    input  logic [108:0]                            i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld,
    output logic [146:0]                            o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld,
    input  logic [686:0]                            i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld,
    output logic [182:0]                            o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data,
    output logic                                    o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head,
    input  logic                                    i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy,
    output logic                                    o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail,
    output logic                                    o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld,
    input  logic [182:0]                            i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data,
    input  logic                                    i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head,
    output logic                                    o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy,
    input  logic                                    i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail,
    input  logic                                    i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld,
    input  logic                                    i_l2_addr_mode_port_b0,
    input  logic                                    i_l2_addr_mode_port_b1,
    input  logic                                    i_l2_intr_mode_port_b0,
    input  logic                                    i_l2_intr_mode_port_b1,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e0_req_mainpde,
    output logic                                    lnk_buff_dec_128_to_256_ddr_e0_req_mainprn,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e0_req_mainret,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e0_req_mainse,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainpde,
    output logic                                    lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainprn,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainret,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainse,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e1_req_mainpde,
    output logic                                    lnk_buff_dec_128_to_256_ddr_e1_req_mainprn,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e1_req_mainret,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e1_req_mainse,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainpde,
    output logic                                    lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainprn,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainret,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainse,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e2_req_mainpde,
    output logic                                    lnk_buff_dec_128_to_256_ddr_e2_req_mainprn,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e2_req_mainret,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e2_req_mainse,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainpde,
    output logic                                    lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainprn,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainret,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainse,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e3_req_mainpde,
    output logic                                    lnk_buff_dec_128_to_256_ddr_e3_req_mainprn,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e3_req_mainret,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e3_req_mainse,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainpde,
    output logic                                    lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainprn,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainret,
    input  logic                                    lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainse,
    input  logic                                    lnk_buff_soc_128_to_256_lt_req_mainpde,
    output logic                                    lnk_buff_soc_128_to_256_lt_req_mainprn,
    input  logic                                    lnk_buff_soc_128_to_256_lt_req_mainret,
    input  logic                                    lnk_buff_soc_128_to_256_lt_req_mainse,
    input  logic                                    lnk_buff_soc_128_to_256_lt_req_resp_mainpde,
    output logic                                    lnk_buff_soc_128_to_256_lt_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_128_to_256_lt_req_resp_mainret,
    input  logic                                    lnk_buff_soc_128_to_256_lt_req_resp_mainse,
    input  logic                                    lnk_buff_soc_128_to_256_rd_req_resp_mainpde,
    output logic                                    lnk_buff_soc_128_to_256_rd_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_128_to_256_rd_req_resp_mainret,
    input  logic                                    lnk_buff_soc_128_to_256_rd_req_resp_mainse,
    input  logic                                    lnk_buff_soc_128_to_256_wr_req_mainpde,
    output logic                                    lnk_buff_soc_128_to_256_wr_req_mainprn,
    input  logic                                    lnk_buff_soc_128_to_256_wr_req_mainret,
    input  logic                                    lnk_buff_soc_128_to_256_wr_req_mainse,
    input  logic                                    lnk_buff_soc_128_to_64_req_mainpde,
    output logic                                    lnk_buff_soc_128_to_64_req_mainprn,
    input  logic                                    lnk_buff_soc_128_to_64_req_mainret,
    input  logic                                    lnk_buff_soc_128_to_64_req_mainse,
    input  logic                                    lnk_buff_soc_128_to_64_req_resp_mainpde,
    output logic                                    lnk_buff_soc_128_to_64_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_128_to_64_req_resp_mainret,
    input  logic                                    lnk_buff_soc_128_to_64_req_resp_mainse,
    input  logic                                    lnk_buff_soc_256_to_128_rd_req_resp_mainpde,
    output logic                                    lnk_buff_soc_256_to_128_rd_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_256_to_128_rd_req_resp_mainret,
    input  logic                                    lnk_buff_soc_256_to_128_rd_req_resp_mainse,
    input  logic                                    lnk_buff_soc_256_to_128_wr_req_mainpde,
    output logic                                    lnk_buff_soc_256_to_128_wr_req_mainprn,
    input  logic                                    lnk_buff_soc_256_to_128_wr_req_mainret,
    input  logic                                    lnk_buff_soc_256_to_128_wr_req_mainse,
    input  logic                                    lnk_buff_soc_256_to_512_rd_req_resp_mainpde,
    output logic                                    lnk_buff_soc_256_to_512_rd_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_256_to_512_rd_req_resp_mainret,
    input  logic                                    lnk_buff_soc_256_to_512_rd_req_resp_mainse,
    input  logic                                    lnk_buff_soc_256_to_512_wr_req_mainpde,
    output logic                                    lnk_buff_soc_256_to_512_wr_req_mainprn,
    input  logic                                    lnk_buff_soc_256_to_512_wr_req_mainret,
    input  logic                                    lnk_buff_soc_256_to_512_wr_req_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e0_req_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_ddr_e0_req_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e0_req_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e0_req_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e1_req_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_ddr_e1_req_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e1_req_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e1_req_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e2_req_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_ddr_e2_req_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e2_req_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e2_req_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e3_req_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_ddr_e3_req_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e3_req_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e3_req_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_rd_req_resp_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_rd_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_rd_req_resp_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_rd_req_resp_mainse,
    input  logic                                    lnk_buff_soc_512_to_256_wr_req_mainpde,
    output logic                                    lnk_buff_soc_512_to_256_wr_req_mainprn,
    input  logic                                    lnk_buff_soc_512_to_256_wr_req_mainret,
    input  logic                                    lnk_buff_soc_512_to_256_wr_req_mainse,
    input  logic                                    lnk_buff_soc_64_to_128_lt_req_mainpde,
    output logic                                    lnk_buff_soc_64_to_128_lt_req_mainprn,
    input  logic                                    lnk_buff_soc_64_to_128_lt_req_mainret,
    input  logic                                    lnk_buff_soc_64_to_128_lt_req_mainse,
    input  logic                                    lnk_buff_soc_64_to_128_lt_req_resp_mainpde,
    output logic                                    lnk_buff_soc_64_to_128_lt_req_resp_mainprn,
    input  logic                                    lnk_buff_soc_64_to_128_lt_req_resp_mainret,
    input  logic                                    lnk_buff_soc_64_to_128_lt_req_resp_mainse,
    input  logic                                    i_lpddr_graph_addr_mode_port_b0,
    input  logic                                    i_lpddr_graph_addr_mode_port_b1,
    input  logic                                    i_lpddr_graph_intr_mode_port_b0,
    input  logic                                    i_lpddr_graph_intr_mode_port_b1,
    input  logic                                    i_lpddr_ppp_addr_mode_port_b0,
    input  logic                                    i_lpddr_ppp_addr_mode_port_b1,
    input  logic                                    i_lpddr_ppp_intr_mode_port_b0,
    input  logic                                    i_lpddr_ppp_intr_mode_port_b1,
    input  wire                                     i_noc_clk,
    input  wire                                     i_noc_rst_n,
    input  wire                                     i_pcie_aon_clk,
    input  wire                                     i_pcie_aon_rst_n,
    input  wire                                     i_pcie_init_mt_clk,
    input  wire                                     i_pcie_init_mt_clken,
    output logic                                    o_pcie_init_mt_pwr_idle_val,
    output logic                                    o_pcie_init_mt_pwr_idle_ack,
    input  logic                                    i_pcie_init_mt_pwr_idle_req,
    input  chip_pkg::chip_axi_addr_t                i_pcie_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pcie_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pcie_init_mt_axi_s_arcache,
    input  pcie_pkg::pcie_init_mt_axi_id_t          i_pcie_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pcie_init_mt_axi_s_arlen,
    input  logic                                    i_pcie_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pcie_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_pcie_init_mt_axi_s_arqos,
    output logic                                    o_pcie_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pcie_init_mt_axi_s_arsize,
    input  logic                                    i_pcie_init_mt_axi_s_arvalid,
    output pcie_pkg::pcie_init_mt_axi_data_t        o_pcie_init_mt_axi_s_rdata,
    output pcie_pkg::pcie_init_mt_axi_id_t          o_pcie_init_mt_axi_s_rid,
    output logic                                    o_pcie_init_mt_axi_s_rlast,
    input  logic                                    i_pcie_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pcie_init_mt_axi_s_rresp,
    output logic                                    o_pcie_init_mt_axi_s_rvalid,
    input  wire                                     i_pcie_init_mt_rst_n,
    input  chip_pkg::chip_axi_addr_t                i_pcie_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pcie_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pcie_init_mt_axi_s_awcache,
    input  pcie_pkg::pcie_init_mt_axi_id_t          i_pcie_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pcie_init_mt_axi_s_awlen,
    input  logic                                    i_pcie_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pcie_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_pcie_init_mt_axi_s_awqos,
    output logic                                    o_pcie_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pcie_init_mt_axi_s_awsize,
    input  logic                                    i_pcie_init_mt_axi_s_awvalid,
    output pcie_pkg::pcie_init_mt_axi_id_t          o_pcie_init_mt_axi_s_bid,
    input  logic                                    i_pcie_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pcie_init_mt_axi_s_bresp,
    output logic                                    o_pcie_init_mt_axi_s_bvalid,
    input  pcie_pkg::pcie_init_mt_axi_data_t        i_pcie_init_mt_axi_s_wdata,
    input  logic                                    i_pcie_init_mt_axi_s_wlast,
    output logic                                    o_pcie_init_mt_axi_s_wready,
    input  pcie_pkg::pcie_init_mt_axi_strb_t        i_pcie_init_mt_axi_s_wstrb,
    input  logic                                    i_pcie_init_mt_axi_s_wvalid,
    output pcie_pkg::pcie_targ_cfg_apb3_addr_t      o_pcie_targ_cfg_apb_m_paddr,
    output logic                                    o_pcie_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_pcie_targ_cfg_apb_m_pprot,
    input  pcie_pkg::pcie_targ_cfg_apb3_data_t      i_pcie_targ_cfg_apb_m_prdata,
    input  logic                                    i_pcie_targ_cfg_apb_m_pready,
    output logic                                    o_pcie_targ_cfg_apb_m_psel,
    input  logic                                    i_pcie_targ_cfg_apb_m_pslverr,
    output logic [3:0]                              o_pcie_targ_cfg_apb_m_pstrb,
    output pcie_pkg::pcie_targ_cfg_apb3_data_t      o_pcie_targ_cfg_apb_m_pwdata,
    output logic                                    o_pcie_targ_cfg_apb_m_pwrite,
    input  wire                                     i_pcie_targ_cfg_clk,
    input  wire                                     i_pcie_targ_cfg_clken,
    output chip_pkg::chip_axi_addr_t                o_pcie_targ_cfg_dbi_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_pcie_targ_cfg_dbi_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_pcie_targ_cfg_dbi_axi_m_arcache,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_id_t     o_pcie_targ_cfg_dbi_axi_m_arid,
    output axi_pkg::axi_len_t                       o_pcie_targ_cfg_dbi_axi_m_arlen,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_pcie_targ_cfg_dbi_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_pcie_targ_cfg_dbi_axi_m_arqos,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_arready,
    output axi_pkg::axi_size_t                      o_pcie_targ_cfg_dbi_axi_m_arsize,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_pcie_targ_cfg_dbi_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_pcie_targ_cfg_dbi_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_pcie_targ_cfg_dbi_axi_m_awcache,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_id_t     o_pcie_targ_cfg_dbi_axi_m_awid,
    output axi_pkg::axi_len_t                       o_pcie_targ_cfg_dbi_axi_m_awlen,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_pcie_targ_cfg_dbi_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_pcie_targ_cfg_dbi_axi_m_awqos,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_awready,
    output axi_pkg::axi_size_t                      o_pcie_targ_cfg_dbi_axi_m_awsize,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_awvalid,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_id_t     i_pcie_targ_cfg_dbi_axi_m_bid,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_pcie_targ_cfg_dbi_axi_m_bresp,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_bvalid,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_data_t   i_pcie_targ_cfg_dbi_axi_m_rdata,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_id_t     i_pcie_targ_cfg_dbi_axi_m_rid,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_rlast,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_pcie_targ_cfg_dbi_axi_m_rresp,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_rvalid,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_data_t   o_pcie_targ_cfg_dbi_axi_m_wdata,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_wlast,
    input  logic                                    i_pcie_targ_cfg_dbi_axi_m_wready,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_strb_t   o_pcie_targ_cfg_dbi_axi_m_wstrb,
    output logic                                    o_pcie_targ_cfg_dbi_axi_m_wvalid,
    input  wire                                     i_pcie_targ_cfg_dbi_clk,
    input  wire                                     i_pcie_targ_cfg_dbi_clken,
    output logic                                    o_pcie_targ_cfg_dbi_pwr_idle_val,
    output logic                                    o_pcie_targ_cfg_dbi_pwr_idle_ack,
    input  logic                                    i_pcie_targ_cfg_dbi_pwr_idle_req,
    input  wire                                     i_pcie_targ_cfg_dbi_rst_n,
    output logic                                    o_pcie_targ_cfg_pwr_idle_val,
    output logic                                    o_pcie_targ_cfg_pwr_idle_ack,
    input  logic                                    i_pcie_targ_cfg_pwr_idle_req,
    input  wire                                     i_pcie_targ_cfg_rst_n,
    input  wire                                     i_pcie_targ_mt_clk,
    input  wire                                     i_pcie_targ_mt_clken,
    output logic                                    o_pcie_targ_mt_pwr_idle_val,
    output logic                                    o_pcie_targ_mt_pwr_idle_ack,
    input  logic                                    i_pcie_targ_mt_pwr_idle_req,
    output chip_pkg::chip_axi_addr_t                o_pcie_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_pcie_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_pcie_targ_mt_axi_m_arcache,
    output pcie_pkg::pcie_targ_mt_axi_id_t          o_pcie_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_pcie_targ_mt_axi_m_arlen,
    output logic                                    o_pcie_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_pcie_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_pcie_targ_mt_axi_m_arqos,
    input  logic                                    i_pcie_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_pcie_targ_mt_axi_m_arsize,
    output logic                                    o_pcie_targ_mt_axi_m_arvalid,
    input  pcie_pkg::pcie_targ_mt_axi_data_t        i_pcie_targ_mt_axi_m_rdata,
    input  pcie_pkg::pcie_targ_mt_axi_id_t          i_pcie_targ_mt_axi_m_rid,
    input  logic                                    i_pcie_targ_mt_axi_m_rlast,
    output logic                                    o_pcie_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_pcie_targ_mt_axi_m_rresp,
    input  logic                                    i_pcie_targ_mt_axi_m_rvalid,
    input  wire                                     i_pcie_targ_mt_rst_n,
    output chip_pkg::chip_axi_addr_t                o_pcie_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_pcie_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_pcie_targ_mt_axi_m_awcache,
    output pcie_pkg::pcie_targ_mt_axi_id_t          o_pcie_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_pcie_targ_mt_axi_m_awlen,
    output logic                                    o_pcie_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_pcie_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_pcie_targ_mt_axi_m_awqos,
    input  logic                                    i_pcie_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_pcie_targ_mt_axi_m_awsize,
    output logic                                    o_pcie_targ_mt_axi_m_awvalid,
    input  pcie_pkg::pcie_targ_mt_axi_id_t          i_pcie_targ_mt_axi_m_bid,
    output logic                                    o_pcie_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_pcie_targ_mt_axi_m_bresp,
    input  logic                                    i_pcie_targ_mt_axi_m_bvalid,
    output pcie_pkg::pcie_targ_mt_axi_data_t        o_pcie_targ_mt_axi_m_wdata,
    output logic                                    o_pcie_targ_mt_axi_m_wlast,
    input  logic                                    i_pcie_targ_mt_axi_m_wready,
    output pcie_pkg::pcie_targ_mt_axi_strb_t        o_pcie_targ_mt_axi_m_wstrb,
    output logic                                    o_pcie_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_pcie_targ_syscfg_apb_m_paddr,
    output logic                                    o_pcie_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_pcie_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_pcie_targ_syscfg_apb_m_prdata,
    input  logic                                    i_pcie_targ_syscfg_apb_m_pready,
    output logic                                    o_pcie_targ_syscfg_apb_m_psel,
    input  logic                                    i_pcie_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_pcie_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_pcie_targ_syscfg_apb_m_pwdata,
    output logic                                    o_pcie_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_pve_0_aon_clk,
    input  wire                                     i_pve_0_aon_rst_n,
    input  wire                                     i_pve_0_clk,
    input  wire                                     i_pve_0_clken,
    input  chip_pkg::chip_axi_addr_t                i_pve_0_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pve_0_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pve_0_init_ht_axi_s_arcache,
    input  pve_pkg::pve_ht_axi_m_id_t               i_pve_0_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pve_0_init_ht_axi_s_arlen,
    input  logic                                    i_pve_0_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pve_0_init_ht_axi_s_arprot,
    output logic                                    o_pve_0_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pve_0_init_ht_axi_s_arsize,
    input  logic                                    i_pve_0_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t             o_pve_0_init_ht_axi_s_rdata,
    output pve_pkg::pve_ht_axi_m_id_t               o_pve_0_init_ht_axi_s_rid,
    output logic                                    o_pve_0_init_ht_axi_s_rlast,
    input  logic                                    i_pve_0_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pve_0_init_ht_axi_s_rresp,
    output logic                                    o_pve_0_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_0_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pve_0_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pve_0_init_ht_axi_s_awcache,
    input  pve_pkg::pve_ht_axi_m_id_t               i_pve_0_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pve_0_init_ht_axi_s_awlen,
    input  logic                                    i_pve_0_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pve_0_init_ht_axi_s_awprot,
    output logic                                    o_pve_0_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pve_0_init_ht_axi_s_awsize,
    input  logic                                    i_pve_0_init_ht_axi_s_awvalid,
    output pve_pkg::pve_ht_axi_m_id_t               o_pve_0_init_ht_axi_s_bid,
    input  logic                                    i_pve_0_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pve_0_init_ht_axi_s_bresp,
    output logic                                    o_pve_0_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t             i_pve_0_init_ht_axi_s_wdata,
    input  logic                                    i_pve_0_init_ht_axi_s_wlast,
    output logic                                    o_pve_0_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t            i_pve_0_init_ht_axi_s_wstrb,
    input  logic                                    i_pve_0_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_0_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pve_0_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pve_0_init_lt_axi_s_arcache,
    input  pve_pkg::pve_lt_axi_m_id_t               i_pve_0_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pve_0_init_lt_axi_s_arlen,
    input  logic                                    i_pve_0_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pve_0_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_pve_0_init_lt_axi_s_arqos,
    output logic                                    o_pve_0_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pve_0_init_lt_axi_s_arsize,
    input  logic                                    i_pve_0_init_lt_axi_s_arvalid,
    output chip_pkg::chip_axi_lt_data_t             o_pve_0_init_lt_axi_s_rdata,
    output pve_pkg::pve_lt_axi_m_id_t               o_pve_0_init_lt_axi_s_rid,
    output logic                                    o_pve_0_init_lt_axi_s_rlast,
    input  logic                                    i_pve_0_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pve_0_init_lt_axi_s_rresp,
    output logic                                    o_pve_0_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_0_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pve_0_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pve_0_init_lt_axi_s_awcache,
    input  pve_pkg::pve_lt_axi_m_id_t               i_pve_0_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pve_0_init_lt_axi_s_awlen,
    input  logic                                    i_pve_0_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pve_0_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_pve_0_init_lt_axi_s_awqos,
    output logic                                    o_pve_0_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pve_0_init_lt_axi_s_awsize,
    input  logic                                    i_pve_0_init_lt_axi_s_awvalid,
    output pve_pkg::pve_lt_axi_m_id_t               o_pve_0_init_lt_axi_s_bid,
    input  logic                                    i_pve_0_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pve_0_init_lt_axi_s_bresp,
    output logic                                    o_pve_0_init_lt_axi_s_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_pve_0_init_lt_axi_s_wdata,
    input  logic                                    i_pve_0_init_lt_axi_s_wlast,
    output logic                                    o_pve_0_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t            i_pve_0_init_lt_axi_s_wstrb,
    input  logic                                    i_pve_0_init_lt_axi_s_wvalid,
    output logic                                    o_pve_0_pwr_idle_val,
    output logic                                    o_pve_0_pwr_idle_ack,
    input  logic                                    i_pve_0_pwr_idle_req,
    input  wire                                     i_pve_0_rst_n,
    output chip_pkg::chip_axi_addr_t                o_pve_0_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_pve_0_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_pve_0_targ_lt_axi_m_arcache,
    output pve_pkg::pve_lt_axi_s_id_t               o_pve_0_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_pve_0_targ_lt_axi_m_arlen,
    output logic                                    o_pve_0_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_pve_0_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_pve_0_targ_lt_axi_m_arqos,
    input  logic                                    i_pve_0_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_pve_0_targ_lt_axi_m_arsize,
    output logic                                    o_pve_0_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_pve_0_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_pve_0_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_pve_0_targ_lt_axi_m_awcache,
    output pve_pkg::pve_lt_axi_s_id_t               o_pve_0_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_pve_0_targ_lt_axi_m_awlen,
    output logic                                    o_pve_0_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_pve_0_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_pve_0_targ_lt_axi_m_awqos,
    input  logic                                    i_pve_0_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_pve_0_targ_lt_axi_m_awsize,
    output logic                                    o_pve_0_targ_lt_axi_m_awvalid,
    input  pve_pkg::pve_lt_axi_s_id_t               i_pve_0_targ_lt_axi_m_bid,
    output logic                                    o_pve_0_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_pve_0_targ_lt_axi_m_bresp,
    input  logic                                    i_pve_0_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_pve_0_targ_lt_axi_m_rdata,
    input  pve_pkg::pve_lt_axi_s_id_t               i_pve_0_targ_lt_axi_m_rid,
    input  logic                                    i_pve_0_targ_lt_axi_m_rlast,
    output logic                                    o_pve_0_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_pve_0_targ_lt_axi_m_rresp,
    input  logic                                    i_pve_0_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_pve_0_targ_lt_axi_m_wdata,
    output logic                                    o_pve_0_targ_lt_axi_m_wlast,
    input  logic                                    i_pve_0_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_pve_0_targ_lt_axi_m_wstrb,
    output logic                                    o_pve_0_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_pve_0_targ_syscfg_apb_m_paddr,
    output logic                                    o_pve_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_pve_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_pve_0_targ_syscfg_apb_m_prdata,
    input  logic                                    i_pve_0_targ_syscfg_apb_m_pready,
    output logic                                    o_pve_0_targ_syscfg_apb_m_psel,
    input  logic                                    i_pve_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_pve_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_pve_0_targ_syscfg_apb_m_pwdata,
    output logic                                    o_pve_0_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_pve_1_aon_clk,
    input  wire                                     i_pve_1_aon_rst_n,
    input  wire                                     i_pve_1_clk,
    input  wire                                     i_pve_1_clken,
    input  chip_pkg::chip_axi_addr_t                i_pve_1_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pve_1_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pve_1_init_ht_axi_s_arcache,
    input  pve_pkg::pve_ht_axi_m_id_t               i_pve_1_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pve_1_init_ht_axi_s_arlen,
    input  logic                                    i_pve_1_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pve_1_init_ht_axi_s_arprot,
    output logic                                    o_pve_1_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pve_1_init_ht_axi_s_arsize,
    input  logic                                    i_pve_1_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t             o_pve_1_init_ht_axi_s_rdata,
    output pve_pkg::pve_ht_axi_m_id_t               o_pve_1_init_ht_axi_s_rid,
    output logic                                    o_pve_1_init_ht_axi_s_rlast,
    input  logic                                    i_pve_1_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pve_1_init_ht_axi_s_rresp,
    output logic                                    o_pve_1_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_1_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pve_1_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pve_1_init_ht_axi_s_awcache,
    input  pve_pkg::pve_ht_axi_m_id_t               i_pve_1_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pve_1_init_ht_axi_s_awlen,
    input  logic                                    i_pve_1_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pve_1_init_ht_axi_s_awprot,
    output logic                                    o_pve_1_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pve_1_init_ht_axi_s_awsize,
    input  logic                                    i_pve_1_init_ht_axi_s_awvalid,
    output pve_pkg::pve_ht_axi_m_id_t               o_pve_1_init_ht_axi_s_bid,
    input  logic                                    i_pve_1_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pve_1_init_ht_axi_s_bresp,
    output logic                                    o_pve_1_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t             i_pve_1_init_ht_axi_s_wdata,
    input  logic                                    i_pve_1_init_ht_axi_s_wlast,
    output logic                                    o_pve_1_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t            i_pve_1_init_ht_axi_s_wstrb,
    input  logic                                    i_pve_1_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_1_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_pve_1_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_pve_1_init_lt_axi_s_arcache,
    input  pve_pkg::pve_lt_axi_m_id_t               i_pve_1_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_pve_1_init_lt_axi_s_arlen,
    input  logic                                    i_pve_1_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_pve_1_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_pve_1_init_lt_axi_s_arqos,
    output logic                                    o_pve_1_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_pve_1_init_lt_axi_s_arsize,
    input  logic                                    i_pve_1_init_lt_axi_s_arvalid,
    output chip_pkg::chip_axi_lt_data_t             o_pve_1_init_lt_axi_s_rdata,
    output pve_pkg::pve_lt_axi_m_id_t               o_pve_1_init_lt_axi_s_rid,
    output logic                                    o_pve_1_init_lt_axi_s_rlast,
    input  logic                                    i_pve_1_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_pve_1_init_lt_axi_s_rresp,
    output logic                                    o_pve_1_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                i_pve_1_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_pve_1_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_pve_1_init_lt_axi_s_awcache,
    input  pve_pkg::pve_lt_axi_m_id_t               i_pve_1_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_pve_1_init_lt_axi_s_awlen,
    input  logic                                    i_pve_1_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_pve_1_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_pve_1_init_lt_axi_s_awqos,
    output logic                                    o_pve_1_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_pve_1_init_lt_axi_s_awsize,
    input  logic                                    i_pve_1_init_lt_axi_s_awvalid,
    output pve_pkg::pve_lt_axi_m_id_t               o_pve_1_init_lt_axi_s_bid,
    input  logic                                    i_pve_1_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_pve_1_init_lt_axi_s_bresp,
    output logic                                    o_pve_1_init_lt_axi_s_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_pve_1_init_lt_axi_s_wdata,
    input  logic                                    i_pve_1_init_lt_axi_s_wlast,
    output logic                                    o_pve_1_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t            i_pve_1_init_lt_axi_s_wstrb,
    input  logic                                    i_pve_1_init_lt_axi_s_wvalid,
    output logic                                    o_pve_1_pwr_idle_val,
    output logic                                    o_pve_1_pwr_idle_ack,
    input  logic                                    i_pve_1_pwr_idle_req,
    input  wire                                     i_pve_1_rst_n,
    output chip_pkg::chip_axi_addr_t                o_pve_1_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_pve_1_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_pve_1_targ_lt_axi_m_arcache,
    output pve_pkg::pve_lt_axi_s_id_t               o_pve_1_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_pve_1_targ_lt_axi_m_arlen,
    output logic                                    o_pve_1_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_pve_1_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_pve_1_targ_lt_axi_m_arqos,
    input  logic                                    i_pve_1_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_pve_1_targ_lt_axi_m_arsize,
    output logic                                    o_pve_1_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_pve_1_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_pve_1_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_pve_1_targ_lt_axi_m_awcache,
    output pve_pkg::pve_lt_axi_s_id_t               o_pve_1_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_pve_1_targ_lt_axi_m_awlen,
    output logic                                    o_pve_1_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_pve_1_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_pve_1_targ_lt_axi_m_awqos,
    input  logic                                    i_pve_1_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_pve_1_targ_lt_axi_m_awsize,
    output logic                                    o_pve_1_targ_lt_axi_m_awvalid,
    input  pve_pkg::pve_lt_axi_s_id_t               i_pve_1_targ_lt_axi_m_bid,
    output logic                                    o_pve_1_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_pve_1_targ_lt_axi_m_bresp,
    input  logic                                    i_pve_1_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_pve_1_targ_lt_axi_m_rdata,
    input  pve_pkg::pve_lt_axi_s_id_t               i_pve_1_targ_lt_axi_m_rid,
    input  logic                                    i_pve_1_targ_lt_axi_m_rlast,
    output logic                                    o_pve_1_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_pve_1_targ_lt_axi_m_rresp,
    input  logic                                    i_pve_1_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_pve_1_targ_lt_axi_m_wdata,
    output logic                                    o_pve_1_targ_lt_axi_m_wlast,
    input  logic                                    i_pve_1_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_pve_1_targ_lt_axi_m_wstrb,
    output logic                                    o_pve_1_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_pve_1_targ_syscfg_apb_m_paddr,
    output logic                                    o_pve_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_pve_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_pve_1_targ_syscfg_apb_m_prdata,
    input  logic                                    i_pve_1_targ_syscfg_apb_m_pready,
    output logic                                    o_pve_1_targ_syscfg_apb_m_psel,
    input  logic                                    i_pve_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_pve_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_pve_1_targ_syscfg_apb_m_pwdata,
    output logic                                    o_pve_1_targ_syscfg_apb_m_pwrite,
    input  logic                                    scan_en,
    input  wire                                     i_soc_mgmt_aon_clk,
    input  wire                                     i_soc_mgmt_aon_rst_n,
    input  wire                                     i_soc_mgmt_clk,
    input  wire                                     i_soc_mgmt_clken,
    input  chip_pkg::chip_axi_addr_t                i_soc_mgmt_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                     i_soc_mgmt_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                     i_soc_mgmt_init_lt_axi_s_arcache,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t     i_soc_mgmt_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                       i_soc_mgmt_init_lt_axi_s_arlen,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                      i_soc_mgmt_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                       i_soc_mgmt_init_lt_axi_s_arqos,
    output logic                                    o_soc_mgmt_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                      i_soc_mgmt_init_lt_axi_s_arsize,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                i_soc_mgmt_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                     i_soc_mgmt_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                     i_soc_mgmt_init_lt_axi_s_awcache,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t     i_soc_mgmt_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                       i_soc_mgmt_init_lt_axi_s_awlen,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                      i_soc_mgmt_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                       i_soc_mgmt_init_lt_axi_s_awqos,
    output logic                                    o_soc_mgmt_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                      i_soc_mgmt_init_lt_axi_s_awsize,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_awvalid,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t     o_soc_mgmt_init_lt_axi_s_bid,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                      o_soc_mgmt_init_lt_axi_s_bresp,
    output logic                                    o_soc_mgmt_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t             o_soc_mgmt_init_lt_axi_s_rdata,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t     o_soc_mgmt_init_lt_axi_s_rid,
    output logic                                    o_soc_mgmt_init_lt_axi_s_rlast,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                      o_soc_mgmt_init_lt_axi_s_rresp,
    output logic                                    o_soc_mgmt_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_soc_mgmt_init_lt_axi_s_wdata,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_wlast,
    output logic                                    o_soc_mgmt_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t            i_soc_mgmt_init_lt_axi_s_wstrb,
    input  logic                                    i_soc_mgmt_init_lt_axi_s_wvalid,
    output logic                                    o_soc_mgmt_pwr_idle_val,
    output logic                                    o_soc_mgmt_pwr_idle_ack,
    input  logic                                    i_soc_mgmt_pwr_idle_req,
    input  wire                                     i_soc_mgmt_rst_n,
    output chip_pkg::chip_axi_addr_t                o_soc_mgmt_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_soc_mgmt_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_soc_mgmt_targ_lt_axi_m_arcache,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t     o_soc_mgmt_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_soc_mgmt_targ_lt_axi_m_arlen,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_soc_mgmt_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_soc_mgmt_targ_lt_axi_m_arqos,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_soc_mgmt_targ_lt_axi_m_arsize,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_soc_mgmt_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_soc_mgmt_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_soc_mgmt_targ_lt_axi_m_awcache,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t     o_soc_mgmt_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_soc_mgmt_targ_lt_axi_m_awlen,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_soc_mgmt_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_soc_mgmt_targ_lt_axi_m_awqos,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_soc_mgmt_targ_lt_axi_m_awsize,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_awvalid,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t     i_soc_mgmt_targ_lt_axi_m_bid,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_soc_mgmt_targ_lt_axi_m_bresp,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_soc_mgmt_targ_lt_axi_m_rdata,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t     i_soc_mgmt_targ_lt_axi_m_rid,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_rlast,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_soc_mgmt_targ_lt_axi_m_rresp,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_soc_mgmt_targ_lt_axi_m_wdata,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_wlast,
    input  logic                                    i_soc_mgmt_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_soc_mgmt_targ_lt_axi_m_wstrb,
    output logic                                    o_soc_mgmt_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_soc_mgmt_syscfg_addr_t    o_soc_mgmt_targ_syscfg_apb_m_paddr,
    output logic                                    o_soc_mgmt_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_soc_mgmt_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_soc_mgmt_targ_syscfg_apb_m_prdata,
    input  logic                                    i_soc_mgmt_targ_syscfg_apb_m_pready,
    output logic                                    o_soc_mgmt_targ_syscfg_apb_m_psel,
    input  logic                                    i_soc_mgmt_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_soc_mgmt_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_soc_mgmt_targ_syscfg_apb_m_pwdata,
    output logic                                    o_soc_mgmt_targ_syscfg_apb_m_pwrite,
    input  wire                                     i_sys_spm_aon_clk,
    input  wire                                     i_sys_spm_aon_rst_n,
    input  wire                                     i_sys_spm_clk,
    input  wire                                     i_sys_spm_clken,
    output logic                                    o_sys_spm_pwr_idle_val,
    output logic                                    o_sys_spm_pwr_idle_ack,
    input  logic                                    i_sys_spm_pwr_idle_req,
    input  wire                                     i_sys_spm_rst_n,
    output chip_pkg::chip_axi_addr_t                o_sys_spm_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                     o_sys_spm_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                     o_sys_spm_targ_lt_axi_m_arcache,
    output sys_spm_pkg::sys_spm_targ_lt_axi_id_t    o_sys_spm_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                       o_sys_spm_targ_lt_axi_m_arlen,
    output logic                                    o_sys_spm_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                      o_sys_spm_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                       o_sys_spm_targ_lt_axi_m_arqos,
    input  logic                                    i_sys_spm_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                      o_sys_spm_targ_lt_axi_m_arsize,
    output logic                                    o_sys_spm_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                o_sys_spm_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                     o_sys_spm_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                     o_sys_spm_targ_lt_axi_m_awcache,
    output sys_spm_pkg::sys_spm_targ_lt_axi_id_t    o_sys_spm_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                       o_sys_spm_targ_lt_axi_m_awlen,
    output logic                                    o_sys_spm_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                      o_sys_spm_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                       o_sys_spm_targ_lt_axi_m_awqos,
    input  logic                                    i_sys_spm_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                      o_sys_spm_targ_lt_axi_m_awsize,
    output logic                                    o_sys_spm_targ_lt_axi_m_awvalid,
    input  sys_spm_pkg::sys_spm_targ_lt_axi_id_t    i_sys_spm_targ_lt_axi_m_bid,
    output logic                                    o_sys_spm_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                      i_sys_spm_targ_lt_axi_m_bresp,
    input  logic                                    i_sys_spm_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t             i_sys_spm_targ_lt_axi_m_rdata,
    input  sys_spm_pkg::sys_spm_targ_lt_axi_id_t    i_sys_spm_targ_lt_axi_m_rid,
    input  logic                                    i_sys_spm_targ_lt_axi_m_rlast,
    output logic                                    o_sys_spm_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                      i_sys_spm_targ_lt_axi_m_rresp,
    input  logic                                    i_sys_spm_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t             o_sys_spm_targ_lt_axi_m_wdata,
    output logic                                    o_sys_spm_targ_lt_axi_m_wlast,
    input  logic                                    i_sys_spm_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t            o_sys_spm_targ_lt_axi_m_wstrb,
    output logic                                    o_sys_spm_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t             o_sys_spm_targ_syscfg_apb_m_paddr,
    output logic                                    o_sys_spm_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                  o_sys_spm_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t         i_sys_spm_targ_syscfg_apb_m_prdata,
    input  logic                                    i_sys_spm_targ_syscfg_apb_m_pready,
    output logic                                    o_sys_spm_targ_syscfg_apb_m_psel,
    input  logic                                    i_sys_spm_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t         o_sys_spm_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t         o_sys_spm_targ_syscfg_apb_m_pwdata,
    output logic                                    o_sys_spm_targ_syscfg_apb_m_pwrite
);

    // TODO(psarras/joao; tidy up -- do we keep this patch floating or move to a separate design?)
    // TODO(psarras/joao; assert that Exclusives are only issued for the listed IDs)

    // APU RTL Patch for multiple outstanding Exclusives
    logic [2:0] apu_init_lt_axi_s_aruser;
    logic [2:0] apu_init_lt_axi_s_awuser;

    localparam apu_pkg::apu_axi_lt_m_id_t APU_0_AXID = 'h03;
    localparam apu_pkg::apu_axi_lt_m_id_t APU_1_AXID = 'h07;
    localparam apu_pkg::apu_axi_lt_m_id_t APU_2_AXID = 'h0b;
    localparam apu_pkg::apu_axi_lt_m_id_t APU_3_AXID = 'h0f;
    localparam apu_pkg::apu_axi_lt_m_id_t APU_4_AXID = 'h13;
    localparam apu_pkg::apu_axi_lt_m_id_t APU_5_AXID = 'h17;

    always_comb begin
      case(i_apu_init_lt_axi_s_arid)
        APU_0_AXID : apu_init_lt_axi_s_aruser = 3'h0;
        APU_1_AXID : apu_init_lt_axi_s_aruser = 3'h1;
        APU_2_AXID : apu_init_lt_axi_s_aruser = 3'h2;
        APU_3_AXID : apu_init_lt_axi_s_aruser = 3'h3;
        APU_4_AXID : apu_init_lt_axi_s_aruser = 3'h4;
        APU_5_AXID : apu_init_lt_axi_s_aruser = 3'h5;
        default: apu_init_lt_axi_s_aruser = 3'h0;
      endcase
    end

    always_comb begin
      case(i_apu_init_lt_axi_s_awid)
        APU_0_AXID : apu_init_lt_axi_s_awuser = 3'h0;
        APU_1_AXID : apu_init_lt_axi_s_awuser = 3'h1;
        APU_2_AXID : apu_init_lt_axi_s_awuser = 3'h2;
        APU_3_AXID : apu_init_lt_axi_s_awuser = 3'h3;
        APU_4_AXID : apu_init_lt_axi_s_awuser = 3'h4;
        APU_5_AXID : apu_init_lt_axi_s_awuser = 3'h5;
        default: apu_init_lt_axi_s_awuser = 3'h0;
      endcase
    end

    // PVE RTL Patch for multiple outstanding Exclusives
    // - Applying guidance from : https://git.axelera.ai/prod/europa/-/issues/2166#note_288387
    //      > it seems that pve_fabric does direct 1:1 mapping so 4 MSBs of AxID directly correspond to CPUID. 4 LSBs are 0x0, 0x7 or 0xB typically.

    // - PVE0
    logic [2:0] pve_0_init_lt_axi_s_aruser;
    logic [2:0] pve_0_init_lt_axi_s_awuser;
    logic [2:0] pve_1_init_lt_axi_s_aruser;
    logic [2:0] pve_1_init_lt_axi_s_awuser;

    // --------------------------------------------------
    //              SWITCH FIX ON AND OFF
    // --------------------------------------------------
    localparam EN_EX_PVE_FIX = 1;
    // --------------------------------------------------
    //              SWITCH FIX ON AND OFF
    // --------------------------------------------------

    // ----------
    if(EN_EX_PVE_FIX) begin
        always_comb pve_0_init_lt_axi_s_aruser = i_pve_0_init_lt_axi_s_arid[6:4];
        always_comb pve_0_init_lt_axi_s_awuser = i_pve_0_init_lt_axi_s_awid[6:4];
        always_comb pve_1_init_lt_axi_s_aruser = i_pve_1_init_lt_axi_s_arid[6:4];
        always_comb pve_1_init_lt_axi_s_awuser = i_pve_1_init_lt_axi_s_awid[6:4];
    // ----------
    end else begin
        assign pve_0_init_lt_axi_s_aruser = 3'b000;
        assign pve_0_init_lt_axi_s_awuser = 3'b000;
        assign pve_1_init_lt_axi_s_aruser = 3'b000;
        assign pve_1_init_lt_axi_s_awuser = 3'b000;
    end

    // Automated Address MSB fix: extra nets declaration
    logic[40:0] apu_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] apu_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] apu_init_mt_axi_s_araddr_msb_fixed;
    logic[40:0] apu_init_mt_axi_s_awaddr_msb_fixed;
    logic[40:0] apu_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] apu_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] dcd_dec_0_init_mt_axi_s_araddr_msb_fixed;
    logic[40:0] dcd_dec_0_init_mt_axi_s_awaddr_msb_fixed;
    logic[40:0] dcd_dec_1_init_mt_axi_s_araddr_msb_fixed;
    logic[40:0] dcd_dec_1_init_mt_axi_s_awaddr_msb_fixed;
    logic[40:0] dcd_dec_2_init_mt_axi_s_araddr_msb_fixed;
    logic[40:0] dcd_dec_2_init_mt_axi_s_awaddr_msb_fixed;
    logic[40:0] dcd_mcu_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] dcd_mcu_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] pcie_init_mt_axi_s_araddr_msb_fixed;
    logic[40:0] pcie_init_mt_axi_s_awaddr_msb_fixed;
    logic[40:0] pcie_targ_cfg_dbi_axi_m_araddr_msb_fixed;
    logic[40:0] pcie_targ_cfg_dbi_axi_m_awaddr_msb_fixed;
    logic[40:0] pcie_targ_mt_axi_m_araddr_msb_fixed;
    logic[40:0] pcie_targ_mt_axi_m_awaddr_msb_fixed;
    logic[40:0] pve_0_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] pve_0_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] pve_0_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] pve_0_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] pve_0_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] pve_0_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] pve_1_init_ht_axi_s_araddr_msb_fixed;
    logic[40:0] pve_1_init_ht_axi_s_awaddr_msb_fixed;
    logic[40:0] pve_1_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] pve_1_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] pve_1_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] pve_1_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] soc_mgmt_init_lt_axi_s_araddr_msb_fixed;
    logic[40:0] soc_mgmt_init_lt_axi_s_awaddr_msb_fixed;
    logic[40:0] soc_mgmt_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] soc_mgmt_targ_lt_axi_m_awaddr_msb_fixed;
    logic[40:0] sys_spm_targ_lt_axi_m_araddr_msb_fixed;
    logic[40:0] sys_spm_targ_lt_axi_m_awaddr_msb_fixed;

    // Automated Address MSB fix: Initiator-side assignments to extend addresses by 1 bit
    noc_common_addr_msb_setter u_addr_msb_fix_apu_init_lt (
        .i_axi_araddr_40b (i_apu_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (apu_init_lt_axi_s_araddr_msb_fixed)
    );
    assign apu_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_apu_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_apu_init_mt (
        .i_axi_araddr_40b (i_apu_init_mt_axi_s_araddr),
        .o_axi_araddr_41b (apu_init_mt_axi_s_araddr_msb_fixed)
    );
    assign apu_init_mt_axi_s_awaddr_msb_fixed = {1'b0, i_apu_init_mt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_dcd_dec_0_init_mt (
        .i_axi_araddr_40b (i_dcd_dec_0_init_mt_axi_s_araddr),
        .o_axi_araddr_41b (dcd_dec_0_init_mt_axi_s_araddr_msb_fixed)
    );
    assign dcd_dec_0_init_mt_axi_s_awaddr_msb_fixed = {1'b0, i_dcd_dec_0_init_mt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_dcd_dec_1_init_mt (
        .i_axi_araddr_40b (i_dcd_dec_1_init_mt_axi_s_araddr),
        .o_axi_araddr_41b (dcd_dec_1_init_mt_axi_s_araddr_msb_fixed)
    );
    assign dcd_dec_1_init_mt_axi_s_awaddr_msb_fixed = {1'b0, i_dcd_dec_1_init_mt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_dcd_dec_2_init_mt (
        .i_axi_araddr_40b (i_dcd_dec_2_init_mt_axi_s_araddr),
        .o_axi_araddr_41b (dcd_dec_2_init_mt_axi_s_araddr_msb_fixed)
    );
    assign dcd_dec_2_init_mt_axi_s_awaddr_msb_fixed = {1'b0, i_dcd_dec_2_init_mt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_dcd_mcu_init_lt (
        .i_axi_araddr_40b (i_dcd_mcu_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (dcd_mcu_init_lt_axi_s_araddr_msb_fixed)
    );
    assign dcd_mcu_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_dcd_mcu_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_pcie_init_mt (
        .i_axi_araddr_40b (i_pcie_init_mt_axi_s_araddr),
        .o_axi_araddr_41b (pcie_init_mt_axi_s_araddr_msb_fixed)
    );
    assign pcie_init_mt_axi_s_awaddr_msb_fixed = {1'b0, i_pcie_init_mt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_pve_0_init_ht (
        .i_axi_araddr_40b (i_pve_0_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (pve_0_init_ht_axi_s_araddr_msb_fixed)
    );
    assign pve_0_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_pve_0_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_pve_0_init_lt (
        .i_axi_araddr_40b (i_pve_0_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (pve_0_init_lt_axi_s_araddr_msb_fixed)
    );
    assign pve_0_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_pve_0_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_pve_1_init_ht (
        .i_axi_araddr_40b (i_pve_1_init_ht_axi_s_araddr),
        .o_axi_araddr_41b (pve_1_init_ht_axi_s_araddr_msb_fixed)
    );
    assign pve_1_init_ht_axi_s_awaddr_msb_fixed = {1'b0, i_pve_1_init_ht_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_pve_1_init_lt (
        .i_axi_araddr_40b (i_pve_1_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (pve_1_init_lt_axi_s_araddr_msb_fixed)
    );
    assign pve_1_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_pve_1_init_lt_axi_s_awaddr};
    noc_common_addr_msb_setter u_addr_msb_fix_soc_mgmt_init_lt (
        .i_axi_araddr_40b (i_soc_mgmt_init_lt_axi_s_araddr),
        .o_axi_araddr_41b (soc_mgmt_init_lt_axi_s_araddr_msb_fixed)
    );
    assign soc_mgmt_init_lt_axi_s_awaddr_msb_fixed = {1'b0, i_soc_mgmt_init_lt_axi_s_awaddr};

    // Automated Address MSB fix: Target-side assignments to drop unused MSB
    assign o_apu_targ_lt_axi_m_araddr = apu_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_apu_targ_lt_axi_m_awaddr = apu_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_pcie_targ_cfg_dbi_axi_m_araddr = pcie_targ_cfg_dbi_axi_m_araddr_msb_fixed[39:0];
    assign o_pcie_targ_cfg_dbi_axi_m_awaddr = pcie_targ_cfg_dbi_axi_m_awaddr_msb_fixed[39:0];
    assign o_pcie_targ_mt_axi_m_araddr = pcie_targ_mt_axi_m_araddr_msb_fixed[39:0];
    assign o_pcie_targ_mt_axi_m_awaddr = pcie_targ_mt_axi_m_awaddr_msb_fixed[39:0];
    assign o_pve_0_targ_lt_axi_m_araddr = pve_0_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_pve_0_targ_lt_axi_m_awaddr = pve_0_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_pve_1_targ_lt_axi_m_araddr = pve_1_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_pve_1_targ_lt_axi_m_awaddr = pve_1_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_soc_mgmt_targ_lt_axi_m_araddr = soc_mgmt_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_soc_mgmt_targ_lt_axi_m_awaddr = soc_mgmt_targ_lt_axi_m_awaddr_msb_fixed[39:0];
    assign o_sys_spm_targ_lt_axi_m_araddr = sys_spm_targ_lt_axi_m_araddr_msb_fixed[39:0];
    assign o_sys_spm_targ_lt_axi_m_awaddr = sys_spm_targ_lt_axi_m_awaddr_msb_fixed[39:0];


    noc_art_soc u_noc_art_soc (
    .apu_aon_clk(i_apu_aon_clk),
    .apu_aon_rst_n(i_apu_aon_rst_n),
    .apu_init_lt_Ar_Addr(apu_init_lt_axi_s_araddr_msb_fixed),
    .apu_init_lt_Ar_Burst(i_apu_init_lt_axi_s_arburst),
    .apu_init_lt_Ar_Cache(i_apu_init_lt_axi_s_arcache),
    .apu_init_lt_Ar_Id(i_apu_init_lt_axi_s_arid),
    .apu_init_lt_Ar_Len(i_apu_init_lt_axi_s_arlen),
    .apu_init_lt_Ar_Lock(i_apu_init_lt_axi_s_arlock),
    .apu_init_lt_Ar_Prot(i_apu_init_lt_axi_s_arprot),
    .apu_init_lt_Ar_Qos(i_apu_init_lt_axi_s_arqos),
    .apu_init_lt_Ar_Ready(o_apu_init_lt_axi_s_arready),
    .apu_init_lt_Ar_Size(i_apu_init_lt_axi_s_arsize),
    .apu_init_lt_Ar_User(apu_init_lt_axi_s_aruser),
    .apu_init_lt_Ar_Valid(i_apu_init_lt_axi_s_arvalid),
    .apu_init_lt_Aw_Addr(apu_init_lt_axi_s_awaddr_msb_fixed),
    .apu_init_lt_Aw_Burst(i_apu_init_lt_axi_s_awburst),
    .apu_init_lt_Aw_Cache(i_apu_init_lt_axi_s_awcache),
    .apu_init_lt_Aw_Id(i_apu_init_lt_axi_s_awid),
    .apu_init_lt_Aw_Len(i_apu_init_lt_axi_s_awlen),
    .apu_init_lt_Aw_Lock(i_apu_init_lt_axi_s_awlock),
    .apu_init_lt_Aw_Prot(i_apu_init_lt_axi_s_awprot),
    .apu_init_lt_Aw_Qos(i_apu_init_lt_axi_s_awqos),
    .apu_init_lt_Aw_Ready(o_apu_init_lt_axi_s_awready),
    .apu_init_lt_Aw_Size(i_apu_init_lt_axi_s_awsize),
    .apu_init_lt_Aw_User(apu_init_lt_axi_s_awuser),
    .apu_init_lt_Aw_Valid(i_apu_init_lt_axi_s_awvalid),
    .apu_init_lt_B_Id(o_apu_init_lt_axi_s_bid),
    .apu_init_lt_B_Ready(i_apu_init_lt_axi_s_bready),
    .apu_init_lt_B_Resp(o_apu_init_lt_axi_s_bresp),
    .apu_init_lt_B_Valid(o_apu_init_lt_axi_s_bvalid),
    .apu_init_lt_R_Data(o_apu_init_lt_axi_s_rdata),
    .apu_init_lt_R_Id(o_apu_init_lt_axi_s_rid),
    .apu_init_lt_R_Last(o_apu_init_lt_axi_s_rlast),
    .apu_init_lt_R_Ready(i_apu_init_lt_axi_s_rready),
    .apu_init_lt_R_Resp(o_apu_init_lt_axi_s_rresp),
    .apu_init_lt_R_Valid(o_apu_init_lt_axi_s_rvalid),
    .apu_init_lt_W_Data(i_apu_init_lt_axi_s_wdata),
    .apu_init_lt_W_Last(i_apu_init_lt_axi_s_wlast),
    .apu_init_lt_W_Ready(o_apu_init_lt_axi_s_wready),
    .apu_init_lt_W_Strb(i_apu_init_lt_axi_s_wstrb),
    .apu_init_lt_W_Valid(i_apu_init_lt_axi_s_wvalid),
    .apu_init_mt_rd_Ar_Addr(apu_init_mt_axi_s_araddr_msb_fixed),
    .apu_init_mt_rd_Ar_Burst(i_apu_init_mt_axi_s_arburst),
    .apu_init_mt_rd_Ar_Cache(i_apu_init_mt_axi_s_arcache),
    .apu_init_mt_rd_Ar_Id(i_apu_init_mt_axi_s_arid),
    .apu_init_mt_rd_Ar_Len(i_apu_init_mt_axi_s_arlen),
    .apu_init_mt_rd_Ar_Lock(i_apu_init_mt_axi_s_arlock),
    .apu_init_mt_rd_Ar_Prot(i_apu_init_mt_axi_s_arprot),
    .apu_init_mt_rd_Ar_Qos(i_apu_init_mt_axi_s_arqos),
    .apu_init_mt_rd_Ar_Ready(o_apu_init_mt_axi_s_arready),
    .apu_init_mt_rd_Ar_Size(i_apu_init_mt_axi_s_arsize),
    .apu_init_mt_rd_Ar_Valid(i_apu_init_mt_axi_s_arvalid),
    .apu_init_mt_rd_R_Data(o_apu_init_mt_axi_s_rdata),
    .apu_init_mt_rd_R_Id(o_apu_init_mt_axi_s_rid),
    .apu_init_mt_rd_R_Last(o_apu_init_mt_axi_s_rlast),
    .apu_init_mt_rd_R_Ready(i_apu_init_mt_axi_s_rready),
    .apu_init_mt_rd_R_Resp(o_apu_init_mt_axi_s_rresp),
    .apu_init_mt_rd_R_Valid(o_apu_init_mt_axi_s_rvalid),
    .apu_init_mt_wr_Aw_Addr(apu_init_mt_axi_s_awaddr_msb_fixed),
    .apu_init_mt_wr_Aw_Burst(i_apu_init_mt_axi_s_awburst),
    .apu_init_mt_wr_Aw_Cache(i_apu_init_mt_axi_s_awcache),
    .apu_init_mt_wr_Aw_Id(i_apu_init_mt_axi_s_awid),
    .apu_init_mt_wr_Aw_Len(i_apu_init_mt_axi_s_awlen),
    .apu_init_mt_wr_Aw_Lock(i_apu_init_mt_axi_s_awlock),
    .apu_init_mt_wr_Aw_Prot(i_apu_init_mt_axi_s_awprot),
    .apu_init_mt_wr_Aw_Qos(i_apu_init_mt_axi_s_awqos),
    .apu_init_mt_wr_Aw_Ready(o_apu_init_mt_axi_s_awready),
    .apu_init_mt_wr_Aw_Size(i_apu_init_mt_axi_s_awsize),
    .apu_init_mt_wr_Aw_Valid(i_apu_init_mt_axi_s_awvalid),
    .apu_init_mt_wr_B_Id(o_apu_init_mt_axi_s_bid),
    .apu_init_mt_wr_B_Ready(i_apu_init_mt_axi_s_bready),
    .apu_init_mt_wr_B_Resp(o_apu_init_mt_axi_s_bresp),
    .apu_init_mt_wr_B_Valid(o_apu_init_mt_axi_s_bvalid),
    .apu_init_mt_wr_W_Data(i_apu_init_mt_axi_s_wdata),
    .apu_init_mt_wr_W_Last(i_apu_init_mt_axi_s_wlast),
    .apu_init_mt_wr_W_Ready(o_apu_init_mt_axi_s_wready),
    .apu_init_mt_wr_W_Strb(i_apu_init_mt_axi_s_wstrb),
    .apu_init_mt_wr_W_Valid(i_apu_init_mt_axi_s_wvalid),
    .apu_pwr_Idle(o_apu_pwr_idle_val),
    .apu_pwr_IdleAck(o_apu_pwr_idle_ack),
    .apu_pwr_IdleReq(i_apu_pwr_idle_req),
    .apu_targ_lt_Ar_Addr(apu_targ_lt_axi_m_araddr_msb_fixed),
    .apu_targ_lt_Ar_Burst(o_apu_targ_lt_axi_m_arburst),
    .apu_targ_lt_Ar_Cache(o_apu_targ_lt_axi_m_arcache),
    .apu_targ_lt_Ar_Id(o_apu_targ_lt_axi_m_arid),
    .apu_targ_lt_Ar_Len(o_apu_targ_lt_axi_m_arlen),
    .apu_targ_lt_Ar_Lock(o_apu_targ_lt_axi_m_arlock),
    .apu_targ_lt_Ar_Prot(o_apu_targ_lt_axi_m_arprot),
    .apu_targ_lt_Ar_Qos(o_apu_targ_lt_axi_m_arqos),
    .apu_targ_lt_Ar_Ready(i_apu_targ_lt_axi_m_arready),
    .apu_targ_lt_Ar_Size(o_apu_targ_lt_axi_m_arsize),
    .apu_targ_lt_Ar_Valid(o_apu_targ_lt_axi_m_arvalid),
    .apu_targ_lt_Aw_Addr(apu_targ_lt_axi_m_awaddr_msb_fixed),
    .apu_targ_lt_Aw_Burst(o_apu_targ_lt_axi_m_awburst),
    .apu_targ_lt_Aw_Cache(o_apu_targ_lt_axi_m_awcache),
    .apu_targ_lt_Aw_Id(o_apu_targ_lt_axi_m_awid),
    .apu_targ_lt_Aw_Len(o_apu_targ_lt_axi_m_awlen),
    .apu_targ_lt_Aw_Lock(o_apu_targ_lt_axi_m_awlock),
    .apu_targ_lt_Aw_Prot(o_apu_targ_lt_axi_m_awprot),
    .apu_targ_lt_Aw_Qos(o_apu_targ_lt_axi_m_awqos),
    .apu_targ_lt_Aw_Ready(i_apu_targ_lt_axi_m_awready),
    .apu_targ_lt_Aw_Size(o_apu_targ_lt_axi_m_awsize),
    .apu_targ_lt_Aw_Valid(o_apu_targ_lt_axi_m_awvalid),
    .apu_targ_lt_B_Id(i_apu_targ_lt_axi_m_bid),
    .apu_targ_lt_B_Ready(o_apu_targ_lt_axi_m_bready),
    .apu_targ_lt_B_Resp(i_apu_targ_lt_axi_m_bresp),
    .apu_targ_lt_B_Valid(i_apu_targ_lt_axi_m_bvalid),
    .apu_targ_lt_R_Data(i_apu_targ_lt_axi_m_rdata),
    .apu_targ_lt_R_Id(i_apu_targ_lt_axi_m_rid),
    .apu_targ_lt_R_Last(i_apu_targ_lt_axi_m_rlast),
    .apu_targ_lt_R_Ready(o_apu_targ_lt_axi_m_rready),
    .apu_targ_lt_R_Resp(i_apu_targ_lt_axi_m_rresp),
    .apu_targ_lt_R_Valid(i_apu_targ_lt_axi_m_rvalid),
    .apu_targ_lt_W_Data(o_apu_targ_lt_axi_m_wdata),
    .apu_targ_lt_W_Last(o_apu_targ_lt_axi_m_wlast),
    .apu_targ_lt_W_Ready(i_apu_targ_lt_axi_m_wready),
    .apu_targ_lt_W_Strb(o_apu_targ_lt_axi_m_wstrb),
    .apu_targ_lt_W_Valid(o_apu_targ_lt_axi_m_wvalid),
    .apu_targ_syscfg_PAddr(o_apu_targ_syscfg_apb_m_paddr),
    .apu_targ_syscfg_PEnable(o_apu_targ_syscfg_apb_m_penable),
    .apu_targ_syscfg_PProt(o_apu_targ_syscfg_apb_m_pprot),
    .apu_targ_syscfg_PRData(i_apu_targ_syscfg_apb_m_prdata),
    .apu_targ_syscfg_PReady(i_apu_targ_syscfg_apb_m_pready),
    .apu_targ_syscfg_PSel(o_apu_targ_syscfg_apb_m_psel),
    .apu_targ_syscfg_PSlvErr(i_apu_targ_syscfg_apb_m_pslverr),
    .apu_targ_syscfg_PStrb(o_apu_targ_syscfg_apb_m_pstrb),
    .apu_targ_syscfg_PWData(o_apu_targ_syscfg_apb_m_pwdata),
    .apu_targ_syscfg_PWrite(o_apu_targ_syscfg_apb_m_pwrite),
    .apu_x_clk(i_apu_x_clk),
    .apu_x_clken(i_apu_x_clken),
    .apu_x_rst_n(i_apu_x_rst_n),
    .dcd_aon_clk(i_dcd_aon_clk),
    .dcd_aon_rst_n(i_dcd_aon_rst_n),
    .dcd_codec_clk(i_dcd_codec_clk),
    .dcd_codec_clken(i_dcd_codec_clken),
    .dcd_codec_rst_n(i_dcd_codec_rst_n),
    .dcd_dec_0_init_mt_rd_Ar_Addr(dcd_dec_0_init_mt_axi_s_araddr_msb_fixed),
    .dcd_dec_0_init_mt_rd_Ar_Burst(i_dcd_dec_0_init_mt_axi_s_arburst),
    .dcd_dec_0_init_mt_rd_Ar_Cache(i_dcd_dec_0_init_mt_axi_s_arcache),
    .dcd_dec_0_init_mt_rd_Ar_Id(i_dcd_dec_0_init_mt_axi_s_arid),
    .dcd_dec_0_init_mt_rd_Ar_Len(i_dcd_dec_0_init_mt_axi_s_arlen),
    .dcd_dec_0_init_mt_rd_Ar_Lock(i_dcd_dec_0_init_mt_axi_s_arlock),
    .dcd_dec_0_init_mt_rd_Ar_Prot(i_dcd_dec_0_init_mt_axi_s_arprot),
    .dcd_dec_0_init_mt_rd_Ar_Qos(i_dcd_dec_0_init_mt_axi_s_arqos),
    .dcd_dec_0_init_mt_rd_Ar_Ready(o_dcd_dec_0_init_mt_axi_s_arready),
    .dcd_dec_0_init_mt_rd_Ar_Size(i_dcd_dec_0_init_mt_axi_s_arsize),
    .dcd_dec_0_init_mt_rd_Ar_Valid(i_dcd_dec_0_init_mt_axi_s_arvalid),
    .dcd_dec_0_init_mt_rd_R_Data(o_dcd_dec_0_init_mt_axi_s_rdata),
    .dcd_dec_0_init_mt_rd_R_Id(o_dcd_dec_0_init_mt_axi_s_rid),
    .dcd_dec_0_init_mt_rd_R_Last(o_dcd_dec_0_init_mt_axi_s_rlast),
    .dcd_dec_0_init_mt_rd_R_Ready(i_dcd_dec_0_init_mt_axi_s_rready),
    .dcd_dec_0_init_mt_rd_R_Resp(o_dcd_dec_0_init_mt_axi_s_rresp),
    .dcd_dec_0_init_mt_rd_R_Valid(o_dcd_dec_0_init_mt_axi_s_rvalid),
    .dcd_dec_0_init_mt_wr_Aw_Addr(dcd_dec_0_init_mt_axi_s_awaddr_msb_fixed),
    .dcd_dec_0_init_mt_wr_Aw_Burst(i_dcd_dec_0_init_mt_axi_s_awburst),
    .dcd_dec_0_init_mt_wr_Aw_Cache(i_dcd_dec_0_init_mt_axi_s_awcache),
    .dcd_dec_0_init_mt_wr_Aw_Id(i_dcd_dec_0_init_mt_axi_s_awid),
    .dcd_dec_0_init_mt_wr_Aw_Len(i_dcd_dec_0_init_mt_axi_s_awlen),
    .dcd_dec_0_init_mt_wr_Aw_Lock(i_dcd_dec_0_init_mt_axi_s_awlock),
    .dcd_dec_0_init_mt_wr_Aw_Prot(i_dcd_dec_0_init_mt_axi_s_awprot),
    .dcd_dec_0_init_mt_wr_Aw_Qos(i_dcd_dec_0_init_mt_axi_s_awqos),
    .dcd_dec_0_init_mt_wr_Aw_Ready(o_dcd_dec_0_init_mt_axi_s_awready),
    .dcd_dec_0_init_mt_wr_Aw_Size(i_dcd_dec_0_init_mt_axi_s_awsize),
    .dcd_dec_0_init_mt_wr_Aw_Valid(i_dcd_dec_0_init_mt_axi_s_awvalid),
    .dcd_dec_0_init_mt_wr_B_Id(o_dcd_dec_0_init_mt_axi_s_bid),
    .dcd_dec_0_init_mt_wr_B_Ready(i_dcd_dec_0_init_mt_axi_s_bready),
    .dcd_dec_0_init_mt_wr_B_Resp(o_dcd_dec_0_init_mt_axi_s_bresp),
    .dcd_dec_0_init_mt_wr_B_Valid(o_dcd_dec_0_init_mt_axi_s_bvalid),
    .dcd_dec_0_init_mt_wr_W_Data(i_dcd_dec_0_init_mt_axi_s_wdata),
    .dcd_dec_0_init_mt_wr_W_Last(i_dcd_dec_0_init_mt_axi_s_wlast),
    .dcd_dec_0_init_mt_wr_W_Ready(o_dcd_dec_0_init_mt_axi_s_wready),
    .dcd_dec_0_init_mt_wr_W_Strb(i_dcd_dec_0_init_mt_axi_s_wstrb),
    .dcd_dec_0_init_mt_wr_W_Valid(i_dcd_dec_0_init_mt_axi_s_wvalid),
    .dcd_dec_1_init_mt_rd_Ar_Addr(dcd_dec_1_init_mt_axi_s_araddr_msb_fixed),
    .dcd_dec_1_init_mt_rd_Ar_Burst(i_dcd_dec_1_init_mt_axi_s_arburst),
    .dcd_dec_1_init_mt_rd_Ar_Cache(i_dcd_dec_1_init_mt_axi_s_arcache),
    .dcd_dec_1_init_mt_rd_Ar_Id(i_dcd_dec_1_init_mt_axi_s_arid),
    .dcd_dec_1_init_mt_rd_Ar_Len(i_dcd_dec_1_init_mt_axi_s_arlen),
    .dcd_dec_1_init_mt_rd_Ar_Lock(i_dcd_dec_1_init_mt_axi_s_arlock),
    .dcd_dec_1_init_mt_rd_Ar_Prot(i_dcd_dec_1_init_mt_axi_s_arprot),
    .dcd_dec_1_init_mt_rd_Ar_Qos(i_dcd_dec_1_init_mt_axi_s_arqos),
    .dcd_dec_1_init_mt_rd_Ar_Ready(o_dcd_dec_1_init_mt_axi_s_arready),
    .dcd_dec_1_init_mt_rd_Ar_Size(i_dcd_dec_1_init_mt_axi_s_arsize),
    .dcd_dec_1_init_mt_rd_Ar_Valid(i_dcd_dec_1_init_mt_axi_s_arvalid),
    .dcd_dec_1_init_mt_rd_R_Data(o_dcd_dec_1_init_mt_axi_s_rdata),
    .dcd_dec_1_init_mt_rd_R_Id(o_dcd_dec_1_init_mt_axi_s_rid),
    .dcd_dec_1_init_mt_rd_R_Last(o_dcd_dec_1_init_mt_axi_s_rlast),
    .dcd_dec_1_init_mt_rd_R_Ready(i_dcd_dec_1_init_mt_axi_s_rready),
    .dcd_dec_1_init_mt_rd_R_Resp(o_dcd_dec_1_init_mt_axi_s_rresp),
    .dcd_dec_1_init_mt_rd_R_Valid(o_dcd_dec_1_init_mt_axi_s_rvalid),
    .dcd_dec_1_init_mt_wr_Aw_Addr(dcd_dec_1_init_mt_axi_s_awaddr_msb_fixed),
    .dcd_dec_1_init_mt_wr_Aw_Burst(i_dcd_dec_1_init_mt_axi_s_awburst),
    .dcd_dec_1_init_mt_wr_Aw_Cache(i_dcd_dec_1_init_mt_axi_s_awcache),
    .dcd_dec_1_init_mt_wr_Aw_Id(i_dcd_dec_1_init_mt_axi_s_awid),
    .dcd_dec_1_init_mt_wr_Aw_Len(i_dcd_dec_1_init_mt_axi_s_awlen),
    .dcd_dec_1_init_mt_wr_Aw_Lock(i_dcd_dec_1_init_mt_axi_s_awlock),
    .dcd_dec_1_init_mt_wr_Aw_Prot(i_dcd_dec_1_init_mt_axi_s_awprot),
    .dcd_dec_1_init_mt_wr_Aw_Qos(i_dcd_dec_1_init_mt_axi_s_awqos),
    .dcd_dec_1_init_mt_wr_Aw_Ready(o_dcd_dec_1_init_mt_axi_s_awready),
    .dcd_dec_1_init_mt_wr_Aw_Size(i_dcd_dec_1_init_mt_axi_s_awsize),
    .dcd_dec_1_init_mt_wr_Aw_Valid(i_dcd_dec_1_init_mt_axi_s_awvalid),
    .dcd_dec_1_init_mt_wr_B_Id(o_dcd_dec_1_init_mt_axi_s_bid),
    .dcd_dec_1_init_mt_wr_B_Ready(i_dcd_dec_1_init_mt_axi_s_bready),
    .dcd_dec_1_init_mt_wr_B_Resp(o_dcd_dec_1_init_mt_axi_s_bresp),
    .dcd_dec_1_init_mt_wr_B_Valid(o_dcd_dec_1_init_mt_axi_s_bvalid),
    .dcd_dec_1_init_mt_wr_W_Data(i_dcd_dec_1_init_mt_axi_s_wdata),
    .dcd_dec_1_init_mt_wr_W_Last(i_dcd_dec_1_init_mt_axi_s_wlast),
    .dcd_dec_1_init_mt_wr_W_Ready(o_dcd_dec_1_init_mt_axi_s_wready),
    .dcd_dec_1_init_mt_wr_W_Strb(i_dcd_dec_1_init_mt_axi_s_wstrb),
    .dcd_dec_1_init_mt_wr_W_Valid(i_dcd_dec_1_init_mt_axi_s_wvalid),
    .dcd_dec_2_init_mt_rd_Ar_Addr(dcd_dec_2_init_mt_axi_s_araddr_msb_fixed),
    .dcd_dec_2_init_mt_rd_Ar_Burst(i_dcd_dec_2_init_mt_axi_s_arburst),
    .dcd_dec_2_init_mt_rd_Ar_Cache(i_dcd_dec_2_init_mt_axi_s_arcache),
    .dcd_dec_2_init_mt_rd_Ar_Id(i_dcd_dec_2_init_mt_axi_s_arid),
    .dcd_dec_2_init_mt_rd_Ar_Len(i_dcd_dec_2_init_mt_axi_s_arlen),
    .dcd_dec_2_init_mt_rd_Ar_Lock(i_dcd_dec_2_init_mt_axi_s_arlock),
    .dcd_dec_2_init_mt_rd_Ar_Prot(i_dcd_dec_2_init_mt_axi_s_arprot),
    .dcd_dec_2_init_mt_rd_Ar_Qos(i_dcd_dec_2_init_mt_axi_s_arqos),
    .dcd_dec_2_init_mt_rd_Ar_Ready(o_dcd_dec_2_init_mt_axi_s_arready),
    .dcd_dec_2_init_mt_rd_Ar_Size(i_dcd_dec_2_init_mt_axi_s_arsize),
    .dcd_dec_2_init_mt_rd_Ar_Valid(i_dcd_dec_2_init_mt_axi_s_arvalid),
    .dcd_dec_2_init_mt_rd_R_Data(o_dcd_dec_2_init_mt_axi_s_rdata),
    .dcd_dec_2_init_mt_rd_R_Id(o_dcd_dec_2_init_mt_axi_s_rid),
    .dcd_dec_2_init_mt_rd_R_Last(o_dcd_dec_2_init_mt_axi_s_rlast),
    .dcd_dec_2_init_mt_rd_R_Ready(i_dcd_dec_2_init_mt_axi_s_rready),
    .dcd_dec_2_init_mt_rd_R_Resp(o_dcd_dec_2_init_mt_axi_s_rresp),
    .dcd_dec_2_init_mt_rd_R_Valid(o_dcd_dec_2_init_mt_axi_s_rvalid),
    .dcd_dec_2_init_mt_wr_Aw_Addr(dcd_dec_2_init_mt_axi_s_awaddr_msb_fixed),
    .dcd_dec_2_init_mt_wr_Aw_Burst(i_dcd_dec_2_init_mt_axi_s_awburst),
    .dcd_dec_2_init_mt_wr_Aw_Cache(i_dcd_dec_2_init_mt_axi_s_awcache),
    .dcd_dec_2_init_mt_wr_Aw_Id(i_dcd_dec_2_init_mt_axi_s_awid),
    .dcd_dec_2_init_mt_wr_Aw_Len(i_dcd_dec_2_init_mt_axi_s_awlen),
    .dcd_dec_2_init_mt_wr_Aw_Lock(i_dcd_dec_2_init_mt_axi_s_awlock),
    .dcd_dec_2_init_mt_wr_Aw_Prot(i_dcd_dec_2_init_mt_axi_s_awprot),
    .dcd_dec_2_init_mt_wr_Aw_Qos(i_dcd_dec_2_init_mt_axi_s_awqos),
    .dcd_dec_2_init_mt_wr_Aw_Ready(o_dcd_dec_2_init_mt_axi_s_awready),
    .dcd_dec_2_init_mt_wr_Aw_Size(i_dcd_dec_2_init_mt_axi_s_awsize),
    .dcd_dec_2_init_mt_wr_Aw_Valid(i_dcd_dec_2_init_mt_axi_s_awvalid),
    .dcd_dec_2_init_mt_wr_B_Id(o_dcd_dec_2_init_mt_axi_s_bid),
    .dcd_dec_2_init_mt_wr_B_Ready(i_dcd_dec_2_init_mt_axi_s_bready),
    .dcd_dec_2_init_mt_wr_B_Resp(o_dcd_dec_2_init_mt_axi_s_bresp),
    .dcd_dec_2_init_mt_wr_B_Valid(o_dcd_dec_2_init_mt_axi_s_bvalid),
    .dcd_dec_2_init_mt_wr_W_Data(i_dcd_dec_2_init_mt_axi_s_wdata),
    .dcd_dec_2_init_mt_wr_W_Last(i_dcd_dec_2_init_mt_axi_s_wlast),
    .dcd_dec_2_init_mt_wr_W_Ready(o_dcd_dec_2_init_mt_axi_s_wready),
    .dcd_dec_2_init_mt_wr_W_Strb(i_dcd_dec_2_init_mt_axi_s_wstrb),
    .dcd_dec_2_init_mt_wr_W_Valid(i_dcd_dec_2_init_mt_axi_s_wvalid),
    .dcd_mcu_clk(i_dcd_mcu_clk),
    .dcd_mcu_clken(i_dcd_mcu_clken),
    .dcd_mcu_init_lt_rd_Ar_Addr(dcd_mcu_init_lt_axi_s_araddr_msb_fixed),
    .dcd_mcu_init_lt_rd_Ar_Burst(i_dcd_mcu_init_lt_axi_s_arburst),
    .dcd_mcu_init_lt_rd_Ar_Cache(i_dcd_mcu_init_lt_axi_s_arcache),
    .dcd_mcu_init_lt_rd_Ar_Id(i_dcd_mcu_init_lt_axi_s_arid),
    .dcd_mcu_init_lt_rd_Ar_Len(i_dcd_mcu_init_lt_axi_s_arlen),
    .dcd_mcu_init_lt_rd_Ar_Lock(i_dcd_mcu_init_lt_axi_s_arlock),
    .dcd_mcu_init_lt_rd_Ar_Prot(i_dcd_mcu_init_lt_axi_s_arprot),
    .dcd_mcu_init_lt_rd_Ar_Qos(i_dcd_mcu_init_lt_axi_s_arqos),
    .dcd_mcu_init_lt_rd_Ar_Ready(o_dcd_mcu_init_lt_axi_s_arready),
    .dcd_mcu_init_lt_rd_Ar_Size(i_dcd_mcu_init_lt_axi_s_arsize),
    .dcd_mcu_init_lt_rd_Ar_Valid(i_dcd_mcu_init_lt_axi_s_arvalid),
    .dcd_mcu_init_lt_rd_R_Data(o_dcd_mcu_init_lt_axi_s_rdata),
    .dcd_mcu_init_lt_rd_R_Id(o_dcd_mcu_init_lt_axi_s_rid),
    .dcd_mcu_init_lt_rd_R_Last(o_dcd_mcu_init_lt_axi_s_rlast),
    .dcd_mcu_init_lt_rd_R_Ready(i_dcd_mcu_init_lt_axi_s_rready),
    .dcd_mcu_init_lt_rd_R_Resp(o_dcd_mcu_init_lt_axi_s_rresp),
    .dcd_mcu_init_lt_rd_R_Valid(o_dcd_mcu_init_lt_axi_s_rvalid),
    .dcd_mcu_init_lt_wr_Aw_Addr(dcd_mcu_init_lt_axi_s_awaddr_msb_fixed),
    .dcd_mcu_init_lt_wr_Aw_Burst(i_dcd_mcu_init_lt_axi_s_awburst),
    .dcd_mcu_init_lt_wr_Aw_Cache(i_dcd_mcu_init_lt_axi_s_awcache),
    .dcd_mcu_init_lt_wr_Aw_Id(i_dcd_mcu_init_lt_axi_s_awid),
    .dcd_mcu_init_lt_wr_Aw_Len(i_dcd_mcu_init_lt_axi_s_awlen),
    .dcd_mcu_init_lt_wr_Aw_Lock(i_dcd_mcu_init_lt_axi_s_awlock),
    .dcd_mcu_init_lt_wr_Aw_Prot(i_dcd_mcu_init_lt_axi_s_awprot),
    .dcd_mcu_init_lt_wr_Aw_Qos(i_dcd_mcu_init_lt_axi_s_awqos),
    .dcd_mcu_init_lt_wr_Aw_Ready(o_dcd_mcu_init_lt_axi_s_awready),
    .dcd_mcu_init_lt_wr_Aw_Size(i_dcd_mcu_init_lt_axi_s_awsize),
    .dcd_mcu_init_lt_wr_Aw_Valid(i_dcd_mcu_init_lt_axi_s_awvalid),
    .dcd_mcu_init_lt_wr_B_Id(o_dcd_mcu_init_lt_axi_s_bid),
    .dcd_mcu_init_lt_wr_B_Ready(i_dcd_mcu_init_lt_axi_s_bready),
    .dcd_mcu_init_lt_wr_B_Resp(o_dcd_mcu_init_lt_axi_s_bresp),
    .dcd_mcu_init_lt_wr_B_Valid(o_dcd_mcu_init_lt_axi_s_bvalid),
    .dcd_mcu_init_lt_wr_W_Data(i_dcd_mcu_init_lt_axi_s_wdata),
    .dcd_mcu_init_lt_wr_W_Last(i_dcd_mcu_init_lt_axi_s_wlast),
    .dcd_mcu_init_lt_wr_W_Ready(o_dcd_mcu_init_lt_axi_s_wready),
    .dcd_mcu_init_lt_wr_W_Strb(i_dcd_mcu_init_lt_axi_s_wstrb),
    .dcd_mcu_init_lt_wr_W_Valid(i_dcd_mcu_init_lt_axi_s_wvalid),
    .dcd_mcu_pwr_Idle(o_dcd_mcu_pwr_idle_val),
    .dcd_mcu_pwr_IdleAck(o_dcd_mcu_pwr_idle_ack),
    .dcd_mcu_pwr_IdleReq(i_dcd_mcu_pwr_idle_req),
    .dcd_mcu_rst_n(i_dcd_mcu_rst_n),
    .dcd_pwr_Idle(o_dcd_pwr_idle_val),
    .dcd_pwr_IdleAck(o_dcd_pwr_idle_ack),
    .dcd_pwr_IdleReq(i_dcd_pwr_idle_req),
    .dcd_targ_cfg_PAddr(o_dcd_targ_cfg_apb_m_paddr),
    .dcd_targ_cfg_PEnable(o_dcd_targ_cfg_apb_m_penable),
    .dcd_targ_cfg_PProt(o_dcd_targ_cfg_apb_m_pprot),
    .dcd_targ_cfg_PRData(i_dcd_targ_cfg_apb_m_prdata),
    .dcd_targ_cfg_PReady(i_dcd_targ_cfg_apb_m_pready),
    .dcd_targ_cfg_PSel(o_dcd_targ_cfg_apb_m_psel),
    .dcd_targ_cfg_PSlvErr(i_dcd_targ_cfg_apb_m_pslverr),
    .dcd_targ_cfg_PStrb(o_dcd_targ_cfg_apb_m_pstrb),
    .dcd_targ_cfg_PWData(o_dcd_targ_cfg_apb_m_pwdata),
    .dcd_targ_cfg_PWrite(o_dcd_targ_cfg_apb_m_pwrite),
    .dcd_targ_syscfg_PAddr(o_dcd_targ_syscfg_apb_m_paddr),
    .dcd_targ_syscfg_PEnable(o_dcd_targ_syscfg_apb_m_penable),
    .dcd_targ_syscfg_PProt(o_dcd_targ_syscfg_apb_m_pprot),
    .dcd_targ_syscfg_PRData(i_dcd_targ_syscfg_apb_m_prdata),
    .dcd_targ_syscfg_PReady(i_dcd_targ_syscfg_apb_m_pready),
    .dcd_targ_syscfg_PSel(o_dcd_targ_syscfg_apb_m_psel),
    .dcd_targ_syscfg_PSlvErr(i_dcd_targ_syscfg_apb_m_pslverr),
    .dcd_targ_syscfg_PStrb(o_dcd_targ_syscfg_apb_m_pstrb),
    .dcd_targ_syscfg_PWData(o_dcd_targ_syscfg_apb_m_pwdata),
    .dcd_targ_syscfg_PWrite(o_dcd_targ_syscfg_apb_m_pwrite),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Data(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Head(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Rdy(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Tail(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_Vld(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Data(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Head(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Rdy(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Tail(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_Vld(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Data(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Head(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Rdy(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Tail(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail),
    .dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_Vld(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Data(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Head(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Rdy(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Tail(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail),
    .dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_Vld(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Data(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Head(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Rdy(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Tail(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail),
    .dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_Vld(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Data(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Head(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Rdy(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Tail(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail),
    .dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_Vld(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Data(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Head(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Rdy(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Tail(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail),
    .dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_Vld(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Data(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Head(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Rdy(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Tail(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail),
    .dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_Vld(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Data(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Head(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Rdy(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Tail(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail),
    .dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_Vld(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Data(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Head(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Rdy(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Tail(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail),
    .dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_Vld(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Data(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Head(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Rdy(o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Tail(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail),
    .dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_Vld(i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Data(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Head(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Rdy(i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Tail(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail),
    .dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_Vld(o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Data(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Head(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Rdy(i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Tail(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_Vld(o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Data(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Head(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Rdy(o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Tail(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_Vld(i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Data(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Head(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Rdy(i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Tail(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_Vld(o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Data(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Head(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Rdy(o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Tail(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_Vld(i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Data(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Head(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Rdy(i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Tail(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_Vld(o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Data(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Head(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Rdy(o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Tail(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_Vld(i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Data(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Head(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Rdy(i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Tail(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_Vld(o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Data(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Head(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Rdy(o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Tail(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_Vld(i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Data(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Head(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Rdy(i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Tail(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail),
    .dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_Vld(o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Data(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Head(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Rdy(o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Tail(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_Vld(i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Data(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Head(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Rdy(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Tail(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail),
    .dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_Vld(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Data(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Head(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Rdy(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Tail(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail),
    .dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_Vld(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Data(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Head(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Rdy(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Tail(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail),
    .dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_Vld(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Data(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Head(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Rdy(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Tail(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail),
    .dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_Vld(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Data(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Head(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Rdy(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Tail(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail),
    .dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_Vld(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Data(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Head(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Rdy(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Tail(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail),
    .dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_Vld(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld),
    .l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
    .l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
    .l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
    .l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
    .lnk_buff_dec_128_to_256_ddr_e0_req_mainpde(lnk_buff_dec_128_to_256_ddr_e0_req_mainpde),
    .lnk_buff_dec_128_to_256_ddr_e0_req_mainprn(lnk_buff_dec_128_to_256_ddr_e0_req_mainprn),
    .lnk_buff_dec_128_to_256_ddr_e0_req_mainret(lnk_buff_dec_128_to_256_ddr_e0_req_mainret),
    .lnk_buff_dec_128_to_256_ddr_e0_req_mainse(lnk_buff_dec_128_to_256_ddr_e0_req_mainse),
    .lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainpde(lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainpde),
    .lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainprn(lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainprn),
    .lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainret(lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainret),
    .lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainse(lnk_buff_dec_128_to_256_ddr_e0_req_resp_mainse),
    .lnk_buff_dec_128_to_256_ddr_e1_req_mainpde(lnk_buff_dec_128_to_256_ddr_e1_req_mainpde),
    .lnk_buff_dec_128_to_256_ddr_e1_req_mainprn(lnk_buff_dec_128_to_256_ddr_e1_req_mainprn),
    .lnk_buff_dec_128_to_256_ddr_e1_req_mainret(lnk_buff_dec_128_to_256_ddr_e1_req_mainret),
    .lnk_buff_dec_128_to_256_ddr_e1_req_mainse(lnk_buff_dec_128_to_256_ddr_e1_req_mainse),
    .lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainpde(lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainpde),
    .lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainprn(lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainprn),
    .lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainret(lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainret),
    .lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainse(lnk_buff_dec_128_to_256_ddr_e1_req_resp_mainse),
    .lnk_buff_dec_128_to_256_ddr_e2_req_mainpde(lnk_buff_dec_128_to_256_ddr_e2_req_mainpde),
    .lnk_buff_dec_128_to_256_ddr_e2_req_mainprn(lnk_buff_dec_128_to_256_ddr_e2_req_mainprn),
    .lnk_buff_dec_128_to_256_ddr_e2_req_mainret(lnk_buff_dec_128_to_256_ddr_e2_req_mainret),
    .lnk_buff_dec_128_to_256_ddr_e2_req_mainse(lnk_buff_dec_128_to_256_ddr_e2_req_mainse),
    .lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainpde(lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainpde),
    .lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainprn(lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainprn),
    .lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainret(lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainret),
    .lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainse(lnk_buff_dec_128_to_256_ddr_e2_req_resp_mainse),
    .lnk_buff_dec_128_to_256_ddr_e3_req_mainpde(lnk_buff_dec_128_to_256_ddr_e3_req_mainpde),
    .lnk_buff_dec_128_to_256_ddr_e3_req_mainprn(lnk_buff_dec_128_to_256_ddr_e3_req_mainprn),
    .lnk_buff_dec_128_to_256_ddr_e3_req_mainret(lnk_buff_dec_128_to_256_ddr_e3_req_mainret),
    .lnk_buff_dec_128_to_256_ddr_e3_req_mainse(lnk_buff_dec_128_to_256_ddr_e3_req_mainse),
    .lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainpde(lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainpde),
    .lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainprn(lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainprn),
    .lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainret(lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainret),
    .lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainse(lnk_buff_dec_128_to_256_ddr_e3_req_resp_mainse),
    .lnk_buff_soc_128_to_256_lt_req_mainpde(lnk_buff_soc_128_to_256_lt_req_mainpde),
    .lnk_buff_soc_128_to_256_lt_req_mainprn(lnk_buff_soc_128_to_256_lt_req_mainprn),
    .lnk_buff_soc_128_to_256_lt_req_mainret(lnk_buff_soc_128_to_256_lt_req_mainret),
    .lnk_buff_soc_128_to_256_lt_req_mainse(lnk_buff_soc_128_to_256_lt_req_mainse),
    .lnk_buff_soc_128_to_256_lt_req_resp_mainpde(lnk_buff_soc_128_to_256_lt_req_resp_mainpde),
    .lnk_buff_soc_128_to_256_lt_req_resp_mainprn(lnk_buff_soc_128_to_256_lt_req_resp_mainprn),
    .lnk_buff_soc_128_to_256_lt_req_resp_mainret(lnk_buff_soc_128_to_256_lt_req_resp_mainret),
    .lnk_buff_soc_128_to_256_lt_req_resp_mainse(lnk_buff_soc_128_to_256_lt_req_resp_mainse),
    .lnk_buff_soc_128_to_256_rd_req_resp_mainpde(lnk_buff_soc_128_to_256_rd_req_resp_mainpde),
    .lnk_buff_soc_128_to_256_rd_req_resp_mainprn(lnk_buff_soc_128_to_256_rd_req_resp_mainprn),
    .lnk_buff_soc_128_to_256_rd_req_resp_mainret(lnk_buff_soc_128_to_256_rd_req_resp_mainret),
    .lnk_buff_soc_128_to_256_rd_req_resp_mainse(lnk_buff_soc_128_to_256_rd_req_resp_mainse),
    .lnk_buff_soc_128_to_256_wr_req_mainpde(lnk_buff_soc_128_to_256_wr_req_mainpde),
    .lnk_buff_soc_128_to_256_wr_req_mainprn(lnk_buff_soc_128_to_256_wr_req_mainprn),
    .lnk_buff_soc_128_to_256_wr_req_mainret(lnk_buff_soc_128_to_256_wr_req_mainret),
    .lnk_buff_soc_128_to_256_wr_req_mainse(lnk_buff_soc_128_to_256_wr_req_mainse),
    .lnk_buff_soc_128_to_64_req_mainpde(lnk_buff_soc_128_to_64_req_mainpde),
    .lnk_buff_soc_128_to_64_req_mainprn(lnk_buff_soc_128_to_64_req_mainprn),
    .lnk_buff_soc_128_to_64_req_mainret(lnk_buff_soc_128_to_64_req_mainret),
    .lnk_buff_soc_128_to_64_req_mainse(lnk_buff_soc_128_to_64_req_mainse),
    .lnk_buff_soc_128_to_64_req_resp_mainpde(lnk_buff_soc_128_to_64_req_resp_mainpde),
    .lnk_buff_soc_128_to_64_req_resp_mainprn(lnk_buff_soc_128_to_64_req_resp_mainprn),
    .lnk_buff_soc_128_to_64_req_resp_mainret(lnk_buff_soc_128_to_64_req_resp_mainret),
    .lnk_buff_soc_128_to_64_req_resp_mainse(lnk_buff_soc_128_to_64_req_resp_mainse),
    .lnk_buff_soc_256_to_128_rd_req_resp_mainpde(lnk_buff_soc_256_to_128_rd_req_resp_mainpde),
    .lnk_buff_soc_256_to_128_rd_req_resp_mainprn(lnk_buff_soc_256_to_128_rd_req_resp_mainprn),
    .lnk_buff_soc_256_to_128_rd_req_resp_mainret(lnk_buff_soc_256_to_128_rd_req_resp_mainret),
    .lnk_buff_soc_256_to_128_rd_req_resp_mainse(lnk_buff_soc_256_to_128_rd_req_resp_mainse),
    .lnk_buff_soc_256_to_128_wr_req_mainpde(lnk_buff_soc_256_to_128_wr_req_mainpde),
    .lnk_buff_soc_256_to_128_wr_req_mainprn(lnk_buff_soc_256_to_128_wr_req_mainprn),
    .lnk_buff_soc_256_to_128_wr_req_mainret(lnk_buff_soc_256_to_128_wr_req_mainret),
    .lnk_buff_soc_256_to_128_wr_req_mainse(lnk_buff_soc_256_to_128_wr_req_mainse),
    .lnk_buff_soc_256_to_512_rd_req_resp_mainpde(lnk_buff_soc_256_to_512_rd_req_resp_mainpde),
    .lnk_buff_soc_256_to_512_rd_req_resp_mainprn(lnk_buff_soc_256_to_512_rd_req_resp_mainprn),
    .lnk_buff_soc_256_to_512_rd_req_resp_mainret(lnk_buff_soc_256_to_512_rd_req_resp_mainret),
    .lnk_buff_soc_256_to_512_rd_req_resp_mainse(lnk_buff_soc_256_to_512_rd_req_resp_mainse),
    .lnk_buff_soc_256_to_512_wr_req_mainpde(lnk_buff_soc_256_to_512_wr_req_mainpde),
    .lnk_buff_soc_256_to_512_wr_req_mainprn(lnk_buff_soc_256_to_512_wr_req_mainprn),
    .lnk_buff_soc_256_to_512_wr_req_mainret(lnk_buff_soc_256_to_512_wr_req_mainret),
    .lnk_buff_soc_256_to_512_wr_req_mainse(lnk_buff_soc_256_to_512_wr_req_mainse),
    .lnk_buff_soc_512_to_256_ddr_e0_req_mainpde(lnk_buff_soc_512_to_256_ddr_e0_req_mainpde),
    .lnk_buff_soc_512_to_256_ddr_e0_req_mainprn(lnk_buff_soc_512_to_256_ddr_e0_req_mainprn),
    .lnk_buff_soc_512_to_256_ddr_e0_req_mainret(lnk_buff_soc_512_to_256_ddr_e0_req_mainret),
    .lnk_buff_soc_512_to_256_ddr_e0_req_mainse(lnk_buff_soc_512_to_256_ddr_e0_req_mainse),
    .lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainpde(lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainpde),
    .lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainprn(lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainprn),
    .lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainret(lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainret),
    .lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainse(lnk_buff_soc_512_to_256_ddr_e0_req_resp_mainse),
    .lnk_buff_soc_512_to_256_ddr_e1_req_mainpde(lnk_buff_soc_512_to_256_ddr_e1_req_mainpde),
    .lnk_buff_soc_512_to_256_ddr_e1_req_mainprn(lnk_buff_soc_512_to_256_ddr_e1_req_mainprn),
    .lnk_buff_soc_512_to_256_ddr_e1_req_mainret(lnk_buff_soc_512_to_256_ddr_e1_req_mainret),
    .lnk_buff_soc_512_to_256_ddr_e1_req_mainse(lnk_buff_soc_512_to_256_ddr_e1_req_mainse),
    .lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainpde(lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainpde),
    .lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainprn(lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainprn),
    .lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainret(lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainret),
    .lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainse(lnk_buff_soc_512_to_256_ddr_e1_req_resp_mainse),
    .lnk_buff_soc_512_to_256_ddr_e2_req_mainpde(lnk_buff_soc_512_to_256_ddr_e2_req_mainpde),
    .lnk_buff_soc_512_to_256_ddr_e2_req_mainprn(lnk_buff_soc_512_to_256_ddr_e2_req_mainprn),
    .lnk_buff_soc_512_to_256_ddr_e2_req_mainret(lnk_buff_soc_512_to_256_ddr_e2_req_mainret),
    .lnk_buff_soc_512_to_256_ddr_e2_req_mainse(lnk_buff_soc_512_to_256_ddr_e2_req_mainse),
    .lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainpde(lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainpde),
    .lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainprn(lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainprn),
    .lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainret(lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainret),
    .lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainse(lnk_buff_soc_512_to_256_ddr_e2_req_resp_mainse),
    .lnk_buff_soc_512_to_256_ddr_e3_req_mainpde(lnk_buff_soc_512_to_256_ddr_e3_req_mainpde),
    .lnk_buff_soc_512_to_256_ddr_e3_req_mainprn(lnk_buff_soc_512_to_256_ddr_e3_req_mainprn),
    .lnk_buff_soc_512_to_256_ddr_e3_req_mainret(lnk_buff_soc_512_to_256_ddr_e3_req_mainret),
    .lnk_buff_soc_512_to_256_ddr_e3_req_mainse(lnk_buff_soc_512_to_256_ddr_e3_req_mainse),
    .lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainpde(lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainpde),
    .lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainprn(lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainprn),
    .lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainret(lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainret),
    .lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainse(lnk_buff_soc_512_to_256_ddr_e3_req_resp_mainse),
    .lnk_buff_soc_512_to_256_rd_req_resp_mainpde(lnk_buff_soc_512_to_256_rd_req_resp_mainpde),
    .lnk_buff_soc_512_to_256_rd_req_resp_mainprn(lnk_buff_soc_512_to_256_rd_req_resp_mainprn),
    .lnk_buff_soc_512_to_256_rd_req_resp_mainret(lnk_buff_soc_512_to_256_rd_req_resp_mainret),
    .lnk_buff_soc_512_to_256_rd_req_resp_mainse(lnk_buff_soc_512_to_256_rd_req_resp_mainse),
    .lnk_buff_soc_512_to_256_wr_req_mainpde(lnk_buff_soc_512_to_256_wr_req_mainpde),
    .lnk_buff_soc_512_to_256_wr_req_mainprn(lnk_buff_soc_512_to_256_wr_req_mainprn),
    .lnk_buff_soc_512_to_256_wr_req_mainret(lnk_buff_soc_512_to_256_wr_req_mainret),
    .lnk_buff_soc_512_to_256_wr_req_mainse(lnk_buff_soc_512_to_256_wr_req_mainse),
    .lnk_buff_soc_64_to_128_lt_req_mainpde(lnk_buff_soc_64_to_128_lt_req_mainpde),
    .lnk_buff_soc_64_to_128_lt_req_mainprn(lnk_buff_soc_64_to_128_lt_req_mainprn),
    .lnk_buff_soc_64_to_128_lt_req_mainret(lnk_buff_soc_64_to_128_lt_req_mainret),
    .lnk_buff_soc_64_to_128_lt_req_mainse(lnk_buff_soc_64_to_128_lt_req_mainse),
    .lnk_buff_soc_64_to_128_lt_req_resp_mainpde(lnk_buff_soc_64_to_128_lt_req_resp_mainpde),
    .lnk_buff_soc_64_to_128_lt_req_resp_mainprn(lnk_buff_soc_64_to_128_lt_req_resp_mainprn),
    .lnk_buff_soc_64_to_128_lt_req_resp_mainret(lnk_buff_soc_64_to_128_lt_req_resp_mainret),
    .lnk_buff_soc_64_to_128_lt_req_resp_mainse(lnk_buff_soc_64_to_128_lt_req_resp_mainse),
    .lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
    .lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
    .lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
    .lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
    .lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
    .lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
    .lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
    .lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
    .noc_clk(i_noc_clk),
    .noc_rst_n(i_noc_rst_n),
    .pcie_aon_clk(i_pcie_aon_clk),
    .pcie_aon_rst_n(i_pcie_aon_rst_n),
    .pcie_init_mt_clk(i_pcie_init_mt_clk),
    .pcie_init_mt_clken(i_pcie_init_mt_clken),
    .pcie_init_mt_pwr_Idle(o_pcie_init_mt_pwr_idle_val),
    .pcie_init_mt_pwr_IdleAck(o_pcie_init_mt_pwr_idle_ack),
    .pcie_init_mt_pwr_IdleReq(i_pcie_init_mt_pwr_idle_req),
    .pcie_init_mt_rd_Ar_Addr(pcie_init_mt_axi_s_araddr_msb_fixed),
    .pcie_init_mt_rd_Ar_Burst(i_pcie_init_mt_axi_s_arburst),
    .pcie_init_mt_rd_Ar_Cache(i_pcie_init_mt_axi_s_arcache),
    .pcie_init_mt_rd_Ar_Id(i_pcie_init_mt_axi_s_arid),
    .pcie_init_mt_rd_Ar_Len(i_pcie_init_mt_axi_s_arlen),
    .pcie_init_mt_rd_Ar_Lock(i_pcie_init_mt_axi_s_arlock),
    .pcie_init_mt_rd_Ar_Prot(i_pcie_init_mt_axi_s_arprot),
    .pcie_init_mt_rd_Ar_Qos(i_pcie_init_mt_axi_s_arqos),
    .pcie_init_mt_rd_Ar_Ready(o_pcie_init_mt_axi_s_arready),
    .pcie_init_mt_rd_Ar_Size(i_pcie_init_mt_axi_s_arsize),
    .pcie_init_mt_rd_Ar_Valid(i_pcie_init_mt_axi_s_arvalid),
    .pcie_init_mt_rd_R_Data(o_pcie_init_mt_axi_s_rdata),
    .pcie_init_mt_rd_R_Id(o_pcie_init_mt_axi_s_rid),
    .pcie_init_mt_rd_R_Last(o_pcie_init_mt_axi_s_rlast),
    .pcie_init_mt_rd_R_Ready(i_pcie_init_mt_axi_s_rready),
    .pcie_init_mt_rd_R_Resp(o_pcie_init_mt_axi_s_rresp),
    .pcie_init_mt_rd_R_Valid(o_pcie_init_mt_axi_s_rvalid),
    .pcie_init_mt_rst_n(i_pcie_init_mt_rst_n),
    .pcie_init_mt_wr_Aw_Addr(pcie_init_mt_axi_s_awaddr_msb_fixed),
    .pcie_init_mt_wr_Aw_Burst(i_pcie_init_mt_axi_s_awburst),
    .pcie_init_mt_wr_Aw_Cache(i_pcie_init_mt_axi_s_awcache),
    .pcie_init_mt_wr_Aw_Id(i_pcie_init_mt_axi_s_awid),
    .pcie_init_mt_wr_Aw_Len(i_pcie_init_mt_axi_s_awlen),
    .pcie_init_mt_wr_Aw_Lock(i_pcie_init_mt_axi_s_awlock),
    .pcie_init_mt_wr_Aw_Prot(i_pcie_init_mt_axi_s_awprot),
    .pcie_init_mt_wr_Aw_Qos(i_pcie_init_mt_axi_s_awqos),
    .pcie_init_mt_wr_Aw_Ready(o_pcie_init_mt_axi_s_awready),
    .pcie_init_mt_wr_Aw_Size(i_pcie_init_mt_axi_s_awsize),
    .pcie_init_mt_wr_Aw_Valid(i_pcie_init_mt_axi_s_awvalid),
    .pcie_init_mt_wr_B_Id(o_pcie_init_mt_axi_s_bid),
    .pcie_init_mt_wr_B_Ready(i_pcie_init_mt_axi_s_bready),
    .pcie_init_mt_wr_B_Resp(o_pcie_init_mt_axi_s_bresp),
    .pcie_init_mt_wr_B_Valid(o_pcie_init_mt_axi_s_bvalid),
    .pcie_init_mt_wr_W_Data(i_pcie_init_mt_axi_s_wdata),
    .pcie_init_mt_wr_W_Last(i_pcie_init_mt_axi_s_wlast),
    .pcie_init_mt_wr_W_Ready(o_pcie_init_mt_axi_s_wready),
    .pcie_init_mt_wr_W_Strb(i_pcie_init_mt_axi_s_wstrb),
    .pcie_init_mt_wr_W_Valid(i_pcie_init_mt_axi_s_wvalid),
    .pcie_targ_cfg_PAddr(o_pcie_targ_cfg_apb_m_paddr),
    .pcie_targ_cfg_PEnable(o_pcie_targ_cfg_apb_m_penable),
    .pcie_targ_cfg_PProt(o_pcie_targ_cfg_apb_m_pprot),
    .pcie_targ_cfg_PRData(i_pcie_targ_cfg_apb_m_prdata),
    .pcie_targ_cfg_PReady(i_pcie_targ_cfg_apb_m_pready),
    .pcie_targ_cfg_PSel(o_pcie_targ_cfg_apb_m_psel),
    .pcie_targ_cfg_PSlvErr(i_pcie_targ_cfg_apb_m_pslverr),
    .pcie_targ_cfg_PStrb(o_pcie_targ_cfg_apb_m_pstrb),
    .pcie_targ_cfg_PWData(o_pcie_targ_cfg_apb_m_pwdata),
    .pcie_targ_cfg_PWrite(o_pcie_targ_cfg_apb_m_pwrite),
    .pcie_targ_cfg_clk(i_pcie_targ_cfg_clk),
    .pcie_targ_cfg_clken(i_pcie_targ_cfg_clken),
    .pcie_targ_cfg_dbi_Ar_Addr(pcie_targ_cfg_dbi_axi_m_araddr_msb_fixed),
    .pcie_targ_cfg_dbi_Ar_Burst(o_pcie_targ_cfg_dbi_axi_m_arburst),
    .pcie_targ_cfg_dbi_Ar_Cache(o_pcie_targ_cfg_dbi_axi_m_arcache),
    .pcie_targ_cfg_dbi_Ar_Id(o_pcie_targ_cfg_dbi_axi_m_arid),
    .pcie_targ_cfg_dbi_Ar_Len(o_pcie_targ_cfg_dbi_axi_m_arlen),
    .pcie_targ_cfg_dbi_Ar_Lock(o_pcie_targ_cfg_dbi_axi_m_arlock),
    .pcie_targ_cfg_dbi_Ar_Prot(o_pcie_targ_cfg_dbi_axi_m_arprot),
    .pcie_targ_cfg_dbi_Ar_Qos(o_pcie_targ_cfg_dbi_axi_m_arqos),
    .pcie_targ_cfg_dbi_Ar_Ready(i_pcie_targ_cfg_dbi_axi_m_arready),
    .pcie_targ_cfg_dbi_Ar_Size(o_pcie_targ_cfg_dbi_axi_m_arsize),
    .pcie_targ_cfg_dbi_Ar_Valid(o_pcie_targ_cfg_dbi_axi_m_arvalid),
    .pcie_targ_cfg_dbi_Aw_Addr(pcie_targ_cfg_dbi_axi_m_awaddr_msb_fixed),
    .pcie_targ_cfg_dbi_Aw_Burst(o_pcie_targ_cfg_dbi_axi_m_awburst),
    .pcie_targ_cfg_dbi_Aw_Cache(o_pcie_targ_cfg_dbi_axi_m_awcache),
    .pcie_targ_cfg_dbi_Aw_Id(o_pcie_targ_cfg_dbi_axi_m_awid),
    .pcie_targ_cfg_dbi_Aw_Len(o_pcie_targ_cfg_dbi_axi_m_awlen),
    .pcie_targ_cfg_dbi_Aw_Lock(o_pcie_targ_cfg_dbi_axi_m_awlock),
    .pcie_targ_cfg_dbi_Aw_Prot(o_pcie_targ_cfg_dbi_axi_m_awprot),
    .pcie_targ_cfg_dbi_Aw_Qos(o_pcie_targ_cfg_dbi_axi_m_awqos),
    .pcie_targ_cfg_dbi_Aw_Ready(i_pcie_targ_cfg_dbi_axi_m_awready),
    .pcie_targ_cfg_dbi_Aw_Size(o_pcie_targ_cfg_dbi_axi_m_awsize),
    .pcie_targ_cfg_dbi_Aw_Valid(o_pcie_targ_cfg_dbi_axi_m_awvalid),
    .pcie_targ_cfg_dbi_B_Id(i_pcie_targ_cfg_dbi_axi_m_bid),
    .pcie_targ_cfg_dbi_B_Ready(o_pcie_targ_cfg_dbi_axi_m_bready),
    .pcie_targ_cfg_dbi_B_Resp(i_pcie_targ_cfg_dbi_axi_m_bresp),
    .pcie_targ_cfg_dbi_B_Valid(i_pcie_targ_cfg_dbi_axi_m_bvalid),
    .pcie_targ_cfg_dbi_R_Data(i_pcie_targ_cfg_dbi_axi_m_rdata),
    .pcie_targ_cfg_dbi_R_Id(i_pcie_targ_cfg_dbi_axi_m_rid),
    .pcie_targ_cfg_dbi_R_Last(i_pcie_targ_cfg_dbi_axi_m_rlast),
    .pcie_targ_cfg_dbi_R_Ready(o_pcie_targ_cfg_dbi_axi_m_rready),
    .pcie_targ_cfg_dbi_R_Resp(i_pcie_targ_cfg_dbi_axi_m_rresp),
    .pcie_targ_cfg_dbi_R_Valid(i_pcie_targ_cfg_dbi_axi_m_rvalid),
    .pcie_targ_cfg_dbi_W_Data(o_pcie_targ_cfg_dbi_axi_m_wdata),
    .pcie_targ_cfg_dbi_W_Last(o_pcie_targ_cfg_dbi_axi_m_wlast),
    .pcie_targ_cfg_dbi_W_Ready(i_pcie_targ_cfg_dbi_axi_m_wready),
    .pcie_targ_cfg_dbi_W_Strb(o_pcie_targ_cfg_dbi_axi_m_wstrb),
    .pcie_targ_cfg_dbi_W_Valid(o_pcie_targ_cfg_dbi_axi_m_wvalid),
    .pcie_targ_cfg_dbi_clk(i_pcie_targ_cfg_dbi_clk),
    .pcie_targ_cfg_dbi_clken(i_pcie_targ_cfg_dbi_clken),
    .pcie_targ_cfg_dbi_pwr_Idle(o_pcie_targ_cfg_dbi_pwr_idle_val),
    .pcie_targ_cfg_dbi_pwr_IdleAck(o_pcie_targ_cfg_dbi_pwr_idle_ack),
    .pcie_targ_cfg_dbi_pwr_IdleReq(i_pcie_targ_cfg_dbi_pwr_idle_req),
    .pcie_targ_cfg_dbi_rst_n(i_pcie_targ_cfg_dbi_rst_n),
    .pcie_targ_cfg_pwr_Idle(o_pcie_targ_cfg_pwr_idle_val),
    .pcie_targ_cfg_pwr_IdleAck(o_pcie_targ_cfg_pwr_idle_ack),
    .pcie_targ_cfg_pwr_IdleReq(i_pcie_targ_cfg_pwr_idle_req),
    .pcie_targ_cfg_rst_n(i_pcie_targ_cfg_rst_n),
    .pcie_targ_mt_clk(i_pcie_targ_mt_clk),
    .pcie_targ_mt_clken(i_pcie_targ_mt_clken),
    .pcie_targ_mt_pwr_Idle(o_pcie_targ_mt_pwr_idle_val),
    .pcie_targ_mt_pwr_IdleAck(o_pcie_targ_mt_pwr_idle_ack),
    .pcie_targ_mt_pwr_IdleReq(i_pcie_targ_mt_pwr_idle_req),
    .pcie_targ_mt_rd_Ar_Addr(pcie_targ_mt_axi_m_araddr_msb_fixed),
    .pcie_targ_mt_rd_Ar_Burst(o_pcie_targ_mt_axi_m_arburst),
    .pcie_targ_mt_rd_Ar_Cache(o_pcie_targ_mt_axi_m_arcache),
    .pcie_targ_mt_rd_Ar_Id(o_pcie_targ_mt_axi_m_arid),
    .pcie_targ_mt_rd_Ar_Len(o_pcie_targ_mt_axi_m_arlen),
    .pcie_targ_mt_rd_Ar_Lock(o_pcie_targ_mt_axi_m_arlock),
    .pcie_targ_mt_rd_Ar_Prot(o_pcie_targ_mt_axi_m_arprot),
    .pcie_targ_mt_rd_Ar_Qos(o_pcie_targ_mt_axi_m_arqos),
    .pcie_targ_mt_rd_Ar_Ready(i_pcie_targ_mt_axi_m_arready),
    .pcie_targ_mt_rd_Ar_Size(o_pcie_targ_mt_axi_m_arsize),
    .pcie_targ_mt_rd_Ar_Valid(o_pcie_targ_mt_axi_m_arvalid),
    .pcie_targ_mt_rd_R_Data(i_pcie_targ_mt_axi_m_rdata),
    .pcie_targ_mt_rd_R_Id(i_pcie_targ_mt_axi_m_rid),
    .pcie_targ_mt_rd_R_Last(i_pcie_targ_mt_axi_m_rlast),
    .pcie_targ_mt_rd_R_Ready(o_pcie_targ_mt_axi_m_rready),
    .pcie_targ_mt_rd_R_Resp(i_pcie_targ_mt_axi_m_rresp),
    .pcie_targ_mt_rd_R_Valid(i_pcie_targ_mt_axi_m_rvalid),
    .pcie_targ_mt_rst_n(i_pcie_targ_mt_rst_n),
    .pcie_targ_mt_wr_Aw_Addr(pcie_targ_mt_axi_m_awaddr_msb_fixed),
    .pcie_targ_mt_wr_Aw_Burst(o_pcie_targ_mt_axi_m_awburst),
    .pcie_targ_mt_wr_Aw_Cache(o_pcie_targ_mt_axi_m_awcache),
    .pcie_targ_mt_wr_Aw_Id(o_pcie_targ_mt_axi_m_awid),
    .pcie_targ_mt_wr_Aw_Len(o_pcie_targ_mt_axi_m_awlen),
    .pcie_targ_mt_wr_Aw_Lock(o_pcie_targ_mt_axi_m_awlock),
    .pcie_targ_mt_wr_Aw_Prot(o_pcie_targ_mt_axi_m_awprot),
    .pcie_targ_mt_wr_Aw_Qos(o_pcie_targ_mt_axi_m_awqos),
    .pcie_targ_mt_wr_Aw_Ready(i_pcie_targ_mt_axi_m_awready),
    .pcie_targ_mt_wr_Aw_Size(o_pcie_targ_mt_axi_m_awsize),
    .pcie_targ_mt_wr_Aw_Valid(o_pcie_targ_mt_axi_m_awvalid),
    .pcie_targ_mt_wr_B_Id(i_pcie_targ_mt_axi_m_bid),
    .pcie_targ_mt_wr_B_Ready(o_pcie_targ_mt_axi_m_bready),
    .pcie_targ_mt_wr_B_Resp(i_pcie_targ_mt_axi_m_bresp),
    .pcie_targ_mt_wr_B_Valid(i_pcie_targ_mt_axi_m_bvalid),
    .pcie_targ_mt_wr_W_Data(o_pcie_targ_mt_axi_m_wdata),
    .pcie_targ_mt_wr_W_Last(o_pcie_targ_mt_axi_m_wlast),
    .pcie_targ_mt_wr_W_Ready(i_pcie_targ_mt_axi_m_wready),
    .pcie_targ_mt_wr_W_Strb(o_pcie_targ_mt_axi_m_wstrb),
    .pcie_targ_mt_wr_W_Valid(o_pcie_targ_mt_axi_m_wvalid),
    .pcie_targ_syscfg_PAddr(o_pcie_targ_syscfg_apb_m_paddr),
    .pcie_targ_syscfg_PEnable(o_pcie_targ_syscfg_apb_m_penable),
    .pcie_targ_syscfg_PProt(o_pcie_targ_syscfg_apb_m_pprot),
    .pcie_targ_syscfg_PRData(i_pcie_targ_syscfg_apb_m_prdata),
    .pcie_targ_syscfg_PReady(i_pcie_targ_syscfg_apb_m_pready),
    .pcie_targ_syscfg_PSel(o_pcie_targ_syscfg_apb_m_psel),
    .pcie_targ_syscfg_PSlvErr(i_pcie_targ_syscfg_apb_m_pslverr),
    .pcie_targ_syscfg_PStrb(o_pcie_targ_syscfg_apb_m_pstrb),
    .pcie_targ_syscfg_PWData(o_pcie_targ_syscfg_apb_m_pwdata),
    .pcie_targ_syscfg_PWrite(o_pcie_targ_syscfg_apb_m_pwrite),
    .pve_0_aon_clk(i_pve_0_aon_clk),
    .pve_0_aon_rst_n(i_pve_0_aon_rst_n),
    .pve_0_clk(i_pve_0_clk),
    .pve_0_clken(i_pve_0_clken),
    .pve_0_init_ht_rd_Ar_Addr(pve_0_init_ht_axi_s_araddr_msb_fixed),
    .pve_0_init_ht_rd_Ar_Burst(i_pve_0_init_ht_axi_s_arburst),
    .pve_0_init_ht_rd_Ar_Cache(i_pve_0_init_ht_axi_s_arcache),
    .pve_0_init_ht_rd_Ar_Id(i_pve_0_init_ht_axi_s_arid),
    .pve_0_init_ht_rd_Ar_Len(i_pve_0_init_ht_axi_s_arlen),
    .pve_0_init_ht_rd_Ar_Lock(i_pve_0_init_ht_axi_s_arlock),
    .pve_0_init_ht_rd_Ar_Prot(i_pve_0_init_ht_axi_s_arprot),
    .pve_0_init_ht_rd_Ar_Ready(o_pve_0_init_ht_axi_s_arready),
    .pve_0_init_ht_rd_Ar_Size(i_pve_0_init_ht_axi_s_arsize),
    .pve_0_init_ht_rd_Ar_Valid(i_pve_0_init_ht_axi_s_arvalid),
    .pve_0_init_ht_rd_R_Data(o_pve_0_init_ht_axi_s_rdata),
    .pve_0_init_ht_rd_R_Id(o_pve_0_init_ht_axi_s_rid),
    .pve_0_init_ht_rd_R_Last(o_pve_0_init_ht_axi_s_rlast),
    .pve_0_init_ht_rd_R_Ready(i_pve_0_init_ht_axi_s_rready),
    .pve_0_init_ht_rd_R_Resp(o_pve_0_init_ht_axi_s_rresp),
    .pve_0_init_ht_rd_R_Valid(o_pve_0_init_ht_axi_s_rvalid),
    .pve_0_init_ht_wr_Aw_Addr(pve_0_init_ht_axi_s_awaddr_msb_fixed),
    .pve_0_init_ht_wr_Aw_Burst(i_pve_0_init_ht_axi_s_awburst),
    .pve_0_init_ht_wr_Aw_Cache(i_pve_0_init_ht_axi_s_awcache),
    .pve_0_init_ht_wr_Aw_Id(i_pve_0_init_ht_axi_s_awid),
    .pve_0_init_ht_wr_Aw_Len(i_pve_0_init_ht_axi_s_awlen),
    .pve_0_init_ht_wr_Aw_Lock(i_pve_0_init_ht_axi_s_awlock),
    .pve_0_init_ht_wr_Aw_Prot(i_pve_0_init_ht_axi_s_awprot),
    .pve_0_init_ht_wr_Aw_Ready(o_pve_0_init_ht_axi_s_awready),
    .pve_0_init_ht_wr_Aw_Size(i_pve_0_init_ht_axi_s_awsize),
    .pve_0_init_ht_wr_Aw_Valid(i_pve_0_init_ht_axi_s_awvalid),
    .pve_0_init_ht_wr_B_Id(o_pve_0_init_ht_axi_s_bid),
    .pve_0_init_ht_wr_B_Ready(i_pve_0_init_ht_axi_s_bready),
    .pve_0_init_ht_wr_B_Resp(o_pve_0_init_ht_axi_s_bresp),
    .pve_0_init_ht_wr_B_Valid(o_pve_0_init_ht_axi_s_bvalid),
    .pve_0_init_ht_wr_W_Data(i_pve_0_init_ht_axi_s_wdata),
    .pve_0_init_ht_wr_W_Last(i_pve_0_init_ht_axi_s_wlast),
    .pve_0_init_ht_wr_W_Ready(o_pve_0_init_ht_axi_s_wready),
    .pve_0_init_ht_wr_W_Strb(i_pve_0_init_ht_axi_s_wstrb),
    .pve_0_init_ht_wr_W_Valid(i_pve_0_init_ht_axi_s_wvalid),
    .pve_0_init_lt_rd_Ar_Addr(pve_0_init_lt_axi_s_araddr_msb_fixed),
    .pve_0_init_lt_rd_Ar_Burst(i_pve_0_init_lt_axi_s_arburst),
    .pve_0_init_lt_rd_Ar_Cache(i_pve_0_init_lt_axi_s_arcache),
    .pve_0_init_lt_rd_Ar_Id(i_pve_0_init_lt_axi_s_arid),
    .pve_0_init_lt_rd_Ar_Len(i_pve_0_init_lt_axi_s_arlen),
    .pve_0_init_lt_rd_Ar_Lock(i_pve_0_init_lt_axi_s_arlock),
    .pve_0_init_lt_rd_Ar_Prot(i_pve_0_init_lt_axi_s_arprot),
    .pve_0_init_lt_rd_Ar_Qos(i_pve_0_init_lt_axi_s_arqos),
    .pve_0_init_lt_rd_Ar_Ready(o_pve_0_init_lt_axi_s_arready),
    .pve_0_init_lt_rd_Ar_Size(i_pve_0_init_lt_axi_s_arsize),
    .pve_0_init_lt_rd_Ar_User(pve_0_init_lt_axi_s_aruser),
    .pve_0_init_lt_rd_Ar_Valid(i_pve_0_init_lt_axi_s_arvalid),
    .pve_0_init_lt_rd_R_Data(o_pve_0_init_lt_axi_s_rdata),
    .pve_0_init_lt_rd_R_Id(o_pve_0_init_lt_axi_s_rid),
    .pve_0_init_lt_rd_R_Last(o_pve_0_init_lt_axi_s_rlast),
    .pve_0_init_lt_rd_R_Ready(i_pve_0_init_lt_axi_s_rready),
    .pve_0_init_lt_rd_R_Resp(o_pve_0_init_lt_axi_s_rresp),
    .pve_0_init_lt_rd_R_Valid(o_pve_0_init_lt_axi_s_rvalid),
    .pve_0_init_lt_wr_Aw_Addr(pve_0_init_lt_axi_s_awaddr_msb_fixed),
    .pve_0_init_lt_wr_Aw_Burst(i_pve_0_init_lt_axi_s_awburst),
    .pve_0_init_lt_wr_Aw_Cache(i_pve_0_init_lt_axi_s_awcache),
    .pve_0_init_lt_wr_Aw_Id(i_pve_0_init_lt_axi_s_awid),
    .pve_0_init_lt_wr_Aw_Len(i_pve_0_init_lt_axi_s_awlen),
    .pve_0_init_lt_wr_Aw_Lock(i_pve_0_init_lt_axi_s_awlock),
    .pve_0_init_lt_wr_Aw_Prot(i_pve_0_init_lt_axi_s_awprot),
    .pve_0_init_lt_wr_Aw_Qos(i_pve_0_init_lt_axi_s_awqos),
    .pve_0_init_lt_wr_Aw_Ready(o_pve_0_init_lt_axi_s_awready),
    .pve_0_init_lt_wr_Aw_Size(i_pve_0_init_lt_axi_s_awsize),
    .pve_0_init_lt_wr_Aw_User(pve_0_init_lt_axi_s_awuser),
    .pve_0_init_lt_wr_Aw_Valid(i_pve_0_init_lt_axi_s_awvalid),
    .pve_0_init_lt_wr_B_Id(o_pve_0_init_lt_axi_s_bid),
    .pve_0_init_lt_wr_B_Ready(i_pve_0_init_lt_axi_s_bready),
    .pve_0_init_lt_wr_B_Resp(o_pve_0_init_lt_axi_s_bresp),
    .pve_0_init_lt_wr_B_Valid(o_pve_0_init_lt_axi_s_bvalid),
    .pve_0_init_lt_wr_W_Data(i_pve_0_init_lt_axi_s_wdata),
    .pve_0_init_lt_wr_W_Last(i_pve_0_init_lt_axi_s_wlast),
    .pve_0_init_lt_wr_W_Ready(o_pve_0_init_lt_axi_s_wready),
    .pve_0_init_lt_wr_W_Strb(i_pve_0_init_lt_axi_s_wstrb),
    .pve_0_init_lt_wr_W_Valid(i_pve_0_init_lt_axi_s_wvalid),
    .pve_0_pwr_Idle(o_pve_0_pwr_idle_val),
    .pve_0_pwr_IdleAck(o_pve_0_pwr_idle_ack),
    .pve_0_pwr_IdleReq(i_pve_0_pwr_idle_req),
    .pve_0_rst_n(i_pve_0_rst_n),
    .pve_0_targ_lt_Ar_Addr(pve_0_targ_lt_axi_m_araddr_msb_fixed),
    .pve_0_targ_lt_Ar_Burst(o_pve_0_targ_lt_axi_m_arburst),
    .pve_0_targ_lt_Ar_Cache(o_pve_0_targ_lt_axi_m_arcache),
    .pve_0_targ_lt_Ar_Id(o_pve_0_targ_lt_axi_m_arid),
    .pve_0_targ_lt_Ar_Len(o_pve_0_targ_lt_axi_m_arlen),
    .pve_0_targ_lt_Ar_Lock(o_pve_0_targ_lt_axi_m_arlock),
    .pve_0_targ_lt_Ar_Prot(o_pve_0_targ_lt_axi_m_arprot),
    .pve_0_targ_lt_Ar_Qos(o_pve_0_targ_lt_axi_m_arqos),
    .pve_0_targ_lt_Ar_Ready(i_pve_0_targ_lt_axi_m_arready),
    .pve_0_targ_lt_Ar_Size(o_pve_0_targ_lt_axi_m_arsize),
    .pve_0_targ_lt_Ar_Valid(o_pve_0_targ_lt_axi_m_arvalid),
    .pve_0_targ_lt_Aw_Addr(pve_0_targ_lt_axi_m_awaddr_msb_fixed),
    .pve_0_targ_lt_Aw_Burst(o_pve_0_targ_lt_axi_m_awburst),
    .pve_0_targ_lt_Aw_Cache(o_pve_0_targ_lt_axi_m_awcache),
    .pve_0_targ_lt_Aw_Id(o_pve_0_targ_lt_axi_m_awid),
    .pve_0_targ_lt_Aw_Len(o_pve_0_targ_lt_axi_m_awlen),
    .pve_0_targ_lt_Aw_Lock(o_pve_0_targ_lt_axi_m_awlock),
    .pve_0_targ_lt_Aw_Prot(o_pve_0_targ_lt_axi_m_awprot),
    .pve_0_targ_lt_Aw_Qos(o_pve_0_targ_lt_axi_m_awqos),
    .pve_0_targ_lt_Aw_Ready(i_pve_0_targ_lt_axi_m_awready),
    .pve_0_targ_lt_Aw_Size(o_pve_0_targ_lt_axi_m_awsize),
    .pve_0_targ_lt_Aw_Valid(o_pve_0_targ_lt_axi_m_awvalid),
    .pve_0_targ_lt_B_Id(i_pve_0_targ_lt_axi_m_bid),
    .pve_0_targ_lt_B_Ready(o_pve_0_targ_lt_axi_m_bready),
    .pve_0_targ_lt_B_Resp(i_pve_0_targ_lt_axi_m_bresp),
    .pve_0_targ_lt_B_Valid(i_pve_0_targ_lt_axi_m_bvalid),
    .pve_0_targ_lt_R_Data(i_pve_0_targ_lt_axi_m_rdata),
    .pve_0_targ_lt_R_Id(i_pve_0_targ_lt_axi_m_rid),
    .pve_0_targ_lt_R_Last(i_pve_0_targ_lt_axi_m_rlast),
    .pve_0_targ_lt_R_Ready(o_pve_0_targ_lt_axi_m_rready),
    .pve_0_targ_lt_R_Resp(i_pve_0_targ_lt_axi_m_rresp),
    .pve_0_targ_lt_R_Valid(i_pve_0_targ_lt_axi_m_rvalid),
    .pve_0_targ_lt_W_Data(o_pve_0_targ_lt_axi_m_wdata),
    .pve_0_targ_lt_W_Last(o_pve_0_targ_lt_axi_m_wlast),
    .pve_0_targ_lt_W_Ready(i_pve_0_targ_lt_axi_m_wready),
    .pve_0_targ_lt_W_Strb(o_pve_0_targ_lt_axi_m_wstrb),
    .pve_0_targ_lt_W_Valid(o_pve_0_targ_lt_axi_m_wvalid),
    .pve_0_targ_syscfg_PAddr(o_pve_0_targ_syscfg_apb_m_paddr),
    .pve_0_targ_syscfg_PEnable(o_pve_0_targ_syscfg_apb_m_penable),
    .pve_0_targ_syscfg_PProt(o_pve_0_targ_syscfg_apb_m_pprot),
    .pve_0_targ_syscfg_PRData(i_pve_0_targ_syscfg_apb_m_prdata),
    .pve_0_targ_syscfg_PReady(i_pve_0_targ_syscfg_apb_m_pready),
    .pve_0_targ_syscfg_PSel(o_pve_0_targ_syscfg_apb_m_psel),
    .pve_0_targ_syscfg_PSlvErr(i_pve_0_targ_syscfg_apb_m_pslverr),
    .pve_0_targ_syscfg_PStrb(o_pve_0_targ_syscfg_apb_m_pstrb),
    .pve_0_targ_syscfg_PWData(o_pve_0_targ_syscfg_apb_m_pwdata),
    .pve_0_targ_syscfg_PWrite(o_pve_0_targ_syscfg_apb_m_pwrite),
    .pve_1_aon_clk(i_pve_1_aon_clk),
    .pve_1_aon_rst_n(i_pve_1_aon_rst_n),
    .pve_1_clk(i_pve_1_clk),
    .pve_1_clken(i_pve_1_clken),
    .pve_1_init_ht_rd_Ar_Addr(pve_1_init_ht_axi_s_araddr_msb_fixed),
    .pve_1_init_ht_rd_Ar_Burst(i_pve_1_init_ht_axi_s_arburst),
    .pve_1_init_ht_rd_Ar_Cache(i_pve_1_init_ht_axi_s_arcache),
    .pve_1_init_ht_rd_Ar_Id(i_pve_1_init_ht_axi_s_arid),
    .pve_1_init_ht_rd_Ar_Len(i_pve_1_init_ht_axi_s_arlen),
    .pve_1_init_ht_rd_Ar_Lock(i_pve_1_init_ht_axi_s_arlock),
    .pve_1_init_ht_rd_Ar_Prot(i_pve_1_init_ht_axi_s_arprot),
    .pve_1_init_ht_rd_Ar_Ready(o_pve_1_init_ht_axi_s_arready),
    .pve_1_init_ht_rd_Ar_Size(i_pve_1_init_ht_axi_s_arsize),
    .pve_1_init_ht_rd_Ar_Valid(i_pve_1_init_ht_axi_s_arvalid),
    .pve_1_init_ht_rd_R_Data(o_pve_1_init_ht_axi_s_rdata),
    .pve_1_init_ht_rd_R_Id(o_pve_1_init_ht_axi_s_rid),
    .pve_1_init_ht_rd_R_Last(o_pve_1_init_ht_axi_s_rlast),
    .pve_1_init_ht_rd_R_Ready(i_pve_1_init_ht_axi_s_rready),
    .pve_1_init_ht_rd_R_Resp(o_pve_1_init_ht_axi_s_rresp),
    .pve_1_init_ht_rd_R_Valid(o_pve_1_init_ht_axi_s_rvalid),
    .pve_1_init_ht_wr_Aw_Addr(pve_1_init_ht_axi_s_awaddr_msb_fixed),
    .pve_1_init_ht_wr_Aw_Burst(i_pve_1_init_ht_axi_s_awburst),
    .pve_1_init_ht_wr_Aw_Cache(i_pve_1_init_ht_axi_s_awcache),
    .pve_1_init_ht_wr_Aw_Id(i_pve_1_init_ht_axi_s_awid),
    .pve_1_init_ht_wr_Aw_Len(i_pve_1_init_ht_axi_s_awlen),
    .pve_1_init_ht_wr_Aw_Lock(i_pve_1_init_ht_axi_s_awlock),
    .pve_1_init_ht_wr_Aw_Prot(i_pve_1_init_ht_axi_s_awprot),
    .pve_1_init_ht_wr_Aw_Ready(o_pve_1_init_ht_axi_s_awready),
    .pve_1_init_ht_wr_Aw_Size(i_pve_1_init_ht_axi_s_awsize),
    .pve_1_init_ht_wr_Aw_Valid(i_pve_1_init_ht_axi_s_awvalid),
    .pve_1_init_ht_wr_B_Id(o_pve_1_init_ht_axi_s_bid),
    .pve_1_init_ht_wr_B_Ready(i_pve_1_init_ht_axi_s_bready),
    .pve_1_init_ht_wr_B_Resp(o_pve_1_init_ht_axi_s_bresp),
    .pve_1_init_ht_wr_B_Valid(o_pve_1_init_ht_axi_s_bvalid),
    .pve_1_init_ht_wr_W_Data(i_pve_1_init_ht_axi_s_wdata),
    .pve_1_init_ht_wr_W_Last(i_pve_1_init_ht_axi_s_wlast),
    .pve_1_init_ht_wr_W_Ready(o_pve_1_init_ht_axi_s_wready),
    .pve_1_init_ht_wr_W_Strb(i_pve_1_init_ht_axi_s_wstrb),
    .pve_1_init_ht_wr_W_Valid(i_pve_1_init_ht_axi_s_wvalid),
    .pve_1_init_lt_rd_Ar_Addr(pve_1_init_lt_axi_s_araddr_msb_fixed),
    .pve_1_init_lt_rd_Ar_Burst(i_pve_1_init_lt_axi_s_arburst),
    .pve_1_init_lt_rd_Ar_Cache(i_pve_1_init_lt_axi_s_arcache),
    .pve_1_init_lt_rd_Ar_Id(i_pve_1_init_lt_axi_s_arid),
    .pve_1_init_lt_rd_Ar_Len(i_pve_1_init_lt_axi_s_arlen),
    .pve_1_init_lt_rd_Ar_Lock(i_pve_1_init_lt_axi_s_arlock),
    .pve_1_init_lt_rd_Ar_Prot(i_pve_1_init_lt_axi_s_arprot),
    .pve_1_init_lt_rd_Ar_Qos(i_pve_1_init_lt_axi_s_arqos),
    .pve_1_init_lt_rd_Ar_Ready(o_pve_1_init_lt_axi_s_arready),
    .pve_1_init_lt_rd_Ar_Size(i_pve_1_init_lt_axi_s_arsize),
    .pve_1_init_lt_rd_Ar_User(pve_1_init_lt_axi_s_aruser),
    .pve_1_init_lt_rd_Ar_Valid(i_pve_1_init_lt_axi_s_arvalid),
    .pve_1_init_lt_rd_R_Data(o_pve_1_init_lt_axi_s_rdata),
    .pve_1_init_lt_rd_R_Id(o_pve_1_init_lt_axi_s_rid),
    .pve_1_init_lt_rd_R_Last(o_pve_1_init_lt_axi_s_rlast),
    .pve_1_init_lt_rd_R_Ready(i_pve_1_init_lt_axi_s_rready),
    .pve_1_init_lt_rd_R_Resp(o_pve_1_init_lt_axi_s_rresp),
    .pve_1_init_lt_rd_R_Valid(o_pve_1_init_lt_axi_s_rvalid),
    .pve_1_init_lt_wr_Aw_Addr(pve_1_init_lt_axi_s_awaddr_msb_fixed),
    .pve_1_init_lt_wr_Aw_Burst(i_pve_1_init_lt_axi_s_awburst),
    .pve_1_init_lt_wr_Aw_Cache(i_pve_1_init_lt_axi_s_awcache),
    .pve_1_init_lt_wr_Aw_Id(i_pve_1_init_lt_axi_s_awid),
    .pve_1_init_lt_wr_Aw_Len(i_pve_1_init_lt_axi_s_awlen),
    .pve_1_init_lt_wr_Aw_Lock(i_pve_1_init_lt_axi_s_awlock),
    .pve_1_init_lt_wr_Aw_Prot(i_pve_1_init_lt_axi_s_awprot),
    .pve_1_init_lt_wr_Aw_Qos(i_pve_1_init_lt_axi_s_awqos),
    .pve_1_init_lt_wr_Aw_Ready(o_pve_1_init_lt_axi_s_awready),
    .pve_1_init_lt_wr_Aw_Size(i_pve_1_init_lt_axi_s_awsize),
    .pve_1_init_lt_wr_Aw_User(pve_1_init_lt_axi_s_awuser),
    .pve_1_init_lt_wr_Aw_Valid(i_pve_1_init_lt_axi_s_awvalid),
    .pve_1_init_lt_wr_B_Id(o_pve_1_init_lt_axi_s_bid),
    .pve_1_init_lt_wr_B_Ready(i_pve_1_init_lt_axi_s_bready),
    .pve_1_init_lt_wr_B_Resp(o_pve_1_init_lt_axi_s_bresp),
    .pve_1_init_lt_wr_B_Valid(o_pve_1_init_lt_axi_s_bvalid),
    .pve_1_init_lt_wr_W_Data(i_pve_1_init_lt_axi_s_wdata),
    .pve_1_init_lt_wr_W_Last(i_pve_1_init_lt_axi_s_wlast),
    .pve_1_init_lt_wr_W_Ready(o_pve_1_init_lt_axi_s_wready),
    .pve_1_init_lt_wr_W_Strb(i_pve_1_init_lt_axi_s_wstrb),
    .pve_1_init_lt_wr_W_Valid(i_pve_1_init_lt_axi_s_wvalid),
    .pve_1_pwr_Idle(o_pve_1_pwr_idle_val),
    .pve_1_pwr_IdleAck(o_pve_1_pwr_idle_ack),
    .pve_1_pwr_IdleReq(i_pve_1_pwr_idle_req),
    .pve_1_rst_n(i_pve_1_rst_n),
    .pve_1_targ_lt_Ar_Addr(pve_1_targ_lt_axi_m_araddr_msb_fixed),
    .pve_1_targ_lt_Ar_Burst(o_pve_1_targ_lt_axi_m_arburst),
    .pve_1_targ_lt_Ar_Cache(o_pve_1_targ_lt_axi_m_arcache),
    .pve_1_targ_lt_Ar_Id(o_pve_1_targ_lt_axi_m_arid),
    .pve_1_targ_lt_Ar_Len(o_pve_1_targ_lt_axi_m_arlen),
    .pve_1_targ_lt_Ar_Lock(o_pve_1_targ_lt_axi_m_arlock),
    .pve_1_targ_lt_Ar_Prot(o_pve_1_targ_lt_axi_m_arprot),
    .pve_1_targ_lt_Ar_Qos(o_pve_1_targ_lt_axi_m_arqos),
    .pve_1_targ_lt_Ar_Ready(i_pve_1_targ_lt_axi_m_arready),
    .pve_1_targ_lt_Ar_Size(o_pve_1_targ_lt_axi_m_arsize),
    .pve_1_targ_lt_Ar_Valid(o_pve_1_targ_lt_axi_m_arvalid),
    .pve_1_targ_lt_Aw_Addr(pve_1_targ_lt_axi_m_awaddr_msb_fixed),
    .pve_1_targ_lt_Aw_Burst(o_pve_1_targ_lt_axi_m_awburst),
    .pve_1_targ_lt_Aw_Cache(o_pve_1_targ_lt_axi_m_awcache),
    .pve_1_targ_lt_Aw_Id(o_pve_1_targ_lt_axi_m_awid),
    .pve_1_targ_lt_Aw_Len(o_pve_1_targ_lt_axi_m_awlen),
    .pve_1_targ_lt_Aw_Lock(o_pve_1_targ_lt_axi_m_awlock),
    .pve_1_targ_lt_Aw_Prot(o_pve_1_targ_lt_axi_m_awprot),
    .pve_1_targ_lt_Aw_Qos(o_pve_1_targ_lt_axi_m_awqos),
    .pve_1_targ_lt_Aw_Ready(i_pve_1_targ_lt_axi_m_awready),
    .pve_1_targ_lt_Aw_Size(o_pve_1_targ_lt_axi_m_awsize),
    .pve_1_targ_lt_Aw_Valid(o_pve_1_targ_lt_axi_m_awvalid),
    .pve_1_targ_lt_B_Id(i_pve_1_targ_lt_axi_m_bid),
    .pve_1_targ_lt_B_Ready(o_pve_1_targ_lt_axi_m_bready),
    .pve_1_targ_lt_B_Resp(i_pve_1_targ_lt_axi_m_bresp),
    .pve_1_targ_lt_B_Valid(i_pve_1_targ_lt_axi_m_bvalid),
    .pve_1_targ_lt_R_Data(i_pve_1_targ_lt_axi_m_rdata),
    .pve_1_targ_lt_R_Id(i_pve_1_targ_lt_axi_m_rid),
    .pve_1_targ_lt_R_Last(i_pve_1_targ_lt_axi_m_rlast),
    .pve_1_targ_lt_R_Ready(o_pve_1_targ_lt_axi_m_rready),
    .pve_1_targ_lt_R_Resp(i_pve_1_targ_lt_axi_m_rresp),
    .pve_1_targ_lt_R_Valid(i_pve_1_targ_lt_axi_m_rvalid),
    .pve_1_targ_lt_W_Data(o_pve_1_targ_lt_axi_m_wdata),
    .pve_1_targ_lt_W_Last(o_pve_1_targ_lt_axi_m_wlast),
    .pve_1_targ_lt_W_Ready(i_pve_1_targ_lt_axi_m_wready),
    .pve_1_targ_lt_W_Strb(o_pve_1_targ_lt_axi_m_wstrb),
    .pve_1_targ_lt_W_Valid(o_pve_1_targ_lt_axi_m_wvalid),
    .pve_1_targ_syscfg_PAddr(o_pve_1_targ_syscfg_apb_m_paddr),
    .pve_1_targ_syscfg_PEnable(o_pve_1_targ_syscfg_apb_m_penable),
    .pve_1_targ_syscfg_PProt(o_pve_1_targ_syscfg_apb_m_pprot),
    .pve_1_targ_syscfg_PRData(i_pve_1_targ_syscfg_apb_m_prdata),
    .pve_1_targ_syscfg_PReady(i_pve_1_targ_syscfg_apb_m_pready),
    .pve_1_targ_syscfg_PSel(o_pve_1_targ_syscfg_apb_m_psel),
    .pve_1_targ_syscfg_PSlvErr(i_pve_1_targ_syscfg_apb_m_pslverr),
    .pve_1_targ_syscfg_PStrb(o_pve_1_targ_syscfg_apb_m_pstrb),
    .pve_1_targ_syscfg_PWData(o_pve_1_targ_syscfg_apb_m_pwdata),
    .pve_1_targ_syscfg_PWrite(o_pve_1_targ_syscfg_apb_m_pwrite),
    .scan_en(scan_en),
    .soc_mgmt_aon_clk(i_soc_mgmt_aon_clk),
    .soc_mgmt_aon_rst_n(i_soc_mgmt_aon_rst_n),
    .soc_mgmt_clk(i_soc_mgmt_clk),
    .soc_mgmt_clken(i_soc_mgmt_clken),
    .soc_mgmt_init_lt_Ar_Addr(soc_mgmt_init_lt_axi_s_araddr_msb_fixed),
    .soc_mgmt_init_lt_Ar_Burst(i_soc_mgmt_init_lt_axi_s_arburst),
    .soc_mgmt_init_lt_Ar_Cache(i_soc_mgmt_init_lt_axi_s_arcache),
    .soc_mgmt_init_lt_Ar_Id(i_soc_mgmt_init_lt_axi_s_arid),
    .soc_mgmt_init_lt_Ar_Len(i_soc_mgmt_init_lt_axi_s_arlen),
    .soc_mgmt_init_lt_Ar_Lock(i_soc_mgmt_init_lt_axi_s_arlock),
    .soc_mgmt_init_lt_Ar_Prot(i_soc_mgmt_init_lt_axi_s_arprot),
    .soc_mgmt_init_lt_Ar_Qos(i_soc_mgmt_init_lt_axi_s_arqos),
    .soc_mgmt_init_lt_Ar_Ready(o_soc_mgmt_init_lt_axi_s_arready),
    .soc_mgmt_init_lt_Ar_Size(i_soc_mgmt_init_lt_axi_s_arsize),
    .soc_mgmt_init_lt_Ar_Valid(i_soc_mgmt_init_lt_axi_s_arvalid),
    .soc_mgmt_init_lt_Aw_Addr(soc_mgmt_init_lt_axi_s_awaddr_msb_fixed),
    .soc_mgmt_init_lt_Aw_Burst(i_soc_mgmt_init_lt_axi_s_awburst),
    .soc_mgmt_init_lt_Aw_Cache(i_soc_mgmt_init_lt_axi_s_awcache),
    .soc_mgmt_init_lt_Aw_Id(i_soc_mgmt_init_lt_axi_s_awid),
    .soc_mgmt_init_lt_Aw_Len(i_soc_mgmt_init_lt_axi_s_awlen),
    .soc_mgmt_init_lt_Aw_Lock(i_soc_mgmt_init_lt_axi_s_awlock),
    .soc_mgmt_init_lt_Aw_Prot(i_soc_mgmt_init_lt_axi_s_awprot),
    .soc_mgmt_init_lt_Aw_Qos(i_soc_mgmt_init_lt_axi_s_awqos),
    .soc_mgmt_init_lt_Aw_Ready(o_soc_mgmt_init_lt_axi_s_awready),
    .soc_mgmt_init_lt_Aw_Size(i_soc_mgmt_init_lt_axi_s_awsize),
    .soc_mgmt_init_lt_Aw_Valid(i_soc_mgmt_init_lt_axi_s_awvalid),
    .soc_mgmt_init_lt_B_Id(o_soc_mgmt_init_lt_axi_s_bid),
    .soc_mgmt_init_lt_B_Ready(i_soc_mgmt_init_lt_axi_s_bready),
    .soc_mgmt_init_lt_B_Resp(o_soc_mgmt_init_lt_axi_s_bresp),
    .soc_mgmt_init_lt_B_Valid(o_soc_mgmt_init_lt_axi_s_bvalid),
    .soc_mgmt_init_lt_R_Data(o_soc_mgmt_init_lt_axi_s_rdata),
    .soc_mgmt_init_lt_R_Id(o_soc_mgmt_init_lt_axi_s_rid),
    .soc_mgmt_init_lt_R_Last(o_soc_mgmt_init_lt_axi_s_rlast),
    .soc_mgmt_init_lt_R_Ready(i_soc_mgmt_init_lt_axi_s_rready),
    .soc_mgmt_init_lt_R_Resp(o_soc_mgmt_init_lt_axi_s_rresp),
    .soc_mgmt_init_lt_R_Valid(o_soc_mgmt_init_lt_axi_s_rvalid),
    .soc_mgmt_init_lt_W_Data(i_soc_mgmt_init_lt_axi_s_wdata),
    .soc_mgmt_init_lt_W_Last(i_soc_mgmt_init_lt_axi_s_wlast),
    .soc_mgmt_init_lt_W_Ready(o_soc_mgmt_init_lt_axi_s_wready),
    .soc_mgmt_init_lt_W_Strb(i_soc_mgmt_init_lt_axi_s_wstrb),
    .soc_mgmt_init_lt_W_Valid(i_soc_mgmt_init_lt_axi_s_wvalid),
    .soc_mgmt_pwr_Idle(o_soc_mgmt_pwr_idle_val),
    .soc_mgmt_pwr_IdleAck(o_soc_mgmt_pwr_idle_ack),
    .soc_mgmt_pwr_IdleReq(i_soc_mgmt_pwr_idle_req),
    .soc_mgmt_rst_n(i_soc_mgmt_rst_n),
    .soc_mgmt_targ_lt_Ar_Addr(soc_mgmt_targ_lt_axi_m_araddr_msb_fixed),
    .soc_mgmt_targ_lt_Ar_Burst(o_soc_mgmt_targ_lt_axi_m_arburst),
    .soc_mgmt_targ_lt_Ar_Cache(o_soc_mgmt_targ_lt_axi_m_arcache),
    .soc_mgmt_targ_lt_Ar_Id(o_soc_mgmt_targ_lt_axi_m_arid),
    .soc_mgmt_targ_lt_Ar_Len(o_soc_mgmt_targ_lt_axi_m_arlen),
    .soc_mgmt_targ_lt_Ar_Lock(o_soc_mgmt_targ_lt_axi_m_arlock),
    .soc_mgmt_targ_lt_Ar_Prot(o_soc_mgmt_targ_lt_axi_m_arprot),
    .soc_mgmt_targ_lt_Ar_Qos(o_soc_mgmt_targ_lt_axi_m_arqos),
    .soc_mgmt_targ_lt_Ar_Ready(i_soc_mgmt_targ_lt_axi_m_arready),
    .soc_mgmt_targ_lt_Ar_Size(o_soc_mgmt_targ_lt_axi_m_arsize),
    .soc_mgmt_targ_lt_Ar_Valid(o_soc_mgmt_targ_lt_axi_m_arvalid),
    .soc_mgmt_targ_lt_Aw_Addr(soc_mgmt_targ_lt_axi_m_awaddr_msb_fixed),
    .soc_mgmt_targ_lt_Aw_Burst(o_soc_mgmt_targ_lt_axi_m_awburst),
    .soc_mgmt_targ_lt_Aw_Cache(o_soc_mgmt_targ_lt_axi_m_awcache),
    .soc_mgmt_targ_lt_Aw_Id(o_soc_mgmt_targ_lt_axi_m_awid),
    .soc_mgmt_targ_lt_Aw_Len(o_soc_mgmt_targ_lt_axi_m_awlen),
    .soc_mgmt_targ_lt_Aw_Lock(o_soc_mgmt_targ_lt_axi_m_awlock),
    .soc_mgmt_targ_lt_Aw_Prot(o_soc_mgmt_targ_lt_axi_m_awprot),
    .soc_mgmt_targ_lt_Aw_Qos(o_soc_mgmt_targ_lt_axi_m_awqos),
    .soc_mgmt_targ_lt_Aw_Ready(i_soc_mgmt_targ_lt_axi_m_awready),
    .soc_mgmt_targ_lt_Aw_Size(o_soc_mgmt_targ_lt_axi_m_awsize),
    .soc_mgmt_targ_lt_Aw_Valid(o_soc_mgmt_targ_lt_axi_m_awvalid),
    .soc_mgmt_targ_lt_B_Id(i_soc_mgmt_targ_lt_axi_m_bid),
    .soc_mgmt_targ_lt_B_Ready(o_soc_mgmt_targ_lt_axi_m_bready),
    .soc_mgmt_targ_lt_B_Resp(i_soc_mgmt_targ_lt_axi_m_bresp),
    .soc_mgmt_targ_lt_B_Valid(i_soc_mgmt_targ_lt_axi_m_bvalid),
    .soc_mgmt_targ_lt_R_Data(i_soc_mgmt_targ_lt_axi_m_rdata),
    .soc_mgmt_targ_lt_R_Id(i_soc_mgmt_targ_lt_axi_m_rid),
    .soc_mgmt_targ_lt_R_Last(i_soc_mgmt_targ_lt_axi_m_rlast),
    .soc_mgmt_targ_lt_R_Ready(o_soc_mgmt_targ_lt_axi_m_rready),
    .soc_mgmt_targ_lt_R_Resp(i_soc_mgmt_targ_lt_axi_m_rresp),
    .soc_mgmt_targ_lt_R_Valid(i_soc_mgmt_targ_lt_axi_m_rvalid),
    .soc_mgmt_targ_lt_W_Data(o_soc_mgmt_targ_lt_axi_m_wdata),
    .soc_mgmt_targ_lt_W_Last(o_soc_mgmt_targ_lt_axi_m_wlast),
    .soc_mgmt_targ_lt_W_Ready(i_soc_mgmt_targ_lt_axi_m_wready),
    .soc_mgmt_targ_lt_W_Strb(o_soc_mgmt_targ_lt_axi_m_wstrb),
    .soc_mgmt_targ_lt_W_Valid(o_soc_mgmt_targ_lt_axi_m_wvalid),
    .soc_mgmt_targ_syscfg_PAddr(o_soc_mgmt_targ_syscfg_apb_m_paddr),
    .soc_mgmt_targ_syscfg_PEnable(o_soc_mgmt_targ_syscfg_apb_m_penable),
    .soc_mgmt_targ_syscfg_PProt(o_soc_mgmt_targ_syscfg_apb_m_pprot),
    .soc_mgmt_targ_syscfg_PRData(i_soc_mgmt_targ_syscfg_apb_m_prdata),
    .soc_mgmt_targ_syscfg_PReady(i_soc_mgmt_targ_syscfg_apb_m_pready),
    .soc_mgmt_targ_syscfg_PSel(o_soc_mgmt_targ_syscfg_apb_m_psel),
    .soc_mgmt_targ_syscfg_PSlvErr(i_soc_mgmt_targ_syscfg_apb_m_pslverr),
    .soc_mgmt_targ_syscfg_PStrb(o_soc_mgmt_targ_syscfg_apb_m_pstrb),
    .soc_mgmt_targ_syscfg_PWData(o_soc_mgmt_targ_syscfg_apb_m_pwdata),
    .soc_mgmt_targ_syscfg_PWrite(o_soc_mgmt_targ_syscfg_apb_m_pwrite),
    .sys_spm_aon_clk(i_sys_spm_aon_clk),
    .sys_spm_aon_rst_n(i_sys_spm_aon_rst_n),
    .sys_spm_clk(i_sys_spm_clk),
    .sys_spm_clken(i_sys_spm_clken),
    .sys_spm_pwr_Idle(o_sys_spm_pwr_idle_val),
    .sys_spm_pwr_IdleAck(o_sys_spm_pwr_idle_ack),
    .sys_spm_pwr_IdleReq(i_sys_spm_pwr_idle_req),
    .sys_spm_rst_n(i_sys_spm_rst_n),
    .sys_spm_targ_lt_Ar_Addr(sys_spm_targ_lt_axi_m_araddr_msb_fixed),
    .sys_spm_targ_lt_Ar_Burst(o_sys_spm_targ_lt_axi_m_arburst),
    .sys_spm_targ_lt_Ar_Cache(o_sys_spm_targ_lt_axi_m_arcache),
    .sys_spm_targ_lt_Ar_Id(o_sys_spm_targ_lt_axi_m_arid),
    .sys_spm_targ_lt_Ar_Len(o_sys_spm_targ_lt_axi_m_arlen),
    .sys_spm_targ_lt_Ar_Lock(o_sys_spm_targ_lt_axi_m_arlock),
    .sys_spm_targ_lt_Ar_Prot(o_sys_spm_targ_lt_axi_m_arprot),
    .sys_spm_targ_lt_Ar_Qos(o_sys_spm_targ_lt_axi_m_arqos),
    .sys_spm_targ_lt_Ar_Ready(i_sys_spm_targ_lt_axi_m_arready),
    .sys_spm_targ_lt_Ar_Size(o_sys_spm_targ_lt_axi_m_arsize),
    .sys_spm_targ_lt_Ar_Valid(o_sys_spm_targ_lt_axi_m_arvalid),
    .sys_spm_targ_lt_Aw_Addr(sys_spm_targ_lt_axi_m_awaddr_msb_fixed),
    .sys_spm_targ_lt_Aw_Burst(o_sys_spm_targ_lt_axi_m_awburst),
    .sys_spm_targ_lt_Aw_Cache(o_sys_spm_targ_lt_axi_m_awcache),
    .sys_spm_targ_lt_Aw_Id(o_sys_spm_targ_lt_axi_m_awid),
    .sys_spm_targ_lt_Aw_Len(o_sys_spm_targ_lt_axi_m_awlen),
    .sys_spm_targ_lt_Aw_Lock(o_sys_spm_targ_lt_axi_m_awlock),
    .sys_spm_targ_lt_Aw_Prot(o_sys_spm_targ_lt_axi_m_awprot),
    .sys_spm_targ_lt_Aw_Qos(o_sys_spm_targ_lt_axi_m_awqos),
    .sys_spm_targ_lt_Aw_Ready(i_sys_spm_targ_lt_axi_m_awready),
    .sys_spm_targ_lt_Aw_Size(o_sys_spm_targ_lt_axi_m_awsize),
    .sys_spm_targ_lt_Aw_Valid(o_sys_spm_targ_lt_axi_m_awvalid),
    .sys_spm_targ_lt_B_Id(i_sys_spm_targ_lt_axi_m_bid),
    .sys_spm_targ_lt_B_Ready(o_sys_spm_targ_lt_axi_m_bready),
    .sys_spm_targ_lt_B_Resp(i_sys_spm_targ_lt_axi_m_bresp),
    .sys_spm_targ_lt_B_Valid(i_sys_spm_targ_lt_axi_m_bvalid),
    .sys_spm_targ_lt_R_Data(i_sys_spm_targ_lt_axi_m_rdata),
    .sys_spm_targ_lt_R_Id(i_sys_spm_targ_lt_axi_m_rid),
    .sys_spm_targ_lt_R_Last(i_sys_spm_targ_lt_axi_m_rlast),
    .sys_spm_targ_lt_R_Ready(o_sys_spm_targ_lt_axi_m_rready),
    .sys_spm_targ_lt_R_Resp(i_sys_spm_targ_lt_axi_m_rresp),
    .sys_spm_targ_lt_R_Valid(i_sys_spm_targ_lt_axi_m_rvalid),
    .sys_spm_targ_lt_W_Data(o_sys_spm_targ_lt_axi_m_wdata),
    .sys_spm_targ_lt_W_Last(o_sys_spm_targ_lt_axi_m_wlast),
    .sys_spm_targ_lt_W_Ready(i_sys_spm_targ_lt_axi_m_wready),
    .sys_spm_targ_lt_W_Strb(o_sys_spm_targ_lt_axi_m_wstrb),
    .sys_spm_targ_lt_W_Valid(o_sys_spm_targ_lt_axi_m_wvalid),
    .sys_spm_targ_syscfg_PAddr(o_sys_spm_targ_syscfg_apb_m_paddr),
    .sys_spm_targ_syscfg_PEnable(o_sys_spm_targ_syscfg_apb_m_penable),
    .sys_spm_targ_syscfg_PProt(o_sys_spm_targ_syscfg_apb_m_pprot),
    .sys_spm_targ_syscfg_PRData(i_sys_spm_targ_syscfg_apb_m_prdata),
    .sys_spm_targ_syscfg_PReady(i_sys_spm_targ_syscfg_apb_m_pready),
    .sys_spm_targ_syscfg_PSel(o_sys_spm_targ_syscfg_apb_m_psel),
    .sys_spm_targ_syscfg_PSlvErr(i_sys_spm_targ_syscfg_apb_m_pslverr),
    .sys_spm_targ_syscfg_PStrb(o_sys_spm_targ_syscfg_apb_m_pstrb),
    .sys_spm_targ_syscfg_PWData(o_sys_spm_targ_syscfg_apb_m_pwdata),
    .sys_spm_targ_syscfg_PWrite(o_sys_spm_targ_syscfg_apb_m_pwrite)
);

endmodule
