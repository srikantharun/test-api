`ifndef SOC_MGMT_UTILS_SVH
`define SOC_MGMT_UTILS_SVH





`endif
