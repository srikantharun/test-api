// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: Wrapper for noc_h_east
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>

module noc_h_east_p (
  input logic [41:0] i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld,
  output logic [41:0] o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data,
  output logic  o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head,
  input logic  i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy,
  output logic  o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail,
  output logic  o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld,
  output logic [31:0] o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data,
  output logic  o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head,
  input logic  i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy,
  output logic  o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail,
  output logic  o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld,
  input logic [41:0] i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data,
  input logic  i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head,
  output logic  o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy,
  input logic  i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail,
  input logic  i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld,
  input logic [31:0] i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data,
  input logic  i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head,
  output logic  o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy,
  input logic  i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail,
  input logic  i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld,

    input  logic [686:0]  i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head,
    output logic          o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld,
    output logic [108:0]  o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head,
    output logic          o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld,
    output logic [108:0]  o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld,
    input  logic [146:0]  i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head,
    output logic          o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld,
    input  logic [146:0]  i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head,
    output logic          o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld,
    output logic [686:0]  o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld,
    input  logic [182:0]  i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data,
    input  logic          i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head,
    output logic          o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy,
    input  logic          i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail,
    input  logic          i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld,
    output logic [182:0]  o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data,
    output logic          o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head,
    input  logic          i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy,
    output logic          o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail,
    output logic          o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld,
    output logic [686:0]  o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data,
    output logic          o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head,
    input  logic          i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail,
    output logic          o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld,
    input  logic [108:0]  i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld,
    output logic [146:0]  o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data,
    output logic          o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head,
    input  logic          i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy,
    output logic          o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail,
    output logic          o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld,
    input  logic [686:0]  i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld,
    output logic [182:0]  o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data,
    output logic          o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head,
    input  logic          i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail,
    output logic          o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld,
    input  logic [182:0]  i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld,
    output logic [686:0]  o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld,
    input  logic [108:0]  i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld,
    output logic [686:0]  o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld,
    input  logic [108:0]  i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld,
    output logic [146:0]  o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld,
    input  logic [686:0]  i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld,
    output logic [146:0]  o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld,
    input  logic [686:0]  i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld,
    output logic [182:0]  o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data,
    output logic          o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head,
    input  logic          i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy,
    output logic          o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail,
    output logic          o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld,
    input  logic [182:0]  i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data,
    input  logic          i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head,
    output logic          o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy,
    input  logic          i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail,
    input  logic          i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld,
    input  logic [686:0]  i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data,
    input  logic          i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head,
    output logic          o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy,
    input  logic          i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail,
    input  logic          i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld,
    output logic [108:0]  o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data,
    output logic          o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head,
    input  logic          i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy,
    output logic          o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail,
    output logic          o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld,
    input  logic [146:0]  i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data,
    input  logic          i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head,
    output logic          o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy,
    input  logic          i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail,
    input  logic          i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld,
    output logic [686:0]  o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data,
    output logic          o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head,
    input  logic          i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy,
    output logic          o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail,
    output logic          o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld,
    input  logic [182:0]  i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data,
    input  logic          i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head,
    output logic          o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy,
    input  logic          i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail,
    input  logic          i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld,
    output logic [182:0]  o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data,
    output logic          o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head,
    input  logic          i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy,
    output logic          o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail,
    output logic          o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld,
    input  wire           i_noc_clk,
    input  wire           i_noc_rst_n,
    // DFT Interface
    input  wire           tck,
    input  wire           trst,
    input  logic          tms,
    input  logic          tdi,
    output logic          tdo_en,
    output logic          tdo,
    input  wire           test_clk,
    input  logic          test_mode,
    input  logic          edt_update,
    input  logic          scan_en,
    input  logic [12-1:0] scan_in,
    output logic [12-1:0] scan_out
);

    noc_h_east u_noc_h_east (
    .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data),
    .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head),
    .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy(o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy),
    .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail),
    .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld(i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld),
    .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data),
    .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head),
    .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy(i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld(o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data),
    .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head),
    .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy(o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy),
    .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail),
    .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld(i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld),
    .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data),
    .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head),
    .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy(i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld(o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data),
    .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head),
    .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy(o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy),
    .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail),
    .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld(i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld),
    .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data),
    .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head),
    .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy(i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld(o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data),
    .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head),
    .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy(o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy),
    .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail),
    .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld(i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld),
    .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data),
    .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head),
    .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy(i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld(o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data),
    .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head),
    .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy(o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy),
    .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail),
    .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld(i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld),
    .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data),
    .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head),
    .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy(i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy),
    .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail),
    .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld(o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld),
    .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data),
    .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head),
    .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy(i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy),
    .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail),
    .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld(o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld),
    .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data),
    .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head),
    .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy(o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld(i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data),
    .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head),
    .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy(i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy),
    .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail),
    .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld(o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld),
    .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data),
    .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head),
    .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy(o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld(i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data),
    .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head),
    .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy(i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy),
    .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail),
    .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld(o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld),
    .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data),
    .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head),
    .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy(o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy),
    .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail),
    .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld(i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld),
    .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data),
    .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head),
    .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy(i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy),
    .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail),
    .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld(o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld),
    .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data),
    .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head),
    .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy(o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld(i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data),
    .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head),
    .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy(i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy),
    .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail),
    .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld(o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld),
    .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data),
    .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head),
    .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy(o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy),
    .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail),
    .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld(i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld),
    .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data),
    .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head),
    .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy(i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy),
    .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail),
    .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld(o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld),
    .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data),
    .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head),
    .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy(o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld(i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data),
    .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head),
    .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy(i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy),
    .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail),
    .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld(o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld),
    .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data),
    .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head),
    .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy(o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy),
    .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail),
    .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld(i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld),
    .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data),
    .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head),
    .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy(i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy),
    .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail),
    .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld(o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld),
    .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data),
    .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head),
    .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy(o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy),
    .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail),
    .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld(i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld),
    .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data),
    .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head),
    .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy(o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy),
    .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail),
    .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld(i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld),
    .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data),
    .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head),
    .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy(i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy),
    .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail),
    .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld(o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld),
    .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data),
    .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head),
    .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy(o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy),
    .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail),
    .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld(i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld),
    .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data),
    .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head),
    .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy(i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy),
    .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail),
    .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld(o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld),
    .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data),
    .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head),
    .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy(o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy),
    .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail),
    .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld(i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld),
    .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data),
    .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head),
    .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy(i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy),
    .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail),
    .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld(o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld),
    .i_noc_clk(i_noc_clk),
    .i_noc_rst_n(i_noc_rst_n),
    .scan_en(scan_en)
    );

noc_tok_h_east u_noc_tok_h_east (
  .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data),
  .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head),
  .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy(o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy),
  .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail),
  .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld(i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld),
  .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data),
  .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head),
  .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy(o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy),
  .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail),
  .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld(i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld),
  .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data),
  .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head),
  .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy(i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy),
  .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail),
  .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld(o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld),
  .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data),
  .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head),
  .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy(i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy),
  .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail),
  .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld(o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld),
  .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data),
  .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head),
  .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy(i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy),
  .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail),
  .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld(o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld),
  .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data),
  .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head),
  .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy(i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy),
  .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail),
  .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld(o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld),
  .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data),
  .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head),
  .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy(o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy),
  .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail),
  .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld(i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld),
  .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data),
  .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head),
  .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy(o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy),
  .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail),
  .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld(i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld),
  .i_noc_clk(i_noc_clk),
  .i_noc_rst_n(i_noc_rst_n),
  .scan_en(scan_en)
);
endmodule
